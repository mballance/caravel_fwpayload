VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1992.330 84.220 1992.650 84.280 ;
        RECT 1995.090 84.220 1995.410 84.280 ;
        RECT 1992.330 84.080 1995.410 84.220 ;
        RECT 1992.330 84.020 1992.650 84.080 ;
        RECT 1995.090 84.020 1995.410 84.080 ;
        RECT 2380.110 84.220 2380.430 84.280 ;
        RECT 2414.610 84.220 2414.930 84.280 ;
        RECT 2380.110 84.080 2414.930 84.220 ;
        RECT 2380.110 84.020 2380.430 84.080 ;
        RECT 2414.610 84.020 2414.930 84.080 ;
        RECT 1800.050 83.880 1800.370 83.940 ;
        RECT 1805.570 83.880 1805.890 83.940 ;
        RECT 1800.050 83.740 1805.890 83.880 ;
        RECT 1800.050 83.680 1800.370 83.740 ;
        RECT 1805.570 83.680 1805.890 83.740 ;
        RECT 2125.270 83.540 2125.590 83.600 ;
        RECT 2172.190 83.540 2172.510 83.600 ;
        RECT 2125.270 83.400 2172.510 83.540 ;
        RECT 2125.270 83.340 2125.590 83.400 ;
        RECT 2172.190 83.340 2172.510 83.400 ;
        RECT 2221.870 83.540 2222.190 83.600 ;
        RECT 2236.130 83.540 2236.450 83.600 ;
        RECT 2221.870 83.400 2236.450 83.540 ;
        RECT 2221.870 83.340 2222.190 83.400 ;
        RECT 2236.130 83.340 2236.450 83.400 ;
      LAYER via ;
        RECT 1992.360 84.020 1992.620 84.280 ;
        RECT 1995.120 84.020 1995.380 84.280 ;
        RECT 2380.140 84.020 2380.400 84.280 ;
        RECT 2414.640 84.020 2414.900 84.280 ;
        RECT 1800.080 83.680 1800.340 83.940 ;
        RECT 1805.600 83.680 1805.860 83.940 ;
        RECT 2125.300 83.340 2125.560 83.600 ;
        RECT 2172.220 83.340 2172.480 83.600 ;
        RECT 2221.900 83.340 2222.160 83.600 ;
        RECT 2236.160 83.340 2236.420 83.600 ;
      LAYER met2 ;
        RECT 1153.705 2796.570 1153.985 2800.000 ;
        RECT 1155.150 2796.570 1155.430 2796.685 ;
        RECT 1153.705 2796.430 1155.430 2796.570 ;
        RECT 1153.705 2796.000 1153.985 2796.430 ;
        RECT 1155.150 2796.315 1155.430 2796.430 ;
        RECT 2359.430 85.155 2359.710 85.525 ;
        RECT 2173.130 84.730 2173.410 84.845 ;
        RECT 2172.280 84.590 2173.410 84.730 ;
        RECT 1992.360 84.165 1992.620 84.310 ;
        RECT 1995.120 84.165 1995.380 84.310 ;
        RECT 1800.070 83.795 1800.350 84.165 ;
        RECT 1805.590 83.795 1805.870 84.165 ;
        RECT 1992.350 83.795 1992.630 84.165 ;
        RECT 1995.110 83.795 1995.390 84.165 ;
        RECT 2089.410 83.795 2089.690 84.165 ;
        RECT 1800.080 83.650 1800.340 83.795 ;
        RECT 1805.600 83.650 1805.860 83.795 ;
        RECT 2089.480 82.125 2089.620 83.795 ;
        RECT 2172.280 83.630 2172.420 84.590 ;
        RECT 2173.130 84.475 2173.410 84.590 ;
        RECT 2236.150 84.475 2236.430 84.845 ;
        RECT 2236.220 83.630 2236.360 84.475 ;
        RECT 2125.300 83.485 2125.560 83.630 ;
        RECT 2125.290 83.115 2125.570 83.485 ;
        RECT 2172.220 83.310 2172.480 83.630 ;
        RECT 2221.900 83.485 2222.160 83.630 ;
        RECT 2221.890 83.115 2222.170 83.485 ;
        RECT 2236.160 83.310 2236.420 83.630 ;
        RECT 2359.500 83.485 2359.640 85.155 ;
        RECT 2414.630 84.475 2414.910 84.845 ;
        RECT 2414.700 84.310 2414.840 84.475 ;
        RECT 2380.140 84.165 2380.400 84.310 ;
        RECT 2380.130 83.795 2380.410 84.165 ;
        RECT 2414.640 83.990 2414.900 84.310 ;
        RECT 2359.430 83.115 2359.710 83.485 ;
        RECT 2089.410 81.755 2089.690 82.125 ;
      LAYER via2 ;
        RECT 1155.150 2796.360 1155.430 2796.640 ;
        RECT 2359.430 85.200 2359.710 85.480 ;
        RECT 1800.070 83.840 1800.350 84.120 ;
        RECT 1805.590 83.840 1805.870 84.120 ;
        RECT 1992.350 83.840 1992.630 84.120 ;
        RECT 1995.110 83.840 1995.390 84.120 ;
        RECT 2089.410 83.840 2089.690 84.120 ;
        RECT 2173.130 84.520 2173.410 84.800 ;
        RECT 2236.150 84.520 2236.430 84.800 ;
        RECT 2125.290 83.160 2125.570 83.440 ;
        RECT 2221.890 83.160 2222.170 83.440 ;
        RECT 2414.630 84.520 2414.910 84.800 ;
        RECT 2380.130 83.840 2380.410 84.120 ;
        RECT 2359.430 83.160 2359.710 83.440 ;
        RECT 2089.410 81.800 2089.690 82.080 ;
      LAYER met3 ;
        RECT 1155.125 2796.650 1155.455 2796.665 ;
        RECT 1158.550 2796.650 1158.930 2796.660 ;
        RECT 1155.125 2796.350 1158.930 2796.650 ;
        RECT 1155.125 2796.335 1155.455 2796.350 ;
        RECT 1158.550 2796.340 1158.930 2796.350 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 2311.310 85.490 2311.690 85.500 ;
        RECT 2359.405 85.490 2359.735 85.505 ;
        RECT 1883.550 85.190 1931.690 85.490 ;
        RECT 1800.045 84.130 1800.375 84.145 ;
        RECT 1752.910 83.830 1800.375 84.130 ;
        RECT 1158.550 83.450 1158.930 83.460 ;
        RECT 1752.910 83.450 1753.210 83.830 ;
        RECT 1800.045 83.815 1800.375 83.830 ;
        RECT 1805.565 84.130 1805.895 84.145 ;
        RECT 1883.550 84.130 1883.850 85.190 ;
        RECT 1805.565 83.830 1835.090 84.130 ;
        RECT 1805.565 83.815 1805.895 83.830 ;
        RECT 1158.550 83.150 1753.210 83.450 ;
        RECT 1834.790 83.450 1835.090 83.830 ;
        RECT 1849.510 83.830 1883.850 84.130 ;
        RECT 1849.510 83.450 1849.810 83.830 ;
        RECT 1834.790 83.150 1849.810 83.450 ;
        RECT 1931.390 83.450 1931.690 85.190 ;
        RECT 2311.310 85.190 2359.735 85.490 ;
        RECT 2311.310 85.180 2311.690 85.190 ;
        RECT 2359.405 85.175 2359.735 85.190 ;
        RECT 2173.105 84.810 2173.435 84.825 ;
        RECT 2236.125 84.810 2236.455 84.825 ;
        RECT 2414.605 84.810 2414.935 84.825 ;
        RECT 2173.105 84.510 2187.450 84.810 ;
        RECT 2173.105 84.495 2173.435 84.510 ;
        RECT 1992.325 84.130 1992.655 84.145 ;
        RECT 1946.110 83.830 1992.655 84.130 ;
        RECT 1946.110 83.450 1946.410 83.830 ;
        RECT 1992.325 83.815 1992.655 83.830 ;
        RECT 1995.085 84.130 1995.415 84.145 ;
        RECT 2089.385 84.130 2089.715 84.145 ;
        RECT 1995.085 83.830 2028.290 84.130 ;
        RECT 1995.085 83.815 1995.415 83.830 ;
        RECT 1931.390 83.150 1946.410 83.450 ;
        RECT 2027.990 83.450 2028.290 83.830 ;
        RECT 2042.710 83.830 2089.715 84.130 ;
        RECT 2042.710 83.450 2043.010 83.830 ;
        RECT 2089.385 83.815 2089.715 83.830 ;
        RECT 2125.265 83.450 2125.595 83.465 ;
        RECT 2027.990 83.150 2043.010 83.450 ;
        RECT 2124.590 83.150 2125.595 83.450 ;
        RECT 2187.150 83.450 2187.450 84.510 ;
        RECT 2236.125 84.510 2294.170 84.810 ;
        RECT 2236.125 84.495 2236.455 84.510 ;
        RECT 2293.870 84.130 2294.170 84.510 ;
        RECT 2414.605 84.510 2449.650 84.810 ;
        RECT 2414.605 84.495 2414.935 84.510 ;
        RECT 2311.310 84.130 2311.690 84.140 ;
        RECT 2380.105 84.130 2380.435 84.145 ;
        RECT 2293.870 83.830 2311.690 84.130 ;
        RECT 2311.310 83.820 2311.690 83.830 ;
        RECT 2366.550 83.830 2380.435 84.130 ;
        RECT 2449.350 84.130 2449.650 84.510 ;
        RECT 2498.110 84.510 2546.250 84.810 ;
        RECT 2449.350 83.830 2497.490 84.130 ;
        RECT 2221.865 83.450 2222.195 83.465 ;
        RECT 2187.150 83.150 2222.195 83.450 ;
        RECT 1158.550 83.140 1158.930 83.150 ;
        RECT 2089.385 82.090 2089.715 82.105 ;
        RECT 2124.590 82.090 2124.890 83.150 ;
        RECT 2125.265 83.135 2125.595 83.150 ;
        RECT 2221.865 83.135 2222.195 83.150 ;
        RECT 2359.405 83.450 2359.735 83.465 ;
        RECT 2366.550 83.450 2366.850 83.830 ;
        RECT 2380.105 83.815 2380.435 83.830 ;
        RECT 2359.405 83.150 2366.850 83.450 ;
        RECT 2497.190 83.450 2497.490 83.830 ;
        RECT 2498.110 83.450 2498.410 84.510 ;
        RECT 2545.950 84.130 2546.250 84.510 ;
        RECT 2594.710 84.510 2642.850 84.810 ;
        RECT 2545.950 83.830 2594.090 84.130 ;
        RECT 2497.190 83.150 2498.410 83.450 ;
        RECT 2593.790 83.450 2594.090 83.830 ;
        RECT 2594.710 83.450 2595.010 84.510 ;
        RECT 2642.550 84.130 2642.850 84.510 ;
        RECT 2691.310 84.510 2739.450 84.810 ;
        RECT 2642.550 83.830 2690.690 84.130 ;
        RECT 2593.790 83.150 2595.010 83.450 ;
        RECT 2690.390 83.450 2690.690 83.830 ;
        RECT 2691.310 83.450 2691.610 84.510 ;
        RECT 2739.150 84.130 2739.450 84.510 ;
        RECT 2787.910 84.510 2836.050 84.810 ;
        RECT 2739.150 83.830 2787.290 84.130 ;
        RECT 2690.390 83.150 2691.610 83.450 ;
        RECT 2786.990 83.450 2787.290 83.830 ;
        RECT 2787.910 83.450 2788.210 84.510 ;
        RECT 2835.750 84.130 2836.050 84.510 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2835.750 83.830 2883.890 84.130 ;
        RECT 2786.990 83.150 2788.210 83.450 ;
        RECT 2883.590 83.450 2883.890 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2883.590 83.150 2884.810 83.450 ;
        RECT 2359.405 83.135 2359.735 83.150 ;
        RECT 2089.385 81.790 2124.890 82.090 ;
        RECT 2089.385 81.775 2089.715 81.790 ;
      LAYER via3 ;
        RECT 1158.580 2796.340 1158.900 2796.660 ;
        RECT 1158.580 83.140 1158.900 83.460 ;
        RECT 2311.340 85.180 2311.660 85.500 ;
        RECT 2311.340 83.820 2311.660 84.140 ;
      LAYER met4 ;
        RECT 1158.575 2796.335 1158.905 2796.665 ;
        RECT 1158.590 83.465 1158.890 2796.335 ;
        RECT 2311.335 85.175 2311.665 85.505 ;
        RECT 2311.350 84.145 2311.650 85.175 ;
        RECT 2311.335 83.815 2311.665 84.145 ;
        RECT 1158.575 83.135 1158.905 83.465 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1443.110 2814.675 1443.390 2815.045 ;
        RECT 1443.180 2800.000 1443.320 2814.675 ;
        RECT 1443.045 2796.000 1443.325 2800.000 ;
      LAYER via2 ;
        RECT 1443.110 2814.720 1443.390 2815.000 ;
      LAYER met3 ;
        RECT 1443.085 2815.010 1443.415 2815.025 ;
        RECT 2231.270 2815.010 2231.650 2815.020 ;
        RECT 1443.085 2814.710 2231.650 2815.010 ;
        RECT 1443.085 2814.695 1443.415 2814.710 ;
        RECT 2231.270 2814.700 2231.650 2814.710 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2916.710 2433.910 2924.800 2434.210 ;
        RECT 2231.270 2430.810 2231.650 2430.820 ;
        RECT 2231.270 2430.510 2256.450 2430.810 ;
        RECT 2231.270 2430.500 2231.650 2430.510 ;
        RECT 2256.150 2430.130 2256.450 2430.510 ;
        RECT 2304.910 2430.510 2353.050 2430.810 ;
        RECT 2256.150 2429.830 2304.290 2430.130 ;
        RECT 2303.990 2429.450 2304.290 2429.830 ;
        RECT 2304.910 2429.450 2305.210 2430.510 ;
        RECT 2352.750 2430.130 2353.050 2430.510 ;
        RECT 2401.510 2430.510 2449.650 2430.810 ;
        RECT 2352.750 2429.830 2400.890 2430.130 ;
        RECT 2303.990 2429.150 2305.210 2429.450 ;
        RECT 2400.590 2429.450 2400.890 2429.830 ;
        RECT 2401.510 2429.450 2401.810 2430.510 ;
        RECT 2449.350 2430.130 2449.650 2430.510 ;
        RECT 2498.110 2430.510 2546.250 2430.810 ;
        RECT 2449.350 2429.830 2497.490 2430.130 ;
        RECT 2400.590 2429.150 2401.810 2429.450 ;
        RECT 2497.190 2429.450 2497.490 2429.830 ;
        RECT 2498.110 2429.450 2498.410 2430.510 ;
        RECT 2545.950 2430.130 2546.250 2430.510 ;
        RECT 2594.710 2430.510 2642.850 2430.810 ;
        RECT 2545.950 2429.830 2594.090 2430.130 ;
        RECT 2497.190 2429.150 2498.410 2429.450 ;
        RECT 2593.790 2429.450 2594.090 2429.830 ;
        RECT 2594.710 2429.450 2595.010 2430.510 ;
        RECT 2642.550 2430.130 2642.850 2430.510 ;
        RECT 2691.310 2430.510 2739.450 2430.810 ;
        RECT 2642.550 2429.830 2690.690 2430.130 ;
        RECT 2593.790 2429.150 2595.010 2429.450 ;
        RECT 2690.390 2429.450 2690.690 2429.830 ;
        RECT 2691.310 2429.450 2691.610 2430.510 ;
        RECT 2739.150 2430.130 2739.450 2430.510 ;
        RECT 2787.910 2430.510 2836.050 2430.810 ;
        RECT 2739.150 2429.830 2787.290 2430.130 ;
        RECT 2690.390 2429.150 2691.610 2429.450 ;
        RECT 2786.990 2429.450 2787.290 2429.830 ;
        RECT 2787.910 2429.450 2788.210 2430.510 ;
        RECT 2835.750 2430.130 2836.050 2430.510 ;
        RECT 2916.710 2430.130 2917.010 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2835.750 2429.830 2883.890 2430.130 ;
        RECT 2786.990 2429.150 2788.210 2429.450 ;
        RECT 2883.590 2429.450 2883.890 2429.830 ;
        RECT 2884.510 2429.830 2917.010 2430.130 ;
        RECT 2884.510 2429.450 2884.810 2429.830 ;
        RECT 2883.590 2429.150 2884.810 2429.450 ;
      LAYER via3 ;
        RECT 2231.300 2814.700 2231.620 2815.020 ;
        RECT 2231.300 2430.500 2231.620 2430.820 ;
      LAYER met4 ;
        RECT 2231.295 2814.695 2231.625 2815.025 ;
        RECT 2231.310 2430.825 2231.610 2814.695 ;
        RECT 2231.295 2430.495 2231.625 2430.825 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2001.145 2803.045 2002.235 2803.215 ;
      LAYER mcon ;
        RECT 2002.065 2803.045 2002.235 2803.215 ;
      LAYER met1 ;
        RECT 1472.070 2803.200 1472.390 2803.260 ;
        RECT 2001.085 2803.200 2001.375 2803.245 ;
        RECT 1472.070 2803.060 2001.375 2803.200 ;
        RECT 1472.070 2803.000 1472.390 2803.060 ;
        RECT 2001.085 2803.015 2001.375 2803.060 ;
        RECT 2002.005 2803.200 2002.295 2803.245 ;
        RECT 2742.590 2803.200 2742.910 2803.260 ;
        RECT 2002.005 2803.060 2742.910 2803.200 ;
        RECT 2002.005 2803.015 2002.295 2803.060 ;
        RECT 2742.590 2803.000 2742.910 2803.060 ;
        RECT 2742.590 2670.260 2742.910 2670.320 ;
        RECT 2898.990 2670.260 2899.310 2670.320 ;
        RECT 2742.590 2670.120 2899.310 2670.260 ;
        RECT 2742.590 2670.060 2742.910 2670.120 ;
        RECT 2898.990 2670.060 2899.310 2670.120 ;
      LAYER via ;
        RECT 1472.100 2803.000 1472.360 2803.260 ;
        RECT 2742.620 2803.000 2742.880 2803.260 ;
        RECT 2742.620 2670.060 2742.880 2670.320 ;
        RECT 2899.020 2670.060 2899.280 2670.320 ;
      LAYER met2 ;
        RECT 1472.100 2802.970 1472.360 2803.290 ;
        RECT 2742.620 2802.970 2742.880 2803.290 ;
        RECT 1472.160 2800.000 1472.300 2802.970 ;
        RECT 1472.025 2796.000 1472.305 2800.000 ;
        RECT 2742.680 2670.350 2742.820 2802.970 ;
        RECT 2742.620 2670.030 2742.880 2670.350 ;
        RECT 2899.020 2670.030 2899.280 2670.350 ;
        RECT 2899.080 2669.525 2899.220 2670.030 ;
        RECT 2899.010 2669.155 2899.290 2669.525 ;
      LAYER via2 ;
        RECT 2899.010 2669.200 2899.290 2669.480 ;
      LAYER met3 ;
        RECT 2898.985 2669.490 2899.315 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2898.985 2669.190 2924.800 2669.490 ;
        RECT 2898.985 2669.175 2899.315 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2125.360 2898.600 2149.420 2898.740 ;
        RECT 1503.350 2898.400 1503.670 2898.460 ;
        RECT 2125.360 2898.400 2125.500 2898.600 ;
        RECT 1503.350 2898.260 2125.500 2898.400 ;
        RECT 2149.280 2898.400 2149.420 2898.600 ;
        RECT 2469.900 2898.600 2471.420 2898.740 ;
        RECT 2469.900 2898.400 2470.040 2898.600 ;
        RECT 2149.280 2898.260 2470.040 2898.400 ;
        RECT 2471.280 2898.400 2471.420 2898.600 ;
        RECT 2777.180 2898.600 2797.100 2898.740 ;
        RECT 2777.180 2898.400 2777.320 2898.600 ;
        RECT 2471.280 2898.260 2777.320 2898.400 ;
        RECT 2796.960 2898.400 2797.100 2898.600 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2796.960 2898.260 2901.150 2898.400 ;
        RECT 1503.350 2898.200 1503.670 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 1503.380 2898.200 1503.640 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1503.380 2898.170 1503.640 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1501.005 2799.970 1501.285 2800.000 ;
        RECT 1503.440 2799.970 1503.580 2898.170 ;
        RECT 1501.005 2799.830 1503.580 2799.970 ;
        RECT 1501.005 2796.000 1501.285 2799.830 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.410 3133.000 1531.730 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1531.410 3132.860 2901.150 3133.000 ;
        RECT 1531.410 3132.800 1531.730 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1531.440 3132.800 1531.700 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1531.440 3132.770 1531.700 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1529.525 2799.970 1529.805 2800.000 ;
        RECT 1531.500 2799.970 1531.640 3132.770 ;
        RECT 1529.525 2799.830 1531.640 2799.970 ;
        RECT 1529.525 2796.000 1529.805 2799.830 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.010 3367.600 1559.330 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1559.010 3367.460 2901.150 3367.600 ;
        RECT 1559.010 3367.400 1559.330 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 1552.570 2825.640 1552.890 2825.700 ;
        RECT 1559.010 2825.640 1559.330 2825.700 ;
        RECT 1552.570 2825.500 1559.330 2825.640 ;
        RECT 1552.570 2825.440 1552.890 2825.500 ;
        RECT 1559.010 2825.440 1559.330 2825.500 ;
        RECT 1552.570 2814.760 1552.890 2814.820 ;
        RECT 1558.550 2814.760 1558.870 2814.820 ;
        RECT 1552.570 2814.620 1558.870 2814.760 ;
        RECT 1552.570 2814.560 1552.890 2814.620 ;
        RECT 1558.550 2814.560 1558.870 2814.620 ;
      LAYER via ;
        RECT 1559.040 3367.400 1559.300 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 1552.600 2825.440 1552.860 2825.700 ;
        RECT 1559.040 2825.440 1559.300 2825.700 ;
        RECT 1552.600 2814.560 1552.860 2814.820 ;
        RECT 1558.580 2814.560 1558.840 2814.820 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1559.040 3367.370 1559.300 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1559.100 2825.730 1559.240 3367.370 ;
        RECT 1552.600 2825.410 1552.860 2825.730 ;
        RECT 1559.040 2825.410 1559.300 2825.730 ;
        RECT 1552.660 2814.850 1552.800 2825.410 ;
        RECT 1552.600 2814.530 1552.860 2814.850 ;
        RECT 1558.580 2814.530 1558.840 2814.850 ;
        RECT 1558.640 2800.000 1558.780 2814.530 ;
        RECT 1558.505 2796.000 1558.785 2800.000 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3422.355 ;
        RECT 2795.565 3008.405 2795.735 3042.915 ;
        RECT 2796.485 2946.525 2796.655 2994.635 ;
        RECT 2796.485 2849.625 2796.655 2898.075 ;
      LAYER mcon ;
        RECT 2796.485 3422.185 2796.655 3422.355 ;
        RECT 2795.565 3042.745 2795.735 3042.915 ;
        RECT 2796.485 2994.465 2796.655 2994.635 ;
        RECT 2796.485 2897.905 2796.655 2898.075 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2796.425 3422.340 2796.715 3422.385 ;
        RECT 2795.030 3422.200 2796.715 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2796.425 3422.155 2796.715 3422.200 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.295 3042.760 2795.810 3042.900 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.505 3008.560 2795.795 3008.605 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.505 3008.420 2796.730 3008.560 ;
        RECT 2795.505 3008.375 2795.795 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2796.215 2994.480 2796.730 2994.620 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2796.425 2946.680 2796.715 2946.725 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2796.425 2946.540 2797.190 2946.680 ;
        RECT 2796.425 2946.495 2796.715 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.410 2898.060 2796.730 2898.120 ;
        RECT 2796.215 2897.920 2796.730 2898.060 ;
        RECT 2796.410 2897.860 2796.730 2897.920 ;
        RECT 2796.425 2849.780 2796.715 2849.825 ;
        RECT 2796.870 2849.780 2797.190 2849.840 ;
        RECT 2796.425 2849.640 2797.190 2849.780 ;
        RECT 2796.425 2849.595 2796.715 2849.640 ;
        RECT 2796.870 2849.580 2797.190 2849.640 ;
        RECT 1587.530 2818.500 1587.850 2818.560 ;
        RECT 2796.870 2818.500 2797.190 2818.560 ;
        RECT 1587.530 2818.360 2797.190 2818.500 ;
        RECT 1587.530 2818.300 1587.850 2818.360 ;
        RECT 2796.870 2818.300 2797.190 2818.360 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.440 2897.860 2796.700 2898.120 ;
        RECT 2796.900 2849.580 2797.160 2849.840 ;
        RECT 1587.560 2818.300 1587.820 2818.560 ;
        RECT 2796.900 2818.300 2797.160 2818.560 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2922.370 2797.100 2946.450 ;
        RECT 2796.040 2922.230 2797.100 2922.370 ;
        RECT 2796.040 2898.570 2796.180 2922.230 ;
        RECT 2796.040 2898.430 2796.640 2898.570 ;
        RECT 2796.500 2898.150 2796.640 2898.430 ;
        RECT 2796.440 2897.830 2796.700 2898.150 ;
        RECT 2796.900 2849.550 2797.160 2849.870 ;
        RECT 2796.960 2818.590 2797.100 2849.550 ;
        RECT 1587.560 2818.270 1587.820 2818.590 ;
        RECT 2796.900 2818.270 2797.160 2818.590 ;
        RECT 1587.620 2800.000 1587.760 2818.270 ;
        RECT 1587.485 2796.000 1587.765 2800.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
        RECT 2470.345 2849.625 2470.515 2898.075 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
        RECT 2470.345 2897.905 2470.515 2898.075 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2470.270 2898.060 2470.590 2898.120 ;
        RECT 2470.075 2897.920 2470.590 2898.060 ;
        RECT 2470.270 2897.860 2470.590 2897.920 ;
        RECT 2470.285 2849.780 2470.575 2849.825 ;
        RECT 2471.190 2849.780 2471.510 2849.840 ;
        RECT 2470.285 2849.640 2471.510 2849.780 ;
        RECT 2470.285 2849.595 2470.575 2849.640 ;
        RECT 2471.190 2849.580 2471.510 2849.640 ;
        RECT 1616.510 2818.840 1616.830 2818.900 ;
        RECT 2471.190 2818.840 2471.510 2818.900 ;
        RECT 1616.510 2818.700 2471.510 2818.840 ;
        RECT 1616.510 2818.640 1616.830 2818.700 ;
        RECT 2471.190 2818.640 2471.510 2818.700 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2470.300 2897.860 2470.560 2898.120 ;
        RECT 2471.220 2849.580 2471.480 2849.840 ;
        RECT 1616.540 2818.640 1616.800 2818.900 ;
        RECT 2471.220 2818.640 2471.480 2818.900 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2898.570 2470.960 2959.630 ;
        RECT 2470.360 2898.430 2470.960 2898.570 ;
        RECT 2470.360 2898.150 2470.500 2898.430 ;
        RECT 2470.300 2897.830 2470.560 2898.150 ;
        RECT 2471.220 2849.550 2471.480 2849.870 ;
        RECT 2471.280 2818.930 2471.420 2849.550 ;
        RECT 1616.540 2818.610 1616.800 2818.930 ;
        RECT 2471.220 2818.610 2471.480 2818.930 ;
        RECT 1616.600 2800.000 1616.740 2818.610 ;
        RECT 1616.465 2796.000 1616.745 2800.000 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3422.355 ;
        RECT 2146.965 3008.405 2147.135 3042.915 ;
        RECT 2147.885 2946.525 2148.055 2994.635 ;
        RECT 2147.425 2849.625 2147.595 2898.075 ;
      LAYER mcon ;
        RECT 2147.885 3422.185 2148.055 3422.355 ;
        RECT 2146.965 3042.745 2147.135 3042.915 ;
        RECT 2147.885 2994.465 2148.055 2994.635 ;
        RECT 2147.425 2897.905 2147.595 2898.075 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.825 3422.340 2148.115 3422.385 ;
        RECT 2146.430 3422.200 2148.115 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.825 3422.155 2148.115 3422.200 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.695 3042.760 2147.210 3042.900 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.905 3008.560 2147.195 3008.605 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.905 3008.420 2148.130 3008.560 ;
        RECT 2146.905 3008.375 2147.195 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2147.810 2994.620 2148.130 2994.680 ;
        RECT 2147.615 2994.480 2148.130 2994.620 ;
        RECT 2147.810 2994.420 2148.130 2994.480 ;
        RECT 2147.825 2946.680 2148.115 2946.725 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2147.825 2946.540 2148.590 2946.680 ;
        RECT 2147.825 2946.495 2148.115 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 2147.365 2898.060 2147.655 2898.105 ;
        RECT 2147.810 2898.060 2148.130 2898.120 ;
        RECT 2147.365 2897.920 2148.130 2898.060 ;
        RECT 2147.365 2897.875 2147.655 2897.920 ;
        RECT 2147.810 2897.860 2148.130 2897.920 ;
        RECT 2147.350 2849.780 2147.670 2849.840 ;
        RECT 2147.155 2849.640 2147.670 2849.780 ;
        RECT 2147.350 2849.580 2147.670 2849.640 ;
        RECT 1642.270 2819.180 1642.590 2819.240 ;
        RECT 2147.350 2819.180 2147.670 2819.240 ;
        RECT 1642.270 2819.040 2147.670 2819.180 ;
        RECT 1642.270 2818.980 1642.590 2819.040 ;
        RECT 2147.350 2818.980 2147.670 2819.040 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2147.840 2994.420 2148.100 2994.680 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 2147.840 2897.860 2148.100 2898.120 ;
        RECT 2147.380 2849.580 2147.640 2849.840 ;
        RECT 1642.300 2818.980 1642.560 2819.240 ;
        RECT 2147.380 2818.980 2147.640 2819.240 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2994.710 2148.040 3008.330 ;
        RECT 2147.840 2994.390 2148.100 2994.710 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2922.370 2148.500 2946.450 ;
        RECT 2147.440 2922.230 2148.500 2922.370 ;
        RECT 2147.440 2898.570 2147.580 2922.230 ;
        RECT 2147.440 2898.430 2148.040 2898.570 ;
        RECT 2147.900 2898.150 2148.040 2898.430 ;
        RECT 2147.840 2897.830 2148.100 2898.150 ;
        RECT 2147.380 2849.550 2147.640 2849.870 ;
        RECT 2147.440 2819.270 2147.580 2849.550 ;
        RECT 1642.300 2818.950 1642.560 2819.270 ;
        RECT 2147.380 2818.950 2147.640 2819.270 ;
        RECT 1642.360 2800.650 1642.500 2818.950 ;
        RECT 1642.360 2800.510 1644.340 2800.650 ;
        RECT 1644.200 2799.970 1644.340 2800.510 ;
        RECT 1645.445 2799.970 1645.725 2800.000 ;
        RECT 1644.200 2799.830 1645.725 2799.970 ;
        RECT 1645.445 2796.000 1645.725 2799.830 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1742.090 3501.220 1742.410 3501.280 ;
        RECT 1824.890 3501.220 1825.210 3501.280 ;
        RECT 1742.090 3501.080 1825.210 3501.220 ;
        RECT 1742.090 3501.020 1742.410 3501.080 ;
        RECT 1824.890 3501.020 1825.210 3501.080 ;
        RECT 1669.870 2819.860 1670.190 2819.920 ;
        RECT 1742.090 2819.860 1742.410 2819.920 ;
        RECT 1669.870 2819.720 1742.410 2819.860 ;
        RECT 1669.870 2819.660 1670.190 2819.720 ;
        RECT 1742.090 2819.660 1742.410 2819.720 ;
      LAYER via ;
        RECT 1742.120 3501.020 1742.380 3501.280 ;
        RECT 1824.920 3501.020 1825.180 3501.280 ;
        RECT 1669.900 2819.660 1670.160 2819.920 ;
        RECT 1742.120 2819.660 1742.380 2819.920 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3501.310 1825.120 3517.600 ;
        RECT 1742.120 3500.990 1742.380 3501.310 ;
        RECT 1824.920 3500.990 1825.180 3501.310 ;
        RECT 1742.180 2819.950 1742.320 3500.990 ;
        RECT 1669.900 2819.630 1670.160 2819.950 ;
        RECT 1742.120 2819.630 1742.380 2819.950 ;
        RECT 1669.960 2800.650 1670.100 2819.630 ;
        RECT 1669.960 2800.510 1672.860 2800.650 ;
        RECT 1672.720 2799.970 1672.860 2800.510 ;
        RECT 1674.425 2799.970 1674.705 2800.000 ;
        RECT 1672.720 2799.830 1674.705 2799.970 ;
        RECT 1674.425 2796.000 1674.705 2799.830 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 2819.520 1504.130 2819.580 ;
        RECT 1703.450 2819.520 1703.770 2819.580 ;
        RECT 1503.810 2819.380 1703.770 2819.520 ;
        RECT 1503.810 2819.320 1504.130 2819.380 ;
        RECT 1703.450 2819.320 1703.770 2819.380 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 2819.320 1504.100 2819.580 ;
        RECT 1703.480 2819.320 1703.740 2819.580 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 2819.610 1504.040 3498.270 ;
        RECT 1503.840 2819.290 1504.100 2819.610 ;
        RECT 1703.480 2819.290 1703.740 2819.610 ;
        RECT 1703.540 2800.000 1703.680 2819.290 ;
        RECT 1703.405 2796.000 1703.685 2800.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1633.990 318.820 1634.310 318.880 ;
        RECT 1676.310 318.820 1676.630 318.880 ;
        RECT 1633.990 318.680 1676.630 318.820 ;
        RECT 1633.990 318.620 1634.310 318.680 ;
        RECT 1676.310 318.620 1676.630 318.680 ;
        RECT 1992.330 318.820 1992.650 318.880 ;
        RECT 1995.090 318.820 1995.410 318.880 ;
        RECT 1992.330 318.680 1995.410 318.820 ;
        RECT 1992.330 318.620 1992.650 318.680 ;
        RECT 1995.090 318.620 1995.410 318.680 ;
        RECT 1797.750 318.480 1798.070 318.540 ;
        RECT 1828.110 318.480 1828.430 318.540 ;
        RECT 1797.750 318.340 1828.430 318.480 ;
        RECT 1797.750 318.280 1798.070 318.340 ;
        RECT 1828.110 318.280 1828.430 318.340 ;
        RECT 2089.390 318.480 2089.710 318.540 ;
        RECT 2098.130 318.480 2098.450 318.540 ;
        RECT 2089.390 318.340 2098.450 318.480 ;
        RECT 2089.390 318.280 2089.710 318.340 ;
        RECT 2098.130 318.280 2098.450 318.340 ;
      LAYER via ;
        RECT 1634.020 318.620 1634.280 318.880 ;
        RECT 1676.340 318.620 1676.600 318.880 ;
        RECT 1992.360 318.620 1992.620 318.880 ;
        RECT 1995.120 318.620 1995.380 318.880 ;
        RECT 1797.780 318.280 1798.040 318.540 ;
        RECT 1828.140 318.280 1828.400 318.540 ;
        RECT 2089.420 318.280 2089.680 318.540 ;
        RECT 2098.160 318.280 2098.420 318.540 ;
      LAYER met2 ;
        RECT 1182.225 2796.570 1182.505 2800.000 ;
        RECT 1183.670 2796.570 1183.950 2796.685 ;
        RECT 1182.225 2796.430 1183.950 2796.570 ;
        RECT 1182.225 2796.000 1182.505 2796.430 ;
        RECT 1183.670 2796.315 1183.950 2796.430 ;
        RECT 2304.230 321.115 2304.510 321.485 ;
        RECT 1741.650 319.755 1741.930 320.125 ;
        RECT 2236.150 319.755 2236.430 320.125 ;
        RECT 1364.910 319.330 1365.190 319.445 ;
        RECT 1365.830 319.330 1366.110 319.445 ;
        RECT 1364.910 319.190 1366.110 319.330 ;
        RECT 1364.910 319.075 1365.190 319.190 ;
        RECT 1365.830 319.075 1366.110 319.190 ;
        RECT 1676.330 319.075 1676.610 319.445 ;
        RECT 1676.400 318.910 1676.540 319.075 ;
        RECT 1634.020 318.765 1634.280 318.910 ;
        RECT 1634.010 318.395 1634.290 318.765 ;
        RECT 1676.340 318.590 1676.600 318.910 ;
        RECT 1741.720 318.765 1741.860 319.755 ;
        RECT 1992.360 318.765 1992.620 318.910 ;
        RECT 1995.120 318.765 1995.380 318.910 ;
        RECT 1741.650 318.395 1741.930 318.765 ;
        RECT 1797.770 318.395 1798.050 318.765 ;
        RECT 1797.780 318.250 1798.040 318.395 ;
        RECT 1828.140 318.250 1828.400 318.570 ;
        RECT 1992.350 318.395 1992.630 318.765 ;
        RECT 1995.110 318.395 1995.390 318.765 ;
        RECT 2089.410 318.395 2089.690 318.765 ;
        RECT 2098.150 318.395 2098.430 318.765 ;
        RECT 2235.690 318.650 2235.970 318.765 ;
        RECT 2236.220 318.650 2236.360 319.755 ;
        RECT 2304.300 319.445 2304.440 321.115 ;
        RECT 2304.230 319.075 2304.510 319.445 ;
        RECT 2235.690 318.510 2236.360 318.650 ;
        RECT 2235.690 318.395 2235.970 318.510 ;
        RECT 2089.420 318.250 2089.680 318.395 ;
        RECT 2098.160 318.250 2098.420 318.395 ;
        RECT 1828.200 318.085 1828.340 318.250 ;
        RECT 1828.130 317.715 1828.410 318.085 ;
      LAYER via2 ;
        RECT 1183.670 2796.360 1183.950 2796.640 ;
        RECT 2304.230 321.160 2304.510 321.440 ;
        RECT 1741.650 319.800 1741.930 320.080 ;
        RECT 2236.150 319.800 2236.430 320.080 ;
        RECT 1364.910 319.120 1365.190 319.400 ;
        RECT 1365.830 319.120 1366.110 319.400 ;
        RECT 1676.330 319.120 1676.610 319.400 ;
        RECT 1634.010 318.440 1634.290 318.720 ;
        RECT 1741.650 318.440 1741.930 318.720 ;
        RECT 1797.770 318.440 1798.050 318.720 ;
        RECT 1992.350 318.440 1992.630 318.720 ;
        RECT 1995.110 318.440 1995.390 318.720 ;
        RECT 2089.410 318.440 2089.690 318.720 ;
        RECT 2098.150 318.440 2098.430 318.720 ;
        RECT 2235.690 318.440 2235.970 318.720 ;
        RECT 2304.230 319.120 2304.510 319.400 ;
        RECT 1828.130 317.760 1828.410 318.040 ;
      LAYER met3 ;
        RECT 1183.645 2796.650 1183.975 2796.665 ;
        RECT 1186.150 2796.650 1186.530 2796.660 ;
        RECT 1183.645 2796.350 1186.530 2796.650 ;
        RECT 1183.645 2796.335 1183.975 2796.350 ;
        RECT 1186.150 2796.340 1186.530 2796.350 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2916.710 322.510 2924.800 322.810 ;
        RECT 2269.910 321.450 2270.290 321.460 ;
        RECT 2304.205 321.450 2304.535 321.465 ;
        RECT 2269.910 321.150 2304.535 321.450 ;
        RECT 2269.910 321.140 2270.290 321.150 ;
        RECT 2304.205 321.135 2304.535 321.150 ;
        RECT 1717.910 320.090 1718.290 320.100 ;
        RECT 1741.625 320.090 1741.955 320.105 ;
        RECT 2236.125 320.090 2236.455 320.105 ;
        RECT 2269.910 320.090 2270.290 320.100 ;
        RECT 1717.910 319.790 1741.955 320.090 ;
        RECT 1717.910 319.780 1718.290 319.790 ;
        RECT 1741.625 319.775 1741.955 319.790 ;
        RECT 1883.550 319.790 1931.690 320.090 ;
        RECT 1364.885 319.410 1365.215 319.425 ;
        RECT 1268.990 319.110 1365.215 319.410 ;
        RECT 1186.150 318.050 1186.530 318.060 ;
        RECT 1268.990 318.050 1269.290 319.110 ;
        RECT 1364.885 319.095 1365.215 319.110 ;
        RECT 1365.805 319.410 1366.135 319.425 ;
        RECT 1676.305 319.410 1676.635 319.425 ;
        RECT 1365.805 319.110 1372.330 319.410 ;
        RECT 1365.805 319.095 1366.135 319.110 ;
        RECT 1372.030 318.730 1372.330 319.110 ;
        RECT 1448.390 319.110 1463.410 319.410 ;
        RECT 1448.390 318.730 1448.690 319.110 ;
        RECT 1372.030 318.430 1448.690 318.730 ;
        RECT 1463.110 318.730 1463.410 319.110 ;
        RECT 1676.305 319.110 1684.210 319.410 ;
        RECT 1676.305 319.095 1676.635 319.110 ;
        RECT 1633.985 318.730 1634.315 318.745 ;
        RECT 1463.110 318.430 1587.610 318.730 ;
        RECT 1186.150 317.750 1269.290 318.050 ;
        RECT 1587.310 318.050 1587.610 318.430 ;
        RECT 1628.710 318.430 1634.315 318.730 ;
        RECT 1683.910 318.730 1684.210 319.110 ;
        RECT 1717.910 318.730 1718.290 318.740 ;
        RECT 1683.910 318.430 1718.290 318.730 ;
        RECT 1628.710 318.050 1629.010 318.430 ;
        RECT 1633.985 318.415 1634.315 318.430 ;
        RECT 1717.910 318.420 1718.290 318.430 ;
        RECT 1741.625 318.730 1741.955 318.745 ;
        RECT 1797.745 318.730 1798.075 318.745 ;
        RECT 1883.550 318.730 1883.850 319.790 ;
        RECT 1741.625 318.430 1798.075 318.730 ;
        RECT 1741.625 318.415 1741.955 318.430 ;
        RECT 1797.745 318.415 1798.075 318.430 ;
        RECT 1849.510 318.430 1883.850 318.730 ;
        RECT 1587.310 317.750 1629.010 318.050 ;
        RECT 1828.105 318.050 1828.435 318.065 ;
        RECT 1849.510 318.050 1849.810 318.430 ;
        RECT 1828.105 317.750 1849.810 318.050 ;
        RECT 1931.390 318.050 1931.690 319.790 ;
        RECT 2236.125 319.790 2270.290 320.090 ;
        RECT 2236.125 319.775 2236.455 319.790 ;
        RECT 2269.910 319.780 2270.290 319.790 ;
        RECT 2304.205 319.410 2304.535 319.425 ;
        RECT 2304.205 319.110 2353.050 319.410 ;
        RECT 2304.205 319.095 2304.535 319.110 ;
        RECT 1992.325 318.730 1992.655 318.745 ;
        RECT 1946.110 318.430 1992.655 318.730 ;
        RECT 1946.110 318.050 1946.410 318.430 ;
        RECT 1992.325 318.415 1992.655 318.430 ;
        RECT 1995.085 318.730 1995.415 318.745 ;
        RECT 2089.385 318.730 2089.715 318.745 ;
        RECT 1995.085 318.430 2028.290 318.730 ;
        RECT 1995.085 318.415 1995.415 318.430 ;
        RECT 1931.390 317.750 1946.410 318.050 ;
        RECT 2027.990 318.050 2028.290 318.430 ;
        RECT 2042.710 318.430 2089.715 318.730 ;
        RECT 2042.710 318.050 2043.010 318.430 ;
        RECT 2089.385 318.415 2089.715 318.430 ;
        RECT 2098.125 318.730 2098.455 318.745 ;
        RECT 2235.665 318.730 2235.995 318.745 ;
        RECT 2098.125 318.430 2124.890 318.730 ;
        RECT 2098.125 318.415 2098.455 318.430 ;
        RECT 2027.990 317.750 2043.010 318.050 ;
        RECT 2124.590 318.050 2124.890 318.430 ;
        RECT 2139.310 318.430 2235.995 318.730 ;
        RECT 2352.750 318.730 2353.050 319.110 ;
        RECT 2401.510 319.110 2449.650 319.410 ;
        RECT 2352.750 318.430 2400.890 318.730 ;
        RECT 2139.310 318.050 2139.610 318.430 ;
        RECT 2235.665 318.415 2235.995 318.430 ;
        RECT 2124.590 317.750 2139.610 318.050 ;
        RECT 2400.590 318.050 2400.890 318.430 ;
        RECT 2401.510 318.050 2401.810 319.110 ;
        RECT 2449.350 318.730 2449.650 319.110 ;
        RECT 2498.110 319.110 2546.250 319.410 ;
        RECT 2449.350 318.430 2497.490 318.730 ;
        RECT 2400.590 317.750 2401.810 318.050 ;
        RECT 2497.190 318.050 2497.490 318.430 ;
        RECT 2498.110 318.050 2498.410 319.110 ;
        RECT 2545.950 318.730 2546.250 319.110 ;
        RECT 2594.710 319.110 2642.850 319.410 ;
        RECT 2545.950 318.430 2594.090 318.730 ;
        RECT 2497.190 317.750 2498.410 318.050 ;
        RECT 2593.790 318.050 2594.090 318.430 ;
        RECT 2594.710 318.050 2595.010 319.110 ;
        RECT 2642.550 318.730 2642.850 319.110 ;
        RECT 2691.310 319.110 2739.450 319.410 ;
        RECT 2642.550 318.430 2690.690 318.730 ;
        RECT 2593.790 317.750 2595.010 318.050 ;
        RECT 2690.390 318.050 2690.690 318.430 ;
        RECT 2691.310 318.050 2691.610 319.110 ;
        RECT 2739.150 318.730 2739.450 319.110 ;
        RECT 2787.910 319.110 2836.050 319.410 ;
        RECT 2739.150 318.430 2787.290 318.730 ;
        RECT 2690.390 317.750 2691.610 318.050 ;
        RECT 2786.990 318.050 2787.290 318.430 ;
        RECT 2787.910 318.050 2788.210 319.110 ;
        RECT 2835.750 318.730 2836.050 319.110 ;
        RECT 2916.710 318.730 2917.010 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2835.750 318.430 2883.890 318.730 ;
        RECT 2786.990 317.750 2788.210 318.050 ;
        RECT 2883.590 318.050 2883.890 318.430 ;
        RECT 2884.510 318.430 2917.010 318.730 ;
        RECT 2884.510 318.050 2884.810 318.430 ;
        RECT 2883.590 317.750 2884.810 318.050 ;
        RECT 1186.150 317.740 1186.530 317.750 ;
        RECT 1828.105 317.735 1828.435 317.750 ;
      LAYER via3 ;
        RECT 1186.180 2796.340 1186.500 2796.660 ;
        RECT 2269.940 321.140 2270.260 321.460 ;
        RECT 1717.940 319.780 1718.260 320.100 ;
        RECT 1186.180 317.740 1186.500 318.060 ;
        RECT 1717.940 318.420 1718.260 318.740 ;
        RECT 2269.940 319.780 2270.260 320.100 ;
      LAYER met4 ;
        RECT 1186.175 2796.335 1186.505 2796.665 ;
        RECT 1186.190 318.065 1186.490 2796.335 ;
        RECT 2269.935 321.135 2270.265 321.465 ;
        RECT 2269.950 320.105 2270.250 321.135 ;
        RECT 1717.935 319.775 1718.265 320.105 ;
        RECT 2269.935 319.775 2270.265 320.105 ;
        RECT 1717.950 318.745 1718.250 319.775 ;
        RECT 1717.935 318.415 1718.265 318.745 ;
        RECT 1186.175 317.735 1186.505 318.065 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3500.200 1176.150 3500.260 ;
        RECT 1731.970 3500.200 1732.290 3500.260 ;
        RECT 1175.830 3500.060 1732.290 3500.200 ;
        RECT 1175.830 3500.000 1176.150 3500.060 ;
        RECT 1731.970 3500.000 1732.290 3500.060 ;
      LAYER via ;
        RECT 1175.860 3500.000 1176.120 3500.260 ;
        RECT 1732.000 3500.000 1732.260 3500.260 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3500.290 1176.060 3517.600 ;
        RECT 1175.860 3499.970 1176.120 3500.290 ;
        RECT 1732.000 3499.970 1732.260 3500.290 ;
        RECT 1732.060 2799.970 1732.200 3499.970 ;
        RECT 1732.385 2799.970 1732.665 2800.000 ;
        RECT 1732.060 2799.830 1732.665 2799.970 ;
        RECT 1732.385 2796.000 1732.665 2799.830 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3504.620 851.850 3504.680 ;
        RECT 1759.570 3504.620 1759.890 3504.680 ;
        RECT 851.530 3504.480 1759.890 3504.620 ;
        RECT 851.530 3504.420 851.850 3504.480 ;
        RECT 1759.570 3504.420 1759.890 3504.480 ;
      LAYER via ;
        RECT 851.560 3504.420 851.820 3504.680 ;
        RECT 1759.600 3504.420 1759.860 3504.680 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3504.710 851.760 3517.600 ;
        RECT 851.560 3504.390 851.820 3504.710 ;
        RECT 1759.600 3504.390 1759.860 3504.710 ;
        RECT 1759.660 2799.970 1759.800 3504.390 ;
        RECT 1761.365 2799.970 1761.645 2800.000 ;
        RECT 1759.660 2799.830 1761.645 2799.970 ;
        RECT 1761.365 2796.000 1761.645 2799.830 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3502.920 527.550 3502.980 ;
        RECT 1787.170 3502.920 1787.490 3502.980 ;
        RECT 527.230 3502.780 1787.490 3502.920 ;
        RECT 527.230 3502.720 527.550 3502.780 ;
        RECT 1787.170 3502.720 1787.490 3502.780 ;
      LAYER via ;
        RECT 527.260 3502.720 527.520 3502.980 ;
        RECT 1787.200 3502.720 1787.460 3502.980 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.010 527.460 3517.600 ;
        RECT 527.260 3502.690 527.520 3503.010 ;
        RECT 1787.200 3502.690 1787.460 3503.010 ;
        RECT 1787.260 2800.650 1787.400 3502.690 ;
        RECT 1787.260 2800.510 1788.780 2800.650 ;
        RECT 1788.640 2799.970 1788.780 2800.510 ;
        RECT 1790.345 2799.970 1790.625 2800.000 ;
        RECT 1788.640 2799.830 1790.625 2799.970 ;
        RECT 1790.345 2796.000 1790.625 2799.830 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 1814.770 3501.900 1815.090 3501.960 ;
        RECT 202.470 3501.760 1815.090 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 1814.770 3501.700 1815.090 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 1814.800 3501.700 1815.060 3501.960 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 1814.800 3501.670 1815.060 3501.990 ;
        RECT 1814.860 2801.330 1815.000 3501.670 ;
        RECT 1814.860 2801.190 1817.760 2801.330 ;
        RECT 1817.620 2799.970 1817.760 2801.190 ;
        RECT 1819.325 2799.970 1819.605 2800.000 ;
        RECT 1817.620 2799.830 1819.605 2799.970 ;
        RECT 1819.325 2796.000 1819.605 2799.830 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1842.370 3408.740 1842.690 3408.800 ;
        RECT 17.550 3408.600 1842.690 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1842.370 3408.540 1842.690 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1842.400 3408.540 1842.660 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1842.400 3408.510 1842.660 3408.830 ;
        RECT 1842.460 2801.330 1842.600 3408.510 ;
        RECT 1842.460 2801.190 1846.280 2801.330 ;
        RECT 1846.140 2799.970 1846.280 2801.190 ;
        RECT 1848.305 2799.970 1848.585 2800.000 ;
        RECT 1846.140 2799.830 1848.585 2799.970 ;
        RECT 1848.305 2796.000 1848.585 2799.830 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 1876.870 3119.060 1877.190 3119.120 ;
        RECT 17.090 3118.920 1877.190 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 1876.870 3118.860 1877.190 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 1876.900 3118.860 1877.160 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 1876.900 3118.830 1877.160 3119.150 ;
        RECT 1876.960 2799.970 1877.100 3118.830 ;
        RECT 1877.285 2799.970 1877.565 2800.000 ;
        RECT 1876.960 2799.830 1877.565 2799.970 ;
        RECT 1877.285 2796.000 1877.565 2799.830 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 1904.470 2836.180 1904.790 2836.240 ;
        RECT 17.090 2836.040 1904.790 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
        RECT 1904.470 2835.980 1904.790 2836.040 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
        RECT 1904.500 2835.980 1904.760 2836.240 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
        RECT 1904.500 2835.950 1904.760 2836.270 ;
        RECT 1904.560 2799.970 1904.700 2835.950 ;
        RECT 1905.805 2799.970 1906.085 2800.000 ;
        RECT 1904.560 2799.830 1906.085 2799.970 ;
        RECT 1905.805 2796.000 1906.085 2799.830 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 2811.700 15.570 2811.760 ;
        RECT 1934.830 2811.700 1935.150 2811.760 ;
        RECT 15.250 2811.560 1935.150 2811.700 ;
        RECT 15.250 2811.500 15.570 2811.560 ;
        RECT 1934.830 2811.500 1935.150 2811.560 ;
      LAYER via ;
        RECT 15.280 2811.500 15.540 2811.760 ;
        RECT 1934.860 2811.500 1935.120 2811.760 ;
      LAYER met2 ;
        RECT 15.280 2811.470 15.540 2811.790 ;
        RECT 1934.860 2811.470 1935.120 2811.790 ;
        RECT 15.340 2549.845 15.480 2811.470 ;
        RECT 1934.920 2800.000 1935.060 2811.470 ;
        RECT 1934.785 2796.000 1935.065 2800.000 ;
        RECT 15.270 2549.475 15.550 2549.845 ;
      LAYER via2 ;
        RECT 15.270 2549.520 15.550 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 15.245 2549.810 15.575 2549.825 ;
        RECT -4.800 2549.510 15.575 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 15.245 2549.495 15.575 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 2811.020 16.030 2811.080 ;
        RECT 1963.810 2811.020 1964.130 2811.080 ;
        RECT 15.710 2810.880 1964.130 2811.020 ;
        RECT 15.710 2810.820 16.030 2810.880 ;
        RECT 1963.810 2810.820 1964.130 2810.880 ;
      LAYER via ;
        RECT 15.740 2810.820 16.000 2811.080 ;
        RECT 1963.840 2810.820 1964.100 2811.080 ;
      LAYER met2 ;
        RECT 15.740 2810.790 16.000 2811.110 ;
        RECT 1963.840 2810.790 1964.100 2811.110 ;
        RECT 15.800 2262.205 15.940 2810.790 ;
        RECT 1963.900 2800.000 1964.040 2810.790 ;
        RECT 1963.765 2796.000 1964.045 2800.000 ;
        RECT 15.730 2261.835 16.010 2262.205 ;
      LAYER via2 ;
        RECT 15.730 2261.880 16.010 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 15.705 2262.170 16.035 2262.185 ;
        RECT -4.800 2261.870 16.035 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 15.705 2261.855 16.035 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2810.000 16.490 2810.060 ;
        RECT 1992.790 2810.000 1993.110 2810.060 ;
        RECT 16.170 2809.860 1993.110 2810.000 ;
        RECT 16.170 2809.800 16.490 2809.860 ;
        RECT 1992.790 2809.800 1993.110 2809.860 ;
      LAYER via ;
        RECT 16.200 2809.800 16.460 2810.060 ;
        RECT 1992.820 2809.800 1993.080 2810.060 ;
      LAYER met2 ;
        RECT 16.200 2809.770 16.460 2810.090 ;
        RECT 1992.820 2809.770 1993.080 2810.090 ;
        RECT 16.260 1975.245 16.400 2809.770 ;
        RECT 1992.880 2800.000 1993.020 2809.770 ;
        RECT 1992.745 2796.000 1993.025 2800.000 ;
        RECT 16.190 1974.875 16.470 1975.245 ;
      LAYER via2 ;
        RECT 16.190 1974.920 16.470 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 16.165 1975.210 16.495 1975.225 ;
        RECT -4.800 1974.910 16.495 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 16.165 1974.895 16.495 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1211.270 2812.635 1211.550 2813.005 ;
        RECT 1211.340 2800.000 1211.480 2812.635 ;
        RECT 2901.770 2811.955 2902.050 2812.325 ;
        RECT 1211.205 2796.000 1211.485 2800.000 ;
        RECT 2901.840 557.445 2901.980 2811.955 ;
        RECT 2901.770 557.075 2902.050 557.445 ;
      LAYER via2 ;
        RECT 1211.270 2812.680 1211.550 2812.960 ;
        RECT 2901.770 2812.000 2902.050 2812.280 ;
        RECT 2901.770 557.120 2902.050 557.400 ;
      LAYER met3 ;
        RECT 1211.245 2812.970 1211.575 2812.985 ;
        RECT 1211.245 2812.670 1220.530 2812.970 ;
        RECT 1211.245 2812.655 1211.575 2812.670 ;
        RECT 1220.230 2812.290 1220.530 2812.670 ;
        RECT 2901.745 2812.290 2902.075 2812.305 ;
        RECT 1220.230 2811.990 2902.075 2812.290 ;
        RECT 2901.745 2811.975 2902.075 2811.990 ;
        RECT 2901.745 557.410 2902.075 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2901.745 557.110 2924.800 557.410 ;
        RECT 2901.745 557.095 2902.075 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2021.790 2813.995 2022.070 2814.365 ;
        RECT 2021.860 2800.000 2022.000 2813.995 ;
        RECT 2021.725 2796.000 2022.005 2800.000 ;
      LAYER via2 ;
        RECT 2021.790 2814.040 2022.070 2814.320 ;
      LAYER met3 ;
        RECT 1184.310 2814.330 1184.690 2814.340 ;
        RECT 2021.765 2814.330 2022.095 2814.345 ;
        RECT 1184.310 2814.030 2022.095 2814.330 ;
        RECT 1184.310 2814.020 1184.690 2814.030 ;
        RECT 2021.765 2814.015 2022.095 2814.030 ;
        RECT 1184.310 1690.290 1184.690 1690.300 ;
        RECT 3.070 1689.990 1184.690 1690.290 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 3.070 1687.570 3.370 1689.990 ;
        RECT 1184.310 1689.980 1184.690 1689.990 ;
        RECT -4.800 1687.270 3.370 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
      LAYER via3 ;
        RECT 1184.340 2814.020 1184.660 2814.340 ;
        RECT 1184.340 1689.980 1184.660 1690.300 ;
      LAYER met4 ;
        RECT 1184.335 2814.015 1184.665 2814.345 ;
        RECT 1184.350 1690.305 1184.650 2814.015 ;
        RECT 1184.335 1689.975 1184.665 1690.305 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1860.845 2802.705 1861.935 2802.875 ;
        RECT 2001.605 2802.705 2002.695 2802.875 ;
      LAYER mcon ;
        RECT 1861.765 2802.705 1861.935 2802.875 ;
        RECT 2002.525 2802.705 2002.695 2802.875 ;
      LAYER met1 ;
        RECT 26.290 2802.860 26.610 2802.920 ;
        RECT 1860.785 2802.860 1861.075 2802.905 ;
        RECT 26.290 2802.720 1861.075 2802.860 ;
        RECT 26.290 2802.660 26.610 2802.720 ;
        RECT 1860.785 2802.675 1861.075 2802.720 ;
        RECT 1861.705 2802.860 1861.995 2802.905 ;
        RECT 2001.545 2802.860 2001.835 2802.905 ;
        RECT 1861.705 2802.720 2001.835 2802.860 ;
        RECT 1861.705 2802.675 1861.995 2802.720 ;
        RECT 2001.545 2802.675 2001.835 2802.720 ;
        RECT 2002.465 2802.860 2002.755 2802.905 ;
        RECT 2050.750 2802.860 2051.070 2802.920 ;
        RECT 2002.465 2802.720 2051.070 2802.860 ;
        RECT 2002.465 2802.675 2002.755 2802.720 ;
        RECT 2050.750 2802.660 2051.070 2802.720 ;
        RECT 13.870 1476.180 14.190 1476.240 ;
        RECT 26.290 1476.180 26.610 1476.240 ;
        RECT 13.870 1476.040 26.610 1476.180 ;
        RECT 13.870 1475.980 14.190 1476.040 ;
        RECT 26.290 1475.980 26.610 1476.040 ;
      LAYER via ;
        RECT 26.320 2802.660 26.580 2802.920 ;
        RECT 2050.780 2802.660 2051.040 2802.920 ;
        RECT 13.900 1475.980 14.160 1476.240 ;
        RECT 26.320 1475.980 26.580 1476.240 ;
      LAYER met2 ;
        RECT 26.320 2802.630 26.580 2802.950 ;
        RECT 2050.780 2802.630 2051.040 2802.950 ;
        RECT 26.380 1476.270 26.520 2802.630 ;
        RECT 2050.840 2800.000 2050.980 2802.630 ;
        RECT 2050.705 2796.000 2050.985 2800.000 ;
        RECT 13.900 1475.950 14.160 1476.270 ;
        RECT 26.320 1475.950 26.580 1476.270 ;
        RECT 13.960 1472.045 14.100 1475.950 ;
        RECT 13.890 1471.675 14.170 1472.045 ;
      LAYER via2 ;
        RECT 13.890 1471.720 14.170 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 13.865 1472.010 14.195 1472.025 ;
        RECT -4.800 1471.710 14.195 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 13.865 1471.695 14.195 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2079.750 2813.315 2080.030 2813.685 ;
        RECT 2079.820 2800.000 2079.960 2813.315 ;
        RECT 2079.685 2796.000 2079.965 2800.000 ;
        RECT 15.730 1262.235 16.010 1262.605 ;
        RECT 15.800 1256.485 15.940 1262.235 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
      LAYER via2 ;
        RECT 2079.750 2813.360 2080.030 2813.640 ;
        RECT 15.730 1262.280 16.010 1262.560 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
        RECT 1182.470 2813.650 1182.850 2813.660 ;
        RECT 2079.725 2813.650 2080.055 2813.665 ;
        RECT 1182.470 2813.350 2080.055 2813.650 ;
        RECT 1182.470 2813.340 1182.850 2813.350 ;
        RECT 2079.725 2813.335 2080.055 2813.350 ;
        RECT 15.705 1262.570 16.035 1262.585 ;
        RECT 1182.470 1262.570 1182.850 1262.580 ;
        RECT 15.705 1262.270 1182.850 1262.570 ;
        RECT 15.705 1262.255 16.035 1262.270 ;
        RECT 1182.470 1262.260 1182.850 1262.270 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
      LAYER via3 ;
        RECT 1182.500 2813.340 1182.820 2813.660 ;
        RECT 1182.500 1262.260 1182.820 1262.580 ;
      LAYER met4 ;
        RECT 1182.495 2813.335 1182.825 2813.665 ;
        RECT 1182.510 1262.585 1182.810 2813.335 ;
        RECT 1182.495 1262.255 1182.825 1262.585 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1861.305 2802.365 1862.395 2802.535 ;
        RECT 2001.145 2802.365 2002.235 2802.535 ;
      LAYER mcon ;
        RECT 1862.225 2802.365 1862.395 2802.535 ;
        RECT 2002.065 2802.365 2002.235 2802.535 ;
      LAYER met1 ;
        RECT 25.830 2802.520 26.150 2802.580 ;
        RECT 1861.245 2802.520 1861.535 2802.565 ;
        RECT 25.830 2802.380 1861.535 2802.520 ;
        RECT 25.830 2802.320 26.150 2802.380 ;
        RECT 1861.245 2802.335 1861.535 2802.380 ;
        RECT 1862.165 2802.520 1862.455 2802.565 ;
        RECT 2001.085 2802.520 2001.375 2802.565 ;
        RECT 1862.165 2802.380 2001.375 2802.520 ;
        RECT 1862.165 2802.335 1862.455 2802.380 ;
        RECT 2001.085 2802.335 2001.375 2802.380 ;
        RECT 2002.005 2802.520 2002.295 2802.565 ;
        RECT 2108.710 2802.520 2109.030 2802.580 ;
        RECT 2002.005 2802.380 2109.030 2802.520 ;
        RECT 2002.005 2802.335 2002.295 2802.380 ;
        RECT 2108.710 2802.320 2109.030 2802.380 ;
        RECT 13.870 1040.980 14.190 1041.040 ;
        RECT 25.830 1040.980 26.150 1041.040 ;
        RECT 13.870 1040.840 26.150 1040.980 ;
        RECT 13.870 1040.780 14.190 1040.840 ;
        RECT 25.830 1040.780 26.150 1040.840 ;
      LAYER via ;
        RECT 25.860 2802.320 26.120 2802.580 ;
        RECT 2108.740 2802.320 2109.000 2802.580 ;
        RECT 13.900 1040.780 14.160 1041.040 ;
        RECT 25.860 1040.780 26.120 1041.040 ;
      LAYER met2 ;
        RECT 25.860 2802.290 26.120 2802.610 ;
        RECT 2108.740 2802.290 2109.000 2802.610 ;
        RECT 25.920 1041.070 26.060 2802.290 ;
        RECT 2108.800 2800.000 2108.940 2802.290 ;
        RECT 2108.665 2796.000 2108.945 2800.000 ;
        RECT 13.900 1040.925 14.160 1041.070 ;
        RECT 13.890 1040.555 14.170 1040.925 ;
        RECT 25.860 1040.750 26.120 1041.070 ;
      LAYER via2 ;
        RECT 13.890 1040.600 14.170 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 13.865 1040.890 14.195 1040.905 ;
        RECT -4.800 1040.590 14.195 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 13.865 1040.575 14.195 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1861.765 2802.025 1862.855 2802.195 ;
        RECT 2001.605 2802.025 2002.695 2802.195 ;
      LAYER mcon ;
        RECT 1862.685 2802.025 1862.855 2802.195 ;
        RECT 2002.525 2802.025 2002.695 2802.195 ;
      LAYER met1 ;
        RECT 24.910 2802.180 25.230 2802.240 ;
        RECT 1861.705 2802.180 1861.995 2802.225 ;
        RECT 24.910 2802.040 1861.995 2802.180 ;
        RECT 24.910 2801.980 25.230 2802.040 ;
        RECT 1861.705 2801.995 1861.995 2802.040 ;
        RECT 1862.625 2802.180 1862.915 2802.225 ;
        RECT 2001.545 2802.180 2001.835 2802.225 ;
        RECT 1862.625 2802.040 2001.835 2802.180 ;
        RECT 1862.625 2801.995 1862.915 2802.040 ;
        RECT 2001.545 2801.995 2001.835 2802.040 ;
        RECT 2002.465 2802.180 2002.755 2802.225 ;
        RECT 2137.690 2802.180 2138.010 2802.240 ;
        RECT 2002.465 2802.040 2138.010 2802.180 ;
        RECT 2002.465 2801.995 2002.755 2802.040 ;
        RECT 2137.690 2801.980 2138.010 2802.040 ;
        RECT 13.870 827.460 14.190 827.520 ;
        RECT 24.910 827.460 25.230 827.520 ;
        RECT 13.870 827.320 25.230 827.460 ;
        RECT 13.870 827.260 14.190 827.320 ;
        RECT 24.910 827.260 25.230 827.320 ;
      LAYER via ;
        RECT 24.940 2801.980 25.200 2802.240 ;
        RECT 2137.720 2801.980 2137.980 2802.240 ;
        RECT 13.900 827.260 14.160 827.520 ;
        RECT 24.940 827.260 25.200 827.520 ;
      LAYER met2 ;
        RECT 24.940 2801.950 25.200 2802.270 ;
        RECT 2137.720 2801.950 2137.980 2802.270 ;
        RECT 25.000 827.550 25.140 2801.950 ;
        RECT 2137.780 2800.000 2137.920 2801.950 ;
        RECT 2137.645 2796.000 2137.925 2800.000 ;
        RECT 13.900 827.230 14.160 827.550 ;
        RECT 24.940 827.230 25.200 827.550 ;
        RECT 13.960 825.365 14.100 827.230 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.800 825.030 14.195 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 2801.840 24.310 2801.900 ;
        RECT 2001.070 2801.840 2001.390 2801.900 ;
        RECT 23.990 2801.700 2001.390 2801.840 ;
        RECT 23.990 2801.640 24.310 2801.700 ;
        RECT 2001.070 2801.640 2001.390 2801.700 ;
        RECT 2002.910 2801.840 2003.230 2801.900 ;
        RECT 2166.670 2801.840 2166.990 2801.900 ;
        RECT 2002.910 2801.700 2166.990 2801.840 ;
        RECT 2002.910 2801.640 2003.230 2801.700 ;
        RECT 2166.670 2801.640 2166.990 2801.700 ;
        RECT 13.870 610.540 14.190 610.600 ;
        RECT 23.990 610.540 24.310 610.600 ;
        RECT 13.870 610.400 24.310 610.540 ;
        RECT 13.870 610.340 14.190 610.400 ;
        RECT 23.990 610.340 24.310 610.400 ;
      LAYER via ;
        RECT 24.020 2801.640 24.280 2801.900 ;
        RECT 2001.100 2801.640 2001.360 2801.900 ;
        RECT 2002.940 2801.640 2003.200 2801.900 ;
        RECT 2166.700 2801.640 2166.960 2801.900 ;
        RECT 13.900 610.340 14.160 610.600 ;
        RECT 24.020 610.340 24.280 610.600 ;
      LAYER met2 ;
        RECT 24.020 2801.610 24.280 2801.930 ;
        RECT 2001.090 2801.755 2001.370 2802.125 ;
        RECT 2002.930 2801.755 2003.210 2802.125 ;
        RECT 2001.100 2801.610 2001.360 2801.755 ;
        RECT 2002.940 2801.610 2003.200 2801.755 ;
        RECT 2166.700 2801.610 2166.960 2801.930 ;
        RECT 24.080 610.630 24.220 2801.610 ;
        RECT 2166.760 2800.000 2166.900 2801.610 ;
        RECT 2166.625 2796.000 2166.905 2800.000 ;
        RECT 13.900 610.485 14.160 610.630 ;
        RECT 13.890 610.115 14.170 610.485 ;
        RECT 24.020 610.310 24.280 610.630 ;
      LAYER via2 ;
        RECT 2001.090 2801.800 2001.370 2802.080 ;
        RECT 2002.930 2801.800 2003.210 2802.080 ;
        RECT 13.890 610.160 14.170 610.440 ;
      LAYER met3 ;
        RECT 2001.065 2802.090 2001.395 2802.105 ;
        RECT 2002.905 2802.090 2003.235 2802.105 ;
        RECT 2001.065 2801.790 2003.235 2802.090 ;
        RECT 2001.065 2801.775 2001.395 2801.790 ;
        RECT 2002.905 2801.775 2003.235 2801.790 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 13.865 610.450 14.195 610.465 ;
        RECT -4.800 610.150 14.195 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 13.865 610.135 14.195 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1861.765 2801.345 1862.855 2801.515 ;
        RECT 2001.605 2801.345 2002.695 2801.515 ;
      LAYER mcon ;
        RECT 1862.685 2801.345 1862.855 2801.515 ;
        RECT 2002.525 2801.345 2002.695 2801.515 ;
      LAYER met1 ;
        RECT 30.890 2801.500 31.210 2801.560 ;
        RECT 1861.705 2801.500 1861.995 2801.545 ;
        RECT 30.890 2801.360 1861.995 2801.500 ;
        RECT 30.890 2801.300 31.210 2801.360 ;
        RECT 1861.705 2801.315 1861.995 2801.360 ;
        RECT 1862.625 2801.500 1862.915 2801.545 ;
        RECT 2001.545 2801.500 2001.835 2801.545 ;
        RECT 1862.625 2801.360 2001.835 2801.500 ;
        RECT 1862.625 2801.315 1862.915 2801.360 ;
        RECT 2001.545 2801.315 2001.835 2801.360 ;
        RECT 2002.465 2801.500 2002.755 2801.545 ;
        RECT 2195.650 2801.500 2195.970 2801.560 ;
        RECT 2002.465 2801.360 2195.970 2801.500 ;
        RECT 2002.465 2801.315 2002.755 2801.360 ;
        RECT 2195.650 2801.300 2195.970 2801.360 ;
        RECT 13.870 397.360 14.190 397.420 ;
        RECT 30.890 397.360 31.210 397.420 ;
        RECT 13.870 397.220 31.210 397.360 ;
        RECT 13.870 397.160 14.190 397.220 ;
        RECT 30.890 397.160 31.210 397.220 ;
      LAYER via ;
        RECT 30.920 2801.300 31.180 2801.560 ;
        RECT 2195.680 2801.300 2195.940 2801.560 ;
        RECT 13.900 397.160 14.160 397.420 ;
        RECT 30.920 397.160 31.180 397.420 ;
      LAYER met2 ;
        RECT 30.920 2801.270 31.180 2801.590 ;
        RECT 2195.680 2801.270 2195.940 2801.590 ;
        RECT 30.980 397.450 31.120 2801.270 ;
        RECT 2195.740 2800.000 2195.880 2801.270 ;
        RECT 2195.605 2796.000 2195.885 2800.000 ;
        RECT 13.900 397.130 14.160 397.450 ;
        RECT 30.920 397.130 31.180 397.450 ;
        RECT 13.960 394.925 14.100 397.130 ;
        RECT 13.890 394.555 14.170 394.925 ;
      LAYER via2 ;
        RECT 13.890 394.600 14.170 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 13.865 394.890 14.195 394.905 ;
        RECT -4.800 394.590 14.195 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 13.865 394.575 14.195 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2222.810 2796.570 2223.090 2796.685 ;
        RECT 2224.585 2796.570 2224.865 2800.000 ;
        RECT 2222.810 2796.430 2224.865 2796.570 ;
        RECT 2222.810 2796.315 2223.090 2796.430 ;
        RECT 2224.585 2796.000 2224.865 2796.430 ;
      LAYER via2 ;
        RECT 2222.810 2796.360 2223.090 2796.640 ;
      LAYER met3 ;
        RECT 2222.070 2796.650 2222.450 2796.660 ;
        RECT 2222.785 2796.650 2223.115 2796.665 ;
        RECT 2222.070 2796.350 2223.115 2796.650 ;
        RECT 2222.070 2796.340 2222.450 2796.350 ;
        RECT 2222.785 2796.335 2223.115 2796.350 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 2222.070 179.330 2222.450 179.340 ;
        RECT -4.800 179.030 2222.450 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 2222.070 179.020 2222.450 179.030 ;
      LAYER via3 ;
        RECT 2222.100 2796.340 2222.420 2796.660 ;
        RECT 2222.100 179.020 2222.420 179.340 ;
      LAYER met4 ;
        RECT 2222.095 2796.335 2222.425 2796.665 ;
        RECT 2222.110 179.345 2222.410 2796.335 ;
        RECT 2222.095 179.015 2222.425 179.345 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1240.250 2812.635 1240.530 2813.005 ;
        RECT 2902.690 2812.635 2902.970 2813.005 ;
        RECT 1240.320 2800.000 1240.460 2812.635 ;
        RECT 1240.185 2796.000 1240.465 2800.000 ;
        RECT 2902.760 792.045 2902.900 2812.635 ;
        RECT 2902.690 791.675 2902.970 792.045 ;
      LAYER via2 ;
        RECT 1240.250 2812.680 1240.530 2812.960 ;
        RECT 2902.690 2812.680 2902.970 2812.960 ;
        RECT 2902.690 791.720 2902.970 792.000 ;
      LAYER met3 ;
        RECT 1240.225 2812.970 1240.555 2812.985 ;
        RECT 2902.665 2812.970 2902.995 2812.985 ;
        RECT 1240.225 2812.670 2902.995 2812.970 ;
        RECT 1240.225 2812.655 1240.555 2812.670 ;
        RECT 2902.665 2812.655 2902.995 2812.670 ;
        RECT 2902.665 792.010 2902.995 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2902.665 791.710 2924.800 792.010 ;
        RECT 2902.665 791.695 2902.995 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2056.730 2802.860 2057.050 2802.920 ;
        RECT 2121.590 2802.860 2121.910 2802.920 ;
        RECT 2056.730 2802.720 2121.910 2802.860 ;
        RECT 2056.730 2802.660 2057.050 2802.720 ;
        RECT 2121.590 2802.660 2121.910 2802.720 ;
      LAYER via ;
        RECT 2056.760 2802.660 2057.020 2802.920 ;
        RECT 2121.620 2802.660 2121.880 2802.920 ;
      LAYER met2 ;
        RECT 1628.490 2804.475 1628.770 2804.845 ;
        RECT 1931.170 2804.475 1931.450 2804.845 ;
        RECT 1628.560 2803.485 1628.700 2804.475 ;
        RECT 1725.090 2803.795 1725.370 2804.165 ;
        RECT 1786.730 2803.795 1787.010 2804.165 ;
        RECT 1835.030 2803.795 1835.310 2804.165 ;
        RECT 1628.490 2803.115 1628.770 2803.485 ;
        RECT 1724.630 2803.115 1724.910 2803.485 ;
        RECT 1724.700 2802.690 1724.840 2803.115 ;
        RECT 1725.160 2802.690 1725.300 2803.795 ;
        RECT 1786.800 2802.805 1786.940 2803.795 ;
        RECT 1835.100 2802.805 1835.240 2803.795 ;
        RECT 1931.240 2802.805 1931.380 2804.475 ;
        RECT 2121.610 2803.795 2121.890 2804.165 ;
        RECT 2159.330 2803.795 2159.610 2804.165 ;
        RECT 2121.680 2802.950 2121.820 2803.795 ;
        RECT 1724.700 2802.550 1725.300 2802.690 ;
        RECT 1786.730 2802.435 1787.010 2802.805 ;
        RECT 1835.030 2802.435 1835.310 2802.805 ;
        RECT 1931.170 2802.435 1931.450 2802.805 ;
        RECT 1932.090 2802.435 1932.370 2802.805 ;
        RECT 1994.650 2802.690 1994.930 2802.805 ;
        RECT 1993.800 2802.550 1994.930 2802.690 ;
        RECT 1269.230 2801.755 1269.510 2802.125 ;
        RECT 1932.160 2802.010 1932.300 2802.435 ;
        RECT 1993.800 2802.125 1993.940 2802.550 ;
        RECT 1994.650 2802.435 1994.930 2802.550 ;
        RECT 2028.690 2802.435 2028.970 2802.805 ;
        RECT 2056.760 2802.630 2057.020 2802.950 ;
        RECT 2121.620 2802.630 2121.880 2802.950 ;
        RECT 2159.400 2802.805 2159.540 2803.795 ;
        RECT 1932.550 2802.010 1932.830 2802.125 ;
        RECT 1932.160 2801.870 1932.830 2802.010 ;
        RECT 1932.550 2801.755 1932.830 2801.870 ;
        RECT 1979.010 2802.010 1979.290 2802.125 ;
        RECT 1979.930 2802.010 1980.210 2802.125 ;
        RECT 1979.010 2801.870 1980.210 2802.010 ;
        RECT 1979.010 2801.755 1979.290 2801.870 ;
        RECT 1979.930 2801.755 1980.210 2801.870 ;
        RECT 1993.730 2801.755 1994.010 2802.125 ;
        RECT 2028.760 2802.010 2028.900 2802.435 ;
        RECT 2029.150 2802.010 2029.430 2802.125 ;
        RECT 2028.760 2801.870 2029.430 2802.010 ;
        RECT 2029.150 2801.755 2029.430 2801.870 ;
        RECT 2056.290 2801.755 2056.570 2802.125 ;
        RECT 1269.300 2800.000 1269.440 2801.755 ;
        RECT 2056.360 2801.330 2056.500 2801.755 ;
        RECT 2056.820 2801.330 2056.960 2802.630 ;
        RECT 2159.330 2802.435 2159.610 2802.805 ;
        RECT 2056.360 2801.190 2056.960 2801.330 ;
        RECT 1269.165 2796.000 1269.445 2800.000 ;
      LAYER via2 ;
        RECT 1628.490 2804.520 1628.770 2804.800 ;
        RECT 1931.170 2804.520 1931.450 2804.800 ;
        RECT 1725.090 2803.840 1725.370 2804.120 ;
        RECT 1786.730 2803.840 1787.010 2804.120 ;
        RECT 1835.030 2803.840 1835.310 2804.120 ;
        RECT 1628.490 2803.160 1628.770 2803.440 ;
        RECT 1724.630 2803.160 1724.910 2803.440 ;
        RECT 2121.610 2803.840 2121.890 2804.120 ;
        RECT 2159.330 2803.840 2159.610 2804.120 ;
        RECT 1786.730 2802.480 1787.010 2802.760 ;
        RECT 1835.030 2802.480 1835.310 2802.760 ;
        RECT 1931.170 2802.480 1931.450 2802.760 ;
        RECT 1932.090 2802.480 1932.370 2802.760 ;
        RECT 1269.230 2801.800 1269.510 2802.080 ;
        RECT 1994.650 2802.480 1994.930 2802.760 ;
        RECT 2028.690 2802.480 2028.970 2802.760 ;
        RECT 1932.550 2801.800 1932.830 2802.080 ;
        RECT 1979.010 2801.800 1979.290 2802.080 ;
        RECT 1979.930 2801.800 1980.210 2802.080 ;
        RECT 1993.730 2801.800 1994.010 2802.080 ;
        RECT 2029.150 2801.800 2029.430 2802.080 ;
        RECT 2056.290 2801.800 2056.570 2802.080 ;
        RECT 2159.330 2802.480 2159.610 2802.760 ;
      LAYER met3 ;
        RECT 1628.465 2804.810 1628.795 2804.825 ;
        RECT 1675.590 2804.810 1675.970 2804.820 ;
        RECT 1628.465 2804.510 1675.970 2804.810 ;
        RECT 1628.465 2804.495 1628.795 2804.510 ;
        RECT 1675.590 2804.500 1675.970 2804.510 ;
        RECT 1883.510 2804.810 1883.890 2804.820 ;
        RECT 1931.145 2804.810 1931.475 2804.825 ;
        RECT 1883.510 2804.510 1931.475 2804.810 ;
        RECT 1883.510 2804.500 1883.890 2804.510 ;
        RECT 1931.145 2804.495 1931.475 2804.510 ;
        RECT 1400.510 2804.130 1400.890 2804.140 ;
        RECT 1725.065 2804.130 1725.395 2804.145 ;
        RECT 1786.705 2804.140 1787.035 2804.145 ;
        RECT 1786.705 2804.130 1787.290 2804.140 ;
        RECT 1835.005 2804.130 1835.335 2804.145 ;
        RECT 1400.510 2803.830 1466.170 2804.130 ;
        RECT 1400.510 2803.820 1400.890 2803.830 ;
        RECT 1400.510 2802.770 1400.890 2802.780 ;
        RECT 1321.430 2802.470 1400.890 2802.770 ;
        RECT 1465.870 2802.770 1466.170 2803.830 ;
        RECT 1497.150 2803.830 1545.290 2804.130 ;
        RECT 1497.150 2802.770 1497.450 2803.830 ;
        RECT 1544.990 2802.780 1545.290 2803.830 ;
        RECT 1725.065 2803.830 1835.335 2804.130 ;
        RECT 1725.065 2803.815 1725.395 2803.830 ;
        RECT 1786.705 2803.820 1787.290 2803.830 ;
        RECT 1786.705 2803.815 1787.035 2803.820 ;
        RECT 1835.005 2803.815 1835.335 2803.830 ;
        RECT 2121.585 2804.130 2121.915 2804.145 ;
        RECT 2159.305 2804.130 2159.635 2804.145 ;
        RECT 2121.585 2803.830 2159.635 2804.130 ;
        RECT 2121.585 2803.815 2121.915 2803.830 ;
        RECT 2159.305 2803.815 2159.635 2803.830 ;
        RECT 1628.465 2803.450 1628.795 2803.465 ;
        RECT 1593.750 2803.150 1628.795 2803.450 ;
        RECT 1465.870 2802.470 1497.450 2802.770 ;
        RECT 1269.205 2802.090 1269.535 2802.105 ;
        RECT 1321.430 2802.090 1321.730 2802.470 ;
        RECT 1400.510 2802.460 1400.890 2802.470 ;
        RECT 1544.950 2802.460 1545.330 2802.780 ;
        RECT 1269.205 2801.790 1321.730 2802.090 ;
        RECT 1544.950 2802.090 1545.330 2802.100 ;
        RECT 1593.750 2802.090 1594.050 2803.150 ;
        RECT 1628.465 2803.135 1628.795 2803.150 ;
        RECT 1676.510 2803.450 1676.890 2803.460 ;
        RECT 1724.605 2803.450 1724.935 2803.465 ;
        RECT 1676.510 2803.150 1724.935 2803.450 ;
        RECT 1676.510 2803.140 1676.890 2803.150 ;
        RECT 1724.605 2803.135 1724.935 2803.150 ;
        RECT 1786.705 2802.780 1787.035 2802.785 ;
        RECT 1786.705 2802.770 1787.290 2802.780 ;
        RECT 1835.005 2802.770 1835.335 2802.785 ;
        RECT 1883.510 2802.770 1883.890 2802.780 ;
        RECT 1786.705 2802.470 1787.670 2802.770 ;
        RECT 1835.005 2802.470 1883.890 2802.770 ;
        RECT 1786.705 2802.460 1787.290 2802.470 ;
        RECT 1786.705 2802.455 1787.035 2802.460 ;
        RECT 1835.005 2802.455 1835.335 2802.470 ;
        RECT 1883.510 2802.460 1883.890 2802.470 ;
        RECT 1931.145 2802.770 1931.475 2802.785 ;
        RECT 1932.065 2802.770 1932.395 2802.785 ;
        RECT 1931.145 2802.470 1932.395 2802.770 ;
        RECT 1931.145 2802.455 1931.475 2802.470 ;
        RECT 1932.065 2802.455 1932.395 2802.470 ;
        RECT 1994.625 2802.770 1994.955 2802.785 ;
        RECT 2028.665 2802.770 2028.995 2802.785 ;
        RECT 1994.625 2802.470 2028.995 2802.770 ;
        RECT 1994.625 2802.455 1994.955 2802.470 ;
        RECT 2028.665 2802.455 2028.995 2802.470 ;
        RECT 2159.305 2802.770 2159.635 2802.785 ;
        RECT 2159.305 2802.470 2208.610 2802.770 ;
        RECT 2159.305 2802.455 2159.635 2802.470 ;
        RECT 1544.950 2801.790 1594.050 2802.090 ;
        RECT 1932.525 2802.090 1932.855 2802.105 ;
        RECT 1978.985 2802.090 1979.315 2802.105 ;
        RECT 1932.525 2801.790 1979.315 2802.090 ;
        RECT 1269.205 2801.775 1269.535 2801.790 ;
        RECT 1544.950 2801.780 1545.330 2801.790 ;
        RECT 1932.525 2801.775 1932.855 2801.790 ;
        RECT 1978.985 2801.775 1979.315 2801.790 ;
        RECT 1979.905 2802.090 1980.235 2802.105 ;
        RECT 1993.705 2802.090 1994.035 2802.105 ;
        RECT 1979.905 2801.790 1994.035 2802.090 ;
        RECT 1979.905 2801.775 1980.235 2801.790 ;
        RECT 1993.705 2801.775 1994.035 2801.790 ;
        RECT 2029.125 2802.090 2029.455 2802.105 ;
        RECT 2056.265 2802.090 2056.595 2802.105 ;
        RECT 2029.125 2801.790 2056.595 2802.090 ;
        RECT 2029.125 2801.775 2029.455 2801.790 ;
        RECT 2056.265 2801.775 2056.595 2801.790 ;
        RECT 2208.310 2801.410 2208.610 2802.470 ;
        RECT 2238.630 2801.410 2239.010 2801.420 ;
        RECT 2208.310 2801.110 2239.010 2801.410 ;
        RECT 2238.630 2801.100 2239.010 2801.110 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2916.710 1026.310 2924.800 1026.610 ;
        RECT 2238.630 1023.210 2239.010 1023.220 ;
        RECT 2238.630 1022.910 2256.450 1023.210 ;
        RECT 2238.630 1022.900 2239.010 1022.910 ;
        RECT 2256.150 1022.530 2256.450 1022.910 ;
        RECT 2304.910 1022.910 2353.050 1023.210 ;
        RECT 2256.150 1022.230 2304.290 1022.530 ;
        RECT 2303.990 1021.850 2304.290 1022.230 ;
        RECT 2304.910 1021.850 2305.210 1022.910 ;
        RECT 2352.750 1022.530 2353.050 1022.910 ;
        RECT 2401.510 1022.910 2449.650 1023.210 ;
        RECT 2352.750 1022.230 2400.890 1022.530 ;
        RECT 2303.990 1021.550 2305.210 1021.850 ;
        RECT 2400.590 1021.850 2400.890 1022.230 ;
        RECT 2401.510 1021.850 2401.810 1022.910 ;
        RECT 2449.350 1022.530 2449.650 1022.910 ;
        RECT 2498.110 1022.910 2546.250 1023.210 ;
        RECT 2449.350 1022.230 2497.490 1022.530 ;
        RECT 2400.590 1021.550 2401.810 1021.850 ;
        RECT 2497.190 1021.850 2497.490 1022.230 ;
        RECT 2498.110 1021.850 2498.410 1022.910 ;
        RECT 2545.950 1022.530 2546.250 1022.910 ;
        RECT 2594.710 1022.910 2642.850 1023.210 ;
        RECT 2545.950 1022.230 2594.090 1022.530 ;
        RECT 2497.190 1021.550 2498.410 1021.850 ;
        RECT 2593.790 1021.850 2594.090 1022.230 ;
        RECT 2594.710 1021.850 2595.010 1022.910 ;
        RECT 2642.550 1022.530 2642.850 1022.910 ;
        RECT 2691.310 1022.910 2739.450 1023.210 ;
        RECT 2642.550 1022.230 2690.690 1022.530 ;
        RECT 2593.790 1021.550 2595.010 1021.850 ;
        RECT 2690.390 1021.850 2690.690 1022.230 ;
        RECT 2691.310 1021.850 2691.610 1022.910 ;
        RECT 2739.150 1022.530 2739.450 1022.910 ;
        RECT 2787.910 1022.910 2836.050 1023.210 ;
        RECT 2739.150 1022.230 2787.290 1022.530 ;
        RECT 2690.390 1021.550 2691.610 1021.850 ;
        RECT 2786.990 1021.850 2787.290 1022.230 ;
        RECT 2787.910 1021.850 2788.210 1022.910 ;
        RECT 2835.750 1022.530 2836.050 1022.910 ;
        RECT 2916.710 1022.530 2917.010 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2835.750 1022.230 2883.890 1022.530 ;
        RECT 2786.990 1021.550 2788.210 1021.850 ;
        RECT 2883.590 1021.850 2883.890 1022.230 ;
        RECT 2884.510 1022.230 2917.010 1022.530 ;
        RECT 2884.510 1021.850 2884.810 1022.230 ;
        RECT 2883.590 1021.550 2884.810 1021.850 ;
      LAYER via3 ;
        RECT 1675.620 2804.500 1675.940 2804.820 ;
        RECT 1883.540 2804.500 1883.860 2804.820 ;
        RECT 1400.540 2803.820 1400.860 2804.140 ;
        RECT 1400.540 2802.460 1400.860 2802.780 ;
        RECT 1786.940 2803.820 1787.260 2804.140 ;
        RECT 1544.980 2802.460 1545.300 2802.780 ;
        RECT 1544.980 2801.780 1545.300 2802.100 ;
        RECT 1676.540 2803.140 1676.860 2803.460 ;
        RECT 1786.940 2802.460 1787.260 2802.780 ;
        RECT 1883.540 2802.460 1883.860 2802.780 ;
        RECT 2238.660 2801.100 2238.980 2801.420 ;
        RECT 2238.660 1022.900 2238.980 1023.220 ;
      LAYER met4 ;
        RECT 1675.615 2804.495 1675.945 2804.825 ;
        RECT 1883.535 2804.495 1883.865 2804.825 ;
        RECT 1400.535 2803.815 1400.865 2804.145 ;
        RECT 1400.550 2802.785 1400.850 2803.815 ;
        RECT 1675.630 2803.450 1675.930 2804.495 ;
        RECT 1786.935 2803.815 1787.265 2804.145 ;
        RECT 1676.535 2803.450 1676.865 2803.465 ;
        RECT 1675.630 2803.150 1676.865 2803.450 ;
        RECT 1676.535 2803.135 1676.865 2803.150 ;
        RECT 1786.950 2802.785 1787.250 2803.815 ;
        RECT 1883.550 2802.785 1883.850 2804.495 ;
        RECT 1400.535 2802.455 1400.865 2802.785 ;
        RECT 1544.975 2802.455 1545.305 2802.785 ;
        RECT 1786.935 2802.455 1787.265 2802.785 ;
        RECT 1883.535 2802.455 1883.865 2802.785 ;
        RECT 1544.990 2802.105 1545.290 2802.455 ;
        RECT 1544.975 2801.775 1545.305 2802.105 ;
        RECT 2238.655 2801.095 2238.985 2801.425 ;
        RECT 2238.670 1023.225 2238.970 2801.095 ;
        RECT 2238.655 1022.895 2238.985 1023.225 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1298.190 2812.380 1298.510 2812.440 ;
        RECT 2904.510 2812.380 2904.830 2812.440 ;
        RECT 1298.190 2812.240 2904.830 2812.380 ;
        RECT 1298.190 2812.180 1298.510 2812.240 ;
        RECT 2904.510 2812.180 2904.830 2812.240 ;
      LAYER via ;
        RECT 1298.220 2812.180 1298.480 2812.440 ;
        RECT 2904.540 2812.180 2904.800 2812.440 ;
      LAYER met2 ;
        RECT 1298.220 2812.150 1298.480 2812.470 ;
        RECT 2904.540 2812.150 2904.800 2812.470 ;
        RECT 1298.280 2800.000 1298.420 2812.150 ;
        RECT 1298.145 2796.000 1298.425 2800.000 ;
        RECT 2904.600 1261.245 2904.740 2812.150 ;
        RECT 2904.530 1260.875 2904.810 1261.245 ;
      LAYER via2 ;
        RECT 2904.530 1260.920 2904.810 1261.200 ;
      LAYER met3 ;
        RECT 2904.505 1261.210 2904.835 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2904.505 1260.910 2924.800 1261.210 ;
        RECT 2904.505 1260.895 2904.835 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1952.845 2799.305 1953.935 2799.475 ;
        RECT 2097.745 2799.305 2098.375 2799.475 ;
      LAYER mcon ;
        RECT 1953.765 2799.305 1953.935 2799.475 ;
        RECT 2098.205 2799.305 2098.375 2799.475 ;
      LAYER met1 ;
        RECT 1329.010 2799.460 1329.330 2799.520 ;
        RECT 1861.230 2799.460 1861.550 2799.520 ;
        RECT 1329.010 2799.320 1861.550 2799.460 ;
        RECT 1329.010 2799.260 1329.330 2799.320 ;
        RECT 1861.230 2799.260 1861.550 2799.320 ;
        RECT 1945.410 2799.460 1945.730 2799.520 ;
        RECT 1952.785 2799.460 1953.075 2799.505 ;
        RECT 1945.410 2799.320 1953.075 2799.460 ;
        RECT 1945.410 2799.260 1945.730 2799.320 ;
        RECT 1952.785 2799.275 1953.075 2799.320 ;
        RECT 1953.705 2799.460 1953.995 2799.505 ;
        RECT 2001.530 2799.460 2001.850 2799.520 ;
        RECT 1953.705 2799.320 2001.850 2799.460 ;
        RECT 1953.705 2799.275 1953.995 2799.320 ;
        RECT 2001.530 2799.260 2001.850 2799.320 ;
        RECT 2003.370 2799.460 2003.690 2799.520 ;
        RECT 2049.370 2799.460 2049.690 2799.520 ;
        RECT 2003.370 2799.320 2049.690 2799.460 ;
        RECT 2003.370 2799.260 2003.690 2799.320 ;
        RECT 2049.370 2799.260 2049.690 2799.320 ;
        RECT 2096.750 2799.460 2097.070 2799.520 ;
        RECT 2097.685 2799.460 2097.975 2799.505 ;
        RECT 2096.750 2799.320 2097.975 2799.460 ;
        RECT 2096.750 2799.260 2097.070 2799.320 ;
        RECT 2097.685 2799.275 2097.975 2799.320 ;
        RECT 2098.145 2799.460 2098.435 2799.505 ;
        RECT 2887.490 2799.460 2887.810 2799.520 ;
        RECT 2098.145 2799.320 2887.810 2799.460 ;
        RECT 2098.145 2799.275 2098.435 2799.320 ;
        RECT 2887.490 2799.260 2887.810 2799.320 ;
        RECT 2887.490 1497.260 2887.810 1497.320 ;
        RECT 2899.450 1497.260 2899.770 1497.320 ;
        RECT 2887.490 1497.120 2899.770 1497.260 ;
        RECT 2887.490 1497.060 2887.810 1497.120 ;
        RECT 2899.450 1497.060 2899.770 1497.120 ;
      LAYER via ;
        RECT 1329.040 2799.260 1329.300 2799.520 ;
        RECT 1861.260 2799.260 1861.520 2799.520 ;
        RECT 1945.440 2799.260 1945.700 2799.520 ;
        RECT 2001.560 2799.260 2001.820 2799.520 ;
        RECT 2003.400 2799.260 2003.660 2799.520 ;
        RECT 2049.400 2799.260 2049.660 2799.520 ;
        RECT 2096.780 2799.260 2097.040 2799.520 ;
        RECT 2887.520 2799.260 2887.780 2799.520 ;
        RECT 2887.520 1497.060 2887.780 1497.320 ;
        RECT 2899.480 1497.060 2899.740 1497.320 ;
      LAYER met2 ;
        RECT 1861.250 2800.395 1861.530 2800.765 ;
        RECT 1945.430 2800.395 1945.710 2800.765 ;
        RECT 1327.125 2799.290 1327.405 2800.000 ;
        RECT 1861.320 2799.550 1861.460 2800.395 ;
        RECT 1945.500 2799.550 1945.640 2800.395 ;
        RECT 1329.040 2799.290 1329.300 2799.550 ;
        RECT 1327.125 2799.230 1329.300 2799.290 ;
        RECT 1861.260 2799.230 1861.520 2799.550 ;
        RECT 1945.440 2799.230 1945.700 2799.550 ;
        RECT 2001.560 2799.405 2001.820 2799.550 ;
        RECT 2003.400 2799.405 2003.660 2799.550 ;
        RECT 2049.400 2799.405 2049.660 2799.550 ;
        RECT 2096.780 2799.405 2097.040 2799.550 ;
        RECT 1327.125 2799.150 1329.240 2799.230 ;
        RECT 1327.125 2796.000 1327.405 2799.150 ;
        RECT 2001.550 2799.035 2001.830 2799.405 ;
        RECT 2003.390 2799.035 2003.670 2799.405 ;
        RECT 2049.390 2799.035 2049.670 2799.405 ;
        RECT 2096.770 2799.035 2097.050 2799.405 ;
        RECT 2887.520 2799.230 2887.780 2799.550 ;
        RECT 2887.580 1497.350 2887.720 2799.230 ;
        RECT 2887.520 1497.030 2887.780 1497.350 ;
        RECT 2899.480 1497.030 2899.740 1497.350 ;
        RECT 2899.540 1495.845 2899.680 1497.030 ;
        RECT 2899.470 1495.475 2899.750 1495.845 ;
      LAYER via2 ;
        RECT 1861.250 2800.440 1861.530 2800.720 ;
        RECT 1945.430 2800.440 1945.710 2800.720 ;
        RECT 2001.550 2799.080 2001.830 2799.360 ;
        RECT 2003.390 2799.080 2003.670 2799.360 ;
        RECT 2049.390 2799.080 2049.670 2799.360 ;
        RECT 2096.770 2799.080 2097.050 2799.360 ;
        RECT 2899.470 1495.520 2899.750 1495.800 ;
      LAYER met3 ;
        RECT 1861.225 2800.730 1861.555 2800.745 ;
        RECT 1945.405 2800.730 1945.735 2800.745 ;
        RECT 1861.225 2800.430 1945.735 2800.730 ;
        RECT 1861.225 2800.415 1861.555 2800.430 ;
        RECT 1945.405 2800.415 1945.735 2800.430 ;
        RECT 2001.525 2799.370 2001.855 2799.385 ;
        RECT 2003.365 2799.370 2003.695 2799.385 ;
        RECT 2001.525 2799.070 2003.695 2799.370 ;
        RECT 2001.525 2799.055 2001.855 2799.070 ;
        RECT 2003.365 2799.055 2003.695 2799.070 ;
        RECT 2049.365 2799.370 2049.695 2799.385 ;
        RECT 2096.745 2799.370 2097.075 2799.385 ;
        RECT 2049.365 2799.070 2097.075 2799.370 ;
        RECT 2049.365 2799.055 2049.695 2799.070 ;
        RECT 2096.745 2799.055 2097.075 2799.070 ;
        RECT 2899.445 1495.810 2899.775 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2899.445 1495.510 2924.800 1495.810 ;
        RECT 2899.445 1495.495 2899.775 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2001.605 2803.385 2002.695 2803.555 ;
      LAYER mcon ;
        RECT 2002.525 2803.385 2002.695 2803.555 ;
      LAYER met1 ;
        RECT 1356.150 2803.540 1356.470 2803.600 ;
        RECT 2001.545 2803.540 2001.835 2803.585 ;
        RECT 1356.150 2803.400 2001.835 2803.540 ;
        RECT 1356.150 2803.340 1356.470 2803.400 ;
        RECT 2001.545 2803.355 2001.835 2803.400 ;
        RECT 2002.465 2803.540 2002.755 2803.585 ;
        RECT 2252.690 2803.540 2253.010 2803.600 ;
        RECT 2002.465 2803.400 2253.010 2803.540 ;
        RECT 2002.465 2803.355 2002.755 2803.400 ;
        RECT 2252.690 2803.340 2253.010 2803.400 ;
        RECT 2252.690 1731.860 2253.010 1731.920 ;
        RECT 2899.450 1731.860 2899.770 1731.920 ;
        RECT 2252.690 1731.720 2899.770 1731.860 ;
        RECT 2252.690 1731.660 2253.010 1731.720 ;
        RECT 2899.450 1731.660 2899.770 1731.720 ;
      LAYER via ;
        RECT 1356.180 2803.340 1356.440 2803.600 ;
        RECT 2252.720 2803.340 2252.980 2803.600 ;
        RECT 2252.720 1731.660 2252.980 1731.920 ;
        RECT 2899.480 1731.660 2899.740 1731.920 ;
      LAYER met2 ;
        RECT 1356.180 2803.310 1356.440 2803.630 ;
        RECT 2252.720 2803.310 2252.980 2803.630 ;
        RECT 1356.240 2800.000 1356.380 2803.310 ;
        RECT 1356.105 2796.000 1356.385 2800.000 ;
        RECT 2252.780 1731.950 2252.920 2803.310 ;
        RECT 2252.720 1731.630 2252.980 1731.950 ;
        RECT 2899.480 1731.630 2899.740 1731.950 ;
        RECT 2899.540 1730.445 2899.680 1731.630 ;
        RECT 2899.470 1730.075 2899.750 1730.445 ;
      LAYER via2 ;
        RECT 2899.470 1730.120 2899.750 1730.400 ;
      LAYER met3 ;
        RECT 2899.445 1730.410 2899.775 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2899.445 1730.110 2924.800 1730.410 ;
        RECT 2899.445 1730.095 2899.775 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1385.130 2803.880 1385.450 2803.940 ;
        RECT 2001.070 2803.880 2001.390 2803.940 ;
        RECT 1385.130 2803.740 2001.390 2803.880 ;
        RECT 1385.130 2803.680 1385.450 2803.740 ;
        RECT 2001.070 2803.680 2001.390 2803.740 ;
        RECT 2002.910 2803.880 2003.230 2803.940 ;
        RECT 2248.090 2803.880 2248.410 2803.940 ;
        RECT 2002.910 2803.740 2248.410 2803.880 ;
        RECT 2002.910 2803.680 2003.230 2803.740 ;
        RECT 2248.090 2803.680 2248.410 2803.740 ;
        RECT 2248.550 1966.460 2248.870 1966.520 ;
        RECT 2898.990 1966.460 2899.310 1966.520 ;
        RECT 2248.550 1966.320 2899.310 1966.460 ;
        RECT 2248.550 1966.260 2248.870 1966.320 ;
        RECT 2898.990 1966.260 2899.310 1966.320 ;
      LAYER via ;
        RECT 1385.160 2803.680 1385.420 2803.940 ;
        RECT 2001.100 2803.680 2001.360 2803.940 ;
        RECT 2002.940 2803.680 2003.200 2803.940 ;
        RECT 2248.120 2803.680 2248.380 2803.940 ;
        RECT 2248.580 1966.260 2248.840 1966.520 ;
        RECT 2899.020 1966.260 2899.280 1966.520 ;
      LAYER met2 ;
        RECT 1385.160 2803.650 1385.420 2803.970 ;
        RECT 2001.090 2803.795 2001.370 2804.165 ;
        RECT 2002.930 2803.795 2003.210 2804.165 ;
        RECT 2001.100 2803.650 2001.360 2803.795 ;
        RECT 2002.940 2803.650 2003.200 2803.795 ;
        RECT 2248.120 2803.650 2248.380 2803.970 ;
        RECT 1385.220 2800.000 1385.360 2803.650 ;
        RECT 1385.085 2796.000 1385.365 2800.000 ;
        RECT 2248.180 1973.090 2248.320 2803.650 ;
        RECT 2248.180 1972.950 2248.780 1973.090 ;
        RECT 2248.640 1966.550 2248.780 1972.950 ;
        RECT 2248.580 1966.230 2248.840 1966.550 ;
        RECT 2899.020 1966.230 2899.280 1966.550 ;
        RECT 2899.080 1965.045 2899.220 1966.230 ;
        RECT 2899.010 1964.675 2899.290 1965.045 ;
      LAYER via2 ;
        RECT 2001.090 2803.840 2001.370 2804.120 ;
        RECT 2002.930 2803.840 2003.210 2804.120 ;
        RECT 2899.010 1964.720 2899.290 1965.000 ;
      LAYER met3 ;
        RECT 2001.065 2804.130 2001.395 2804.145 ;
        RECT 2002.905 2804.130 2003.235 2804.145 ;
        RECT 2001.065 2803.830 2003.235 2804.130 ;
        RECT 2001.065 2803.815 2001.395 2803.830 ;
        RECT 2002.905 2803.815 2003.235 2803.830 ;
        RECT 2898.985 1965.010 2899.315 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.985 1964.710 2924.800 1965.010 ;
        RECT 2898.985 1964.695 2899.315 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2001.605 2804.065 2002.695 2804.235 ;
      LAYER mcon ;
        RECT 2002.525 2804.065 2002.695 2804.235 ;
      LAYER met1 ;
        RECT 1414.110 2804.220 1414.430 2804.280 ;
        RECT 2001.545 2804.220 2001.835 2804.265 ;
        RECT 1414.110 2804.080 2001.835 2804.220 ;
        RECT 1414.110 2804.020 1414.430 2804.080 ;
        RECT 2001.545 2804.035 2001.835 2804.080 ;
        RECT 2002.465 2804.220 2002.755 2804.265 ;
        RECT 2251.310 2804.220 2251.630 2804.280 ;
        RECT 2002.465 2804.080 2251.630 2804.220 ;
        RECT 2002.465 2804.035 2002.755 2804.080 ;
        RECT 2251.310 2804.020 2251.630 2804.080 ;
        RECT 2251.310 2786.540 2251.630 2786.600 ;
        RECT 2254.530 2786.540 2254.850 2786.600 ;
        RECT 2251.310 2786.400 2254.850 2786.540 ;
        RECT 2251.310 2786.340 2251.630 2786.400 ;
        RECT 2254.530 2786.340 2254.850 2786.400 ;
        RECT 2254.530 2201.060 2254.850 2201.120 ;
        RECT 2898.990 2201.060 2899.310 2201.120 ;
        RECT 2254.530 2200.920 2899.310 2201.060 ;
        RECT 2254.530 2200.860 2254.850 2200.920 ;
        RECT 2898.990 2200.860 2899.310 2200.920 ;
      LAYER via ;
        RECT 1414.140 2804.020 1414.400 2804.280 ;
        RECT 2251.340 2804.020 2251.600 2804.280 ;
        RECT 2251.340 2786.340 2251.600 2786.600 ;
        RECT 2254.560 2786.340 2254.820 2786.600 ;
        RECT 2254.560 2200.860 2254.820 2201.120 ;
        RECT 2899.020 2200.860 2899.280 2201.120 ;
      LAYER met2 ;
        RECT 1414.140 2803.990 1414.400 2804.310 ;
        RECT 2251.340 2803.990 2251.600 2804.310 ;
        RECT 1414.200 2800.000 1414.340 2803.990 ;
        RECT 1414.065 2796.000 1414.345 2800.000 ;
        RECT 2251.400 2786.630 2251.540 2803.990 ;
        RECT 2251.340 2786.310 2251.600 2786.630 ;
        RECT 2254.560 2786.310 2254.820 2786.630 ;
        RECT 2254.620 2201.150 2254.760 2786.310 ;
        RECT 2254.560 2200.830 2254.820 2201.150 ;
        RECT 2899.020 2200.830 2899.280 2201.150 ;
        RECT 2899.080 2199.645 2899.220 2200.830 ;
        RECT 2899.010 2199.275 2899.290 2199.645 ;
      LAYER via2 ;
        RECT 2899.010 2199.320 2899.290 2199.600 ;
      LAYER met3 ;
        RECT 2898.985 2199.610 2899.315 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.985 2199.310 2924.800 2199.610 ;
        RECT 2898.985 2199.295 2899.315 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 201.860 1352.790 201.920 ;
        RECT 1402.610 201.860 1402.930 201.920 ;
        RECT 1352.470 201.720 1402.930 201.860 ;
        RECT 1352.470 201.660 1352.790 201.720 ;
        RECT 1402.610 201.660 1402.930 201.720 ;
        RECT 1992.330 201.180 1992.650 201.240 ;
        RECT 1995.090 201.180 1995.410 201.240 ;
        RECT 1992.330 201.040 1995.410 201.180 ;
        RECT 1992.330 200.980 1992.650 201.040 ;
        RECT 1995.090 200.980 1995.410 201.040 ;
        RECT 2089.390 201.180 2089.710 201.240 ;
        RECT 2091.690 201.180 2092.010 201.240 ;
        RECT 2089.390 201.040 2092.010 201.180 ;
        RECT 2089.390 200.980 2089.710 201.040 ;
        RECT 2091.690 200.980 2092.010 201.040 ;
        RECT 1780.270 200.500 1780.590 200.560 ;
        RECT 1828.110 200.500 1828.430 200.560 ;
        RECT 1780.270 200.360 1828.430 200.500 ;
        RECT 1780.270 200.300 1780.590 200.360 ;
        RECT 1828.110 200.300 1828.430 200.360 ;
      LAYER via ;
        RECT 1352.500 201.660 1352.760 201.920 ;
        RECT 1402.640 201.660 1402.900 201.920 ;
        RECT 1992.360 200.980 1992.620 201.240 ;
        RECT 1995.120 200.980 1995.380 201.240 ;
        RECT 2089.420 200.980 2089.680 201.240 ;
        RECT 2091.720 200.980 2091.980 201.240 ;
        RECT 1780.300 200.300 1780.560 200.560 ;
        RECT 1828.140 200.300 1828.400 200.560 ;
      LAYER met2 ;
        RECT 1162.905 2796.570 1163.185 2800.000 ;
        RECT 1164.350 2796.570 1164.630 2796.685 ;
        RECT 1162.905 2796.430 1164.630 2796.570 ;
        RECT 1162.905 2796.000 1163.185 2796.430 ;
        RECT 1164.350 2796.315 1164.630 2796.430 ;
        RECT 2304.230 203.475 2304.510 203.845 ;
        RECT 1641.830 202.795 1642.110 203.165 ;
        RECT 1689.670 202.795 1689.950 203.165 ;
        RECT 1352.500 201.805 1352.760 201.950 ;
        RECT 1402.640 201.805 1402.900 201.950 ;
        RECT 1352.490 201.435 1352.770 201.805 ;
        RECT 1402.630 201.435 1402.910 201.805 ;
        RECT 1487.730 201.435 1488.010 201.805 ;
        RECT 1487.800 200.445 1487.940 201.435 ;
        RECT 1641.900 201.125 1642.040 202.795 ;
        RECT 1641.830 200.755 1642.110 201.125 ;
        RECT 1689.740 200.445 1689.880 202.795 ;
        RECT 2236.150 202.115 2236.430 202.485 ;
        RECT 1992.360 201.125 1992.620 201.270 ;
        RECT 1995.120 201.125 1995.380 201.270 ;
        RECT 2089.420 201.125 2089.680 201.270 ;
        RECT 2091.720 201.125 2091.980 201.270 ;
        RECT 1780.290 200.755 1780.570 201.125 ;
        RECT 1992.350 200.755 1992.630 201.125 ;
        RECT 1995.110 200.755 1995.390 201.125 ;
        RECT 2089.410 200.755 2089.690 201.125 ;
        RECT 2091.710 200.755 2091.990 201.125 ;
        RECT 2235.690 201.010 2235.970 201.125 ;
        RECT 2236.220 201.010 2236.360 202.115 ;
        RECT 2304.300 201.805 2304.440 203.475 ;
        RECT 2304.230 201.435 2304.510 201.805 ;
        RECT 2235.690 200.870 2236.360 201.010 ;
        RECT 2235.690 200.755 2235.970 200.870 ;
        RECT 1780.360 200.590 1780.500 200.755 ;
        RECT 1487.730 200.075 1488.010 200.445 ;
        RECT 1689.670 200.075 1689.950 200.445 ;
        RECT 1780.300 200.270 1780.560 200.590 ;
        RECT 1828.140 200.445 1828.400 200.590 ;
        RECT 1828.130 200.075 1828.410 200.445 ;
      LAYER via2 ;
        RECT 1164.350 2796.360 1164.630 2796.640 ;
        RECT 2304.230 203.520 2304.510 203.800 ;
        RECT 1641.830 202.840 1642.110 203.120 ;
        RECT 1689.670 202.840 1689.950 203.120 ;
        RECT 1352.490 201.480 1352.770 201.760 ;
        RECT 1402.630 201.480 1402.910 201.760 ;
        RECT 1487.730 201.480 1488.010 201.760 ;
        RECT 1641.830 200.800 1642.110 201.080 ;
        RECT 2236.150 202.160 2236.430 202.440 ;
        RECT 1780.290 200.800 1780.570 201.080 ;
        RECT 1992.350 200.800 1992.630 201.080 ;
        RECT 1995.110 200.800 1995.390 201.080 ;
        RECT 2089.410 200.800 2089.690 201.080 ;
        RECT 2091.710 200.800 2091.990 201.080 ;
        RECT 2235.690 200.800 2235.970 201.080 ;
        RECT 2304.230 201.480 2304.510 201.760 ;
        RECT 1487.730 200.120 1488.010 200.400 ;
        RECT 1689.670 200.120 1689.950 200.400 ;
        RECT 1828.130 200.120 1828.410 200.400 ;
      LAYER met3 ;
        RECT 1164.325 2796.650 1164.655 2796.665 ;
        RECT 1164.990 2796.650 1165.370 2796.660 ;
        RECT 1164.325 2796.350 1165.370 2796.650 ;
        RECT 1164.325 2796.335 1164.655 2796.350 ;
        RECT 1164.990 2796.340 1165.370 2796.350 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 2269.910 203.810 2270.290 203.820 ;
        RECT 2304.205 203.810 2304.535 203.825 ;
        RECT 2269.910 203.510 2304.535 203.810 ;
        RECT 2269.910 203.500 2270.290 203.510 ;
        RECT 2304.205 203.495 2304.535 203.510 ;
        RECT 1641.805 203.130 1642.135 203.145 ;
        RECT 1689.645 203.130 1689.975 203.145 ;
        RECT 1641.805 202.830 1689.975 203.130 ;
        RECT 1641.805 202.815 1642.135 202.830 ;
        RECT 1689.645 202.815 1689.975 202.830 ;
        RECT 2236.125 202.450 2236.455 202.465 ;
        RECT 2269.910 202.450 2270.290 202.460 ;
        RECT 1883.550 202.150 1931.690 202.450 ;
        RECT 1248.710 201.770 1249.090 201.780 ;
        RECT 1352.465 201.770 1352.795 201.785 ;
        RECT 1248.710 201.470 1352.795 201.770 ;
        RECT 1248.710 201.460 1249.090 201.470 ;
        RECT 1352.465 201.455 1352.795 201.470 ;
        RECT 1402.605 201.770 1402.935 201.785 ;
        RECT 1487.705 201.770 1488.035 201.785 ;
        RECT 1402.605 201.470 1448.690 201.770 ;
        RECT 1402.605 201.455 1402.935 201.470 ;
        RECT 1448.390 201.090 1448.690 201.470 ;
        RECT 1449.310 201.470 1488.035 201.770 ;
        RECT 1449.310 201.090 1449.610 201.470 ;
        RECT 1487.705 201.455 1488.035 201.470 ;
        RECT 1641.805 201.090 1642.135 201.105 ;
        RECT 1780.265 201.090 1780.595 201.105 ;
        RECT 1883.550 201.090 1883.850 202.150 ;
        RECT 1448.390 200.790 1449.610 201.090 ;
        RECT 1562.470 200.790 1642.135 201.090 ;
        RECT 1164.990 200.410 1165.370 200.420 ;
        RECT 1248.710 200.410 1249.090 200.420 ;
        RECT 1164.990 200.110 1249.090 200.410 ;
        RECT 1164.990 200.100 1165.370 200.110 ;
        RECT 1248.710 200.100 1249.090 200.110 ;
        RECT 1487.705 200.410 1488.035 200.425 ;
        RECT 1562.470 200.410 1562.770 200.790 ;
        RECT 1641.805 200.775 1642.135 200.790 ;
        RECT 1752.910 200.790 1780.595 201.090 ;
        RECT 1487.705 200.110 1562.770 200.410 ;
        RECT 1689.645 200.410 1689.975 200.425 ;
        RECT 1752.910 200.410 1753.210 200.790 ;
        RECT 1780.265 200.775 1780.595 200.790 ;
        RECT 1849.510 200.790 1883.850 201.090 ;
        RECT 1689.645 200.110 1753.210 200.410 ;
        RECT 1828.105 200.410 1828.435 200.425 ;
        RECT 1849.510 200.410 1849.810 200.790 ;
        RECT 1828.105 200.110 1849.810 200.410 ;
        RECT 1931.390 200.410 1931.690 202.150 ;
        RECT 2236.125 202.150 2270.290 202.450 ;
        RECT 2236.125 202.135 2236.455 202.150 ;
        RECT 2269.910 202.140 2270.290 202.150 ;
        RECT 2304.205 201.770 2304.535 201.785 ;
        RECT 2304.205 201.470 2353.050 201.770 ;
        RECT 2304.205 201.455 2304.535 201.470 ;
        RECT 1992.325 201.090 1992.655 201.105 ;
        RECT 1946.110 200.790 1992.655 201.090 ;
        RECT 1946.110 200.410 1946.410 200.790 ;
        RECT 1992.325 200.775 1992.655 200.790 ;
        RECT 1995.085 201.090 1995.415 201.105 ;
        RECT 2089.385 201.090 2089.715 201.105 ;
        RECT 1995.085 200.790 2028.290 201.090 ;
        RECT 1995.085 200.775 1995.415 200.790 ;
        RECT 1931.390 200.110 1946.410 200.410 ;
        RECT 2027.990 200.410 2028.290 200.790 ;
        RECT 2042.710 200.790 2089.715 201.090 ;
        RECT 2042.710 200.410 2043.010 200.790 ;
        RECT 2089.385 200.775 2089.715 200.790 ;
        RECT 2091.685 201.090 2092.015 201.105 ;
        RECT 2235.665 201.090 2235.995 201.105 ;
        RECT 2091.685 200.790 2124.890 201.090 ;
        RECT 2091.685 200.775 2092.015 200.790 ;
        RECT 2027.990 200.110 2043.010 200.410 ;
        RECT 2124.590 200.410 2124.890 200.790 ;
        RECT 2139.310 200.790 2235.995 201.090 ;
        RECT 2352.750 201.090 2353.050 201.470 ;
        RECT 2401.510 201.470 2449.650 201.770 ;
        RECT 2352.750 200.790 2400.890 201.090 ;
        RECT 2139.310 200.410 2139.610 200.790 ;
        RECT 2235.665 200.775 2235.995 200.790 ;
        RECT 2124.590 200.110 2139.610 200.410 ;
        RECT 2400.590 200.410 2400.890 200.790 ;
        RECT 2401.510 200.410 2401.810 201.470 ;
        RECT 2449.350 201.090 2449.650 201.470 ;
        RECT 2498.110 201.470 2546.250 201.770 ;
        RECT 2449.350 200.790 2497.490 201.090 ;
        RECT 2400.590 200.110 2401.810 200.410 ;
        RECT 2497.190 200.410 2497.490 200.790 ;
        RECT 2498.110 200.410 2498.410 201.470 ;
        RECT 2545.950 201.090 2546.250 201.470 ;
        RECT 2594.710 201.470 2642.850 201.770 ;
        RECT 2545.950 200.790 2594.090 201.090 ;
        RECT 2497.190 200.110 2498.410 200.410 ;
        RECT 2593.790 200.410 2594.090 200.790 ;
        RECT 2594.710 200.410 2595.010 201.470 ;
        RECT 2642.550 201.090 2642.850 201.470 ;
        RECT 2691.310 201.470 2739.450 201.770 ;
        RECT 2642.550 200.790 2690.690 201.090 ;
        RECT 2593.790 200.110 2595.010 200.410 ;
        RECT 2690.390 200.410 2690.690 200.790 ;
        RECT 2691.310 200.410 2691.610 201.470 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2690.390 200.110 2691.610 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2883.590 200.110 2884.810 200.410 ;
        RECT 1487.705 200.095 1488.035 200.110 ;
        RECT 1689.645 200.095 1689.975 200.110 ;
        RECT 1828.105 200.095 1828.435 200.110 ;
      LAYER via3 ;
        RECT 1165.020 2796.340 1165.340 2796.660 ;
        RECT 2269.940 203.500 2270.260 203.820 ;
        RECT 1248.740 201.460 1249.060 201.780 ;
        RECT 1165.020 200.100 1165.340 200.420 ;
        RECT 1248.740 200.100 1249.060 200.420 ;
        RECT 2269.940 202.140 2270.260 202.460 ;
      LAYER met4 ;
        RECT 1165.015 2796.335 1165.345 2796.665 ;
        RECT 1165.030 200.425 1165.330 2796.335 ;
        RECT 2269.935 203.495 2270.265 203.825 ;
        RECT 2269.950 202.465 2270.250 203.495 ;
        RECT 2269.935 202.135 2270.265 202.465 ;
        RECT 1248.735 201.455 1249.065 201.785 ;
        RECT 1248.750 200.425 1249.050 201.455 ;
        RECT 1165.015 200.095 1165.345 200.425 ;
        RECT 1248.735 200.095 1249.065 200.425 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2001.145 2804.405 2002.235 2804.575 ;
      LAYER mcon ;
        RECT 2002.065 2804.405 2002.235 2804.575 ;
      LAYER met1 ;
        RECT 1452.750 2804.560 1453.070 2804.620 ;
        RECT 2001.085 2804.560 2001.375 2804.605 ;
        RECT 1452.750 2804.420 2001.375 2804.560 ;
        RECT 1452.750 2804.360 1453.070 2804.420 ;
        RECT 2001.085 2804.375 2001.375 2804.420 ;
        RECT 2002.005 2804.560 2002.295 2804.605 ;
        RECT 2255.910 2804.560 2256.230 2804.620 ;
        RECT 2002.005 2804.420 2256.230 2804.560 ;
        RECT 2002.005 2804.375 2002.295 2804.420 ;
        RECT 2255.910 2804.360 2256.230 2804.420 ;
        RECT 2255.910 2552.960 2256.230 2553.020 ;
        RECT 2898.990 2552.960 2899.310 2553.020 ;
        RECT 2255.910 2552.820 2899.310 2552.960 ;
        RECT 2255.910 2552.760 2256.230 2552.820 ;
        RECT 2898.990 2552.760 2899.310 2552.820 ;
      LAYER via ;
        RECT 1452.780 2804.360 1453.040 2804.620 ;
        RECT 2255.940 2804.360 2256.200 2804.620 ;
        RECT 2255.940 2552.760 2256.200 2553.020 ;
        RECT 2899.020 2552.760 2899.280 2553.020 ;
      LAYER met2 ;
        RECT 1452.780 2804.330 1453.040 2804.650 ;
        RECT 2255.940 2804.330 2256.200 2804.650 ;
        RECT 1452.840 2800.000 1452.980 2804.330 ;
        RECT 1452.705 2796.000 1452.985 2800.000 ;
        RECT 2256.000 2553.050 2256.140 2804.330 ;
        RECT 2255.940 2552.730 2256.200 2553.050 ;
        RECT 2899.020 2552.730 2899.280 2553.050 ;
        RECT 2899.080 2551.885 2899.220 2552.730 ;
        RECT 2899.010 2551.515 2899.290 2551.885 ;
      LAYER via2 ;
        RECT 2899.010 2551.560 2899.290 2551.840 ;
      LAYER met3 ;
        RECT 2898.985 2551.850 2899.315 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2898.985 2551.550 2924.800 2551.850 ;
        RECT 2898.985 2551.535 2899.315 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1481.730 2804.900 1482.050 2804.960 ;
        RECT 2254.070 2804.900 2254.390 2804.960 ;
        RECT 1481.730 2804.760 2254.390 2804.900 ;
        RECT 1481.730 2804.700 1482.050 2804.760 ;
        RECT 2254.070 2804.700 2254.390 2804.760 ;
        RECT 2254.070 2787.560 2254.390 2787.620 ;
        RECT 2898.530 2787.560 2898.850 2787.620 ;
        RECT 2254.070 2787.420 2898.850 2787.560 ;
        RECT 2254.070 2787.360 2254.390 2787.420 ;
        RECT 2898.530 2787.360 2898.850 2787.420 ;
      LAYER via ;
        RECT 1481.760 2804.700 1482.020 2804.960 ;
        RECT 2254.100 2804.700 2254.360 2804.960 ;
        RECT 2254.100 2787.360 2254.360 2787.620 ;
        RECT 2898.560 2787.360 2898.820 2787.620 ;
      LAYER met2 ;
        RECT 1481.760 2804.670 1482.020 2804.990 ;
        RECT 2254.100 2804.670 2254.360 2804.990 ;
        RECT 1481.820 2800.000 1481.960 2804.670 ;
        RECT 1481.685 2796.000 1481.965 2800.000 ;
        RECT 2254.160 2787.650 2254.300 2804.670 ;
        RECT 2254.100 2787.330 2254.360 2787.650 ;
        RECT 2898.560 2787.330 2898.820 2787.650 ;
        RECT 2898.620 2786.485 2898.760 2787.330 ;
        RECT 2898.550 2786.115 2898.830 2786.485 ;
      LAYER via2 ;
        RECT 2898.550 2786.160 2898.830 2786.440 ;
      LAYER met3 ;
        RECT 2898.525 2786.450 2898.855 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2898.525 2786.150 2924.800 2786.450 ;
        RECT 2898.525 2786.135 2898.855 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1510.710 3015.700 1511.030 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1510.710 3015.560 2901.150 3015.700 ;
        RECT 1510.710 3015.500 1511.030 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1510.740 3015.500 1511.000 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1510.740 3015.470 1511.000 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1510.800 2800.000 1510.940 3015.470 ;
        RECT 1510.665 2796.000 1510.945 2800.000 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1545.210 3250.300 1545.530 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1545.210 3250.160 2901.150 3250.300 ;
        RECT 1545.210 3250.100 1545.530 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 1538.770 2825.640 1539.090 2825.700 ;
        RECT 1545.210 2825.640 1545.530 2825.700 ;
        RECT 1538.770 2825.500 1545.530 2825.640 ;
        RECT 1538.770 2825.440 1539.090 2825.500 ;
        RECT 1545.210 2825.440 1545.530 2825.500 ;
      LAYER via ;
        RECT 1545.240 3250.100 1545.500 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 1538.800 2825.440 1539.060 2825.700 ;
        RECT 1545.240 2825.440 1545.500 2825.700 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1545.240 3250.070 1545.500 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1545.300 2825.730 1545.440 3250.070 ;
        RECT 1538.800 2825.410 1539.060 2825.730 ;
        RECT 1545.240 2825.410 1545.500 2825.730 ;
        RECT 1538.860 2799.970 1539.000 2825.410 ;
        RECT 1539.185 2799.970 1539.465 2800.000 ;
        RECT 1538.860 2799.830 1539.465 2799.970 ;
        RECT 1539.185 2796.000 1539.465 2799.830 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1572.810 3484.900 1573.130 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1572.810 3484.760 2901.150 3484.900 ;
        RECT 1572.810 3484.700 1573.130 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 1566.370 2825.640 1566.690 2825.700 ;
        RECT 1572.810 2825.640 1573.130 2825.700 ;
        RECT 1566.370 2825.500 1573.130 2825.640 ;
        RECT 1566.370 2825.440 1566.690 2825.500 ;
        RECT 1572.810 2825.440 1573.130 2825.500 ;
      LAYER via ;
        RECT 1572.840 3484.700 1573.100 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 1566.400 2825.440 1566.660 2825.700 ;
        RECT 1572.840 2825.440 1573.100 2825.700 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1572.840 3484.670 1573.100 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1572.900 2825.730 1573.040 3484.670 ;
        RECT 1566.400 2825.410 1566.660 2825.730 ;
        RECT 1572.840 2825.410 1573.100 2825.730 ;
        RECT 1566.460 2799.970 1566.600 2825.410 ;
        RECT 1568.165 2799.970 1568.445 2800.000 ;
        RECT 1566.460 2799.830 1568.445 2799.970 ;
        RECT 1568.165 2796.000 1568.445 2799.830 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1600.410 3503.940 1600.730 3504.000 ;
        RECT 2635.870 3503.940 2636.190 3504.000 ;
        RECT 1600.410 3503.800 2636.190 3503.940 ;
        RECT 1600.410 3503.740 1600.730 3503.800 ;
        RECT 2635.870 3503.740 2636.190 3503.800 ;
      LAYER via ;
        RECT 1600.440 3503.740 1600.700 3504.000 ;
        RECT 2635.900 3503.740 2636.160 3504.000 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3504.030 2636.100 3517.600 ;
        RECT 1600.440 3503.710 1600.700 3504.030 ;
        RECT 2635.900 3503.710 2636.160 3504.030 ;
        RECT 1600.500 2800.650 1600.640 3503.710 ;
        RECT 1598.660 2800.510 1600.640 2800.650 ;
        RECT 1597.145 2799.970 1597.425 2800.000 ;
        RECT 1598.660 2799.970 1598.800 2800.510 ;
        RECT 1597.145 2799.830 1598.800 2799.970 ;
        RECT 1597.145 2796.000 1597.425 2799.830 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.010 3500.880 1628.330 3500.940 ;
        RECT 2311.570 3500.880 2311.890 3500.940 ;
        RECT 1628.010 3500.740 2311.890 3500.880 ;
        RECT 1628.010 3500.680 1628.330 3500.740 ;
        RECT 2311.570 3500.680 2311.890 3500.740 ;
      LAYER via ;
        RECT 1628.040 3500.680 1628.300 3500.940 ;
        RECT 2311.600 3500.680 2311.860 3500.940 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3500.970 2311.800 3517.600 ;
        RECT 1628.040 3500.650 1628.300 3500.970 ;
        RECT 2311.600 3500.650 2311.860 3500.970 ;
        RECT 1626.125 2799.970 1626.405 2800.000 ;
        RECT 1628.100 2799.970 1628.240 3500.650 ;
        RECT 1626.125 2799.830 1628.240 2799.970 ;
        RECT 1626.125 2796.000 1626.405 2799.830 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.610 3499.180 1655.930 3499.240 ;
        RECT 1987.270 3499.180 1987.590 3499.240 ;
        RECT 1655.610 3499.040 1987.590 3499.180 ;
        RECT 1655.610 3498.980 1655.930 3499.040 ;
        RECT 1987.270 3498.980 1987.590 3499.040 ;
        RECT 1649.170 2825.640 1649.490 2825.700 ;
        RECT 1655.610 2825.640 1655.930 2825.700 ;
        RECT 1649.170 2825.500 1655.930 2825.640 ;
        RECT 1649.170 2825.440 1649.490 2825.500 ;
        RECT 1655.610 2825.440 1655.930 2825.500 ;
      LAYER via ;
        RECT 1655.640 3498.980 1655.900 3499.240 ;
        RECT 1987.300 3498.980 1987.560 3499.240 ;
        RECT 1649.200 2825.440 1649.460 2825.700 ;
        RECT 1655.640 2825.440 1655.900 2825.700 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3499.270 1987.500 3517.600 ;
        RECT 1655.640 3498.950 1655.900 3499.270 ;
        RECT 1987.300 3498.950 1987.560 3499.270 ;
        RECT 1655.700 2825.730 1655.840 3498.950 ;
        RECT 1649.200 2825.410 1649.460 2825.730 ;
        RECT 1655.640 2825.410 1655.900 2825.730 ;
        RECT 1649.260 2800.650 1649.400 2825.410 ;
        RECT 1649.260 2800.510 1653.540 2800.650 ;
        RECT 1653.400 2799.970 1653.540 2800.510 ;
        RECT 1655.105 2799.970 1655.385 2800.000 ;
        RECT 1653.400 2799.830 1655.385 2799.970 ;
        RECT 1655.105 2796.000 1655.385 2799.830 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3498.500 1662.830 3498.560 ;
        RECT 1683.670 3498.500 1683.990 3498.560 ;
        RECT 1662.510 3498.360 1683.990 3498.500 ;
        RECT 1662.510 3498.300 1662.830 3498.360 ;
        RECT 1683.670 3498.300 1683.990 3498.360 ;
      LAYER via ;
        RECT 1662.540 3498.300 1662.800 3498.560 ;
        RECT 1683.700 3498.300 1683.960 3498.560 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3498.590 1662.740 3517.600 ;
        RECT 1662.540 3498.270 1662.800 3498.590 ;
        RECT 1683.700 3498.270 1683.960 3498.590 ;
        RECT 1683.760 2799.970 1683.900 3498.270 ;
        RECT 1684.085 2799.970 1684.365 2800.000 ;
        RECT 1683.760 2799.830 1684.365 2799.970 ;
        RECT 1684.085 2796.000 1684.365 2799.830 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3499.520 1338.530 3499.580 ;
        RECT 1711.270 3499.520 1711.590 3499.580 ;
        RECT 1338.210 3499.380 1711.590 3499.520 ;
        RECT 1338.210 3499.320 1338.530 3499.380 ;
        RECT 1711.270 3499.320 1711.590 3499.380 ;
      LAYER via ;
        RECT 1338.240 3499.320 1338.500 3499.580 ;
        RECT 1711.300 3499.320 1711.560 3499.580 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3499.610 1338.440 3517.600 ;
        RECT 1338.240 3499.290 1338.500 3499.610 ;
        RECT 1711.300 3499.290 1711.560 3499.610 ;
        RECT 1711.360 2799.970 1711.500 3499.290 ;
        RECT 1713.065 2799.970 1713.345 2800.000 ;
        RECT 1711.360 2799.830 1713.345 2799.970 ;
        RECT 1713.065 2796.000 1713.345 2799.830 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1414.110 436.120 1414.430 436.180 ;
        RECT 1463.790 436.120 1464.110 436.180 ;
        RECT 1414.110 435.980 1464.110 436.120 ;
        RECT 1414.110 435.920 1414.430 435.980 ;
        RECT 1463.790 435.920 1464.110 435.980 ;
        RECT 1780.270 435.780 1780.590 435.840 ;
        RECT 1828.110 435.780 1828.430 435.840 ;
        RECT 1780.270 435.640 1828.430 435.780 ;
        RECT 1780.270 435.580 1780.590 435.640 ;
        RECT 1828.110 435.580 1828.430 435.640 ;
        RECT 2089.390 435.780 2089.710 435.840 ;
        RECT 2091.690 435.780 2092.010 435.840 ;
        RECT 2089.390 435.640 2092.010 435.780 ;
        RECT 2089.390 435.580 2089.710 435.640 ;
        RECT 2091.690 435.580 2092.010 435.640 ;
        RECT 1992.330 435.440 1992.650 435.500 ;
        RECT 1994.170 435.440 1994.490 435.500 ;
        RECT 1992.330 435.300 1994.490 435.440 ;
        RECT 1992.330 435.240 1992.650 435.300 ;
        RECT 1994.170 435.240 1994.490 435.300 ;
        RECT 2221.870 435.100 2222.190 435.160 ;
        RECT 2246.250 435.100 2246.570 435.160 ;
        RECT 2221.870 434.960 2246.570 435.100 ;
        RECT 2221.870 434.900 2222.190 434.960 ;
        RECT 2246.250 434.900 2246.570 434.960 ;
        RECT 2318.930 435.100 2319.250 435.160 ;
        RECT 2332.730 435.100 2333.050 435.160 ;
        RECT 2318.930 434.960 2333.050 435.100 ;
        RECT 2318.930 434.900 2319.250 434.960 ;
        RECT 2332.730 434.900 2333.050 434.960 ;
      LAYER via ;
        RECT 1414.140 435.920 1414.400 436.180 ;
        RECT 1463.820 435.920 1464.080 436.180 ;
        RECT 1780.300 435.580 1780.560 435.840 ;
        RECT 1828.140 435.580 1828.400 435.840 ;
        RECT 2089.420 435.580 2089.680 435.840 ;
        RECT 2091.720 435.580 2091.980 435.840 ;
        RECT 1992.360 435.240 1992.620 435.500 ;
        RECT 1994.200 435.240 1994.460 435.500 ;
        RECT 2221.900 434.900 2222.160 435.160 ;
        RECT 2246.280 434.900 2246.540 435.160 ;
        RECT 2318.960 434.900 2319.220 435.160 ;
        RECT 2332.760 434.900 2333.020 435.160 ;
      LAYER met2 ;
        RECT 1191.030 2796.570 1191.310 2796.685 ;
        RECT 1191.885 2796.570 1192.165 2800.000 ;
        RECT 1191.030 2796.430 1192.165 2796.570 ;
        RECT 1191.030 2796.315 1191.310 2796.430 ;
        RECT 1191.885 2796.000 1192.165 2796.430 ;
        RECT 1200.230 455.755 1200.510 456.125 ;
        RECT 1200.300 435.725 1200.440 455.755 ;
        RECT 2318.030 437.395 2318.310 437.765 ;
        RECT 1828.130 436.715 1828.410 437.085 ;
        RECT 1414.130 436.035 1414.410 436.405 ;
        RECT 1463.810 436.035 1464.090 436.405 ;
        RECT 1634.930 436.035 1635.210 436.405 ;
        RECT 1683.230 436.035 1683.510 436.405 ;
        RECT 1414.140 435.890 1414.400 436.035 ;
        RECT 1463.820 435.890 1464.080 436.035 ;
        RECT 1200.230 435.355 1200.510 435.725 ;
        RECT 1268.770 435.610 1269.050 435.725 ;
        RECT 1269.690 435.610 1269.970 435.725 ;
        RECT 1268.770 435.470 1269.970 435.610 ;
        RECT 1268.770 435.355 1269.050 435.470 ;
        RECT 1269.690 435.355 1269.970 435.470 ;
        RECT 1635.000 435.045 1635.140 436.035 ;
        RECT 1683.300 435.045 1683.440 436.035 ;
        RECT 1828.200 435.870 1828.340 436.715 ;
        RECT 2125.750 436.035 2126.030 436.405 ;
        RECT 2246.270 436.035 2246.550 436.405 ;
        RECT 1780.300 435.725 1780.560 435.870 ;
        RECT 1780.290 435.355 1780.570 435.725 ;
        RECT 1828.140 435.550 1828.400 435.870 ;
        RECT 2089.420 435.725 2089.680 435.870 ;
        RECT 2091.720 435.725 2091.980 435.870 ;
        RECT 1992.350 435.355 1992.630 435.725 ;
        RECT 1994.190 435.355 1994.470 435.725 ;
        RECT 2089.410 435.355 2089.690 435.725 ;
        RECT 2091.710 435.355 2091.990 435.725 ;
        RECT 1992.360 435.210 1992.620 435.355 ;
        RECT 1994.200 435.210 1994.460 435.355 ;
        RECT 1634.930 434.675 1635.210 435.045 ;
        RECT 1683.230 434.675 1683.510 435.045 ;
        RECT 2125.290 434.930 2125.570 435.045 ;
        RECT 2125.820 434.930 2125.960 436.035 ;
        RECT 2246.340 435.190 2246.480 436.035 ;
        RECT 2318.100 435.725 2318.240 437.395 ;
        RECT 2318.030 435.355 2318.310 435.725 ;
        RECT 2221.900 435.045 2222.160 435.190 ;
        RECT 2125.290 434.790 2125.960 434.930 ;
        RECT 2125.290 434.675 2125.570 434.790 ;
        RECT 2221.890 434.675 2222.170 435.045 ;
        RECT 2246.280 434.870 2246.540 435.190 ;
        RECT 2318.960 435.045 2319.220 435.190 ;
        RECT 2332.760 435.045 2333.020 435.190 ;
        RECT 2318.950 434.675 2319.230 435.045 ;
        RECT 2332.750 434.675 2333.030 435.045 ;
      LAYER via2 ;
        RECT 1191.030 2796.360 1191.310 2796.640 ;
        RECT 1200.230 455.800 1200.510 456.080 ;
        RECT 2318.030 437.440 2318.310 437.720 ;
        RECT 1828.130 436.760 1828.410 437.040 ;
        RECT 1414.130 436.080 1414.410 436.360 ;
        RECT 1463.810 436.080 1464.090 436.360 ;
        RECT 1634.930 436.080 1635.210 436.360 ;
        RECT 1683.230 436.080 1683.510 436.360 ;
        RECT 1200.230 435.400 1200.510 435.680 ;
        RECT 1268.770 435.400 1269.050 435.680 ;
        RECT 1269.690 435.400 1269.970 435.680 ;
        RECT 2125.750 436.080 2126.030 436.360 ;
        RECT 2246.270 436.080 2246.550 436.360 ;
        RECT 1780.290 435.400 1780.570 435.680 ;
        RECT 1992.350 435.400 1992.630 435.680 ;
        RECT 1994.190 435.400 1994.470 435.680 ;
        RECT 2089.410 435.400 2089.690 435.680 ;
        RECT 2091.710 435.400 2091.990 435.680 ;
        RECT 1634.930 434.720 1635.210 435.000 ;
        RECT 1683.230 434.720 1683.510 435.000 ;
        RECT 2125.290 434.720 2125.570 435.000 ;
        RECT 2318.030 435.400 2318.310 435.680 ;
        RECT 2221.890 434.720 2222.170 435.000 ;
        RECT 2318.950 434.720 2319.230 435.000 ;
        RECT 2332.750 434.720 2333.030 435.000 ;
      LAYER met3 ;
        RECT 1191.005 2796.660 1191.335 2796.665 ;
        RECT 1190.750 2796.650 1191.335 2796.660 ;
        RECT 1190.550 2796.350 1191.335 2796.650 ;
        RECT 1190.750 2796.340 1191.335 2796.350 ;
        RECT 1191.005 2796.335 1191.335 2796.340 ;
        RECT 1190.750 456.090 1191.130 456.100 ;
        RECT 1200.205 456.090 1200.535 456.105 ;
        RECT 1190.750 455.790 1200.535 456.090 ;
        RECT 1190.750 455.780 1191.130 455.790 ;
        RECT 1200.205 455.775 1200.535 455.790 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 1497.110 437.730 1497.490 437.740 ;
        RECT 2269.910 437.730 2270.290 437.740 ;
        RECT 2318.005 437.730 2318.335 437.745 ;
        RECT 1497.110 437.430 1562.770 437.730 ;
        RECT 1497.110 437.420 1497.490 437.430 ;
        RECT 1345.310 436.370 1345.690 436.380 ;
        RECT 1414.105 436.370 1414.435 436.385 ;
        RECT 1272.670 436.070 1318.050 436.370 ;
        RECT 1200.205 435.690 1200.535 435.705 ;
        RECT 1268.745 435.690 1269.075 435.705 ;
        RECT 1200.205 435.390 1269.075 435.690 ;
        RECT 1200.205 435.375 1200.535 435.390 ;
        RECT 1268.745 435.375 1269.075 435.390 ;
        RECT 1269.665 435.690 1269.995 435.705 ;
        RECT 1272.670 435.690 1272.970 436.070 ;
        RECT 1269.665 435.390 1272.970 435.690 ;
        RECT 1269.665 435.375 1269.995 435.390 ;
        RECT 1317.750 435.010 1318.050 436.070 ;
        RECT 1345.310 436.070 1414.435 436.370 ;
        RECT 1345.310 436.060 1345.690 436.070 ;
        RECT 1414.105 436.055 1414.435 436.070 ;
        RECT 1463.785 436.370 1464.115 436.385 ;
        RECT 1497.110 436.370 1497.490 436.380 ;
        RECT 1463.785 436.070 1497.490 436.370 ;
        RECT 1562.470 436.370 1562.770 437.430 ;
        RECT 2269.910 437.430 2318.335 437.730 ;
        RECT 2269.910 437.420 2270.290 437.430 ;
        RECT 2318.005 437.415 2318.335 437.430 ;
        RECT 1828.105 437.050 1828.435 437.065 ;
        RECT 1834.750 437.050 1835.130 437.060 ;
        RECT 1828.105 436.750 1835.130 437.050 ;
        RECT 1828.105 436.735 1828.435 436.750 ;
        RECT 1834.750 436.740 1835.130 436.750 ;
        RECT 1896.430 436.750 1931.690 437.050 ;
        RECT 1587.270 436.370 1587.650 436.380 ;
        RECT 1562.470 436.070 1587.650 436.370 ;
        RECT 1463.785 436.055 1464.115 436.070 ;
        RECT 1497.110 436.060 1497.490 436.070 ;
        RECT 1587.270 436.060 1587.650 436.070 ;
        RECT 1634.905 436.370 1635.235 436.385 ;
        RECT 1683.205 436.370 1683.535 436.385 ;
        RECT 1634.905 436.070 1683.535 436.370 ;
        RECT 1634.905 436.055 1635.235 436.070 ;
        RECT 1683.205 436.055 1683.535 436.070 ;
        RECT 1780.265 435.690 1780.595 435.705 ;
        RECT 1896.430 435.690 1896.730 436.750 ;
        RECT 1702.310 435.390 1780.595 435.690 ;
        RECT 1345.310 435.010 1345.690 435.020 ;
        RECT 1317.750 434.710 1345.690 435.010 ;
        RECT 1345.310 434.700 1345.690 434.710 ;
        RECT 1587.270 435.010 1587.650 435.020 ;
        RECT 1634.905 435.010 1635.235 435.025 ;
        RECT 1587.270 434.710 1635.235 435.010 ;
        RECT 1587.270 434.700 1587.650 434.710 ;
        RECT 1634.905 434.695 1635.235 434.710 ;
        RECT 1683.205 435.010 1683.535 435.025 ;
        RECT 1702.310 435.010 1702.610 435.390 ;
        RECT 1780.265 435.375 1780.595 435.390 ;
        RECT 1849.510 435.390 1896.730 435.690 ;
        RECT 1683.205 434.710 1702.610 435.010 ;
        RECT 1834.750 435.010 1835.130 435.020 ;
        RECT 1849.510 435.010 1849.810 435.390 ;
        RECT 1834.750 434.710 1849.810 435.010 ;
        RECT 1931.390 435.010 1931.690 436.750 ;
        RECT 2125.725 436.370 2126.055 436.385 ;
        RECT 2246.245 436.370 2246.575 436.385 ;
        RECT 2269.910 436.370 2270.290 436.380 ;
        RECT 2125.725 436.070 2187.450 436.370 ;
        RECT 2125.725 436.055 2126.055 436.070 ;
        RECT 1992.325 435.690 1992.655 435.705 ;
        RECT 1946.110 435.390 1992.655 435.690 ;
        RECT 1946.110 435.010 1946.410 435.390 ;
        RECT 1992.325 435.375 1992.655 435.390 ;
        RECT 1994.165 435.690 1994.495 435.705 ;
        RECT 2089.385 435.690 2089.715 435.705 ;
        RECT 1994.165 435.390 2028.290 435.690 ;
        RECT 1994.165 435.375 1994.495 435.390 ;
        RECT 1931.390 434.710 1946.410 435.010 ;
        RECT 2027.990 435.010 2028.290 435.390 ;
        RECT 2042.710 435.390 2089.715 435.690 ;
        RECT 2042.710 435.010 2043.010 435.390 ;
        RECT 2089.385 435.375 2089.715 435.390 ;
        RECT 2091.685 435.690 2092.015 435.705 ;
        RECT 2091.685 435.390 2124.890 435.690 ;
        RECT 2091.685 435.375 2092.015 435.390 ;
        RECT 2027.990 434.710 2043.010 435.010 ;
        RECT 2124.590 435.010 2124.890 435.390 ;
        RECT 2125.265 435.010 2125.595 435.025 ;
        RECT 2124.590 434.710 2125.595 435.010 ;
        RECT 2187.150 435.010 2187.450 436.070 ;
        RECT 2246.245 436.070 2270.290 436.370 ;
        RECT 2246.245 436.055 2246.575 436.070 ;
        RECT 2269.910 436.060 2270.290 436.070 ;
        RECT 2366.510 436.370 2366.890 436.380 ;
        RECT 2366.510 436.070 2449.650 436.370 ;
        RECT 2366.510 436.060 2366.890 436.070 ;
        RECT 2318.005 435.690 2318.335 435.705 ;
        RECT 2449.350 435.690 2449.650 436.070 ;
        RECT 2498.110 436.070 2546.250 436.370 ;
        RECT 2318.005 435.390 2319.010 435.690 ;
        RECT 2449.350 435.390 2497.490 435.690 ;
        RECT 2318.005 435.375 2318.335 435.390 ;
        RECT 2318.710 435.025 2319.010 435.390 ;
        RECT 2221.865 435.010 2222.195 435.025 ;
        RECT 2187.150 434.710 2222.195 435.010 ;
        RECT 2318.710 434.710 2319.255 435.025 ;
        RECT 1683.205 434.695 1683.535 434.710 ;
        RECT 1834.750 434.700 1835.130 434.710 ;
        RECT 2125.265 434.695 2125.595 434.710 ;
        RECT 2221.865 434.695 2222.195 434.710 ;
        RECT 2318.925 434.695 2319.255 434.710 ;
        RECT 2332.725 435.010 2333.055 435.025 ;
        RECT 2366.510 435.010 2366.890 435.020 ;
        RECT 2332.725 434.710 2366.890 435.010 ;
        RECT 2497.190 435.010 2497.490 435.390 ;
        RECT 2498.110 435.010 2498.410 436.070 ;
        RECT 2545.950 435.690 2546.250 436.070 ;
        RECT 2594.710 436.070 2642.850 436.370 ;
        RECT 2545.950 435.390 2594.090 435.690 ;
        RECT 2497.190 434.710 2498.410 435.010 ;
        RECT 2593.790 435.010 2594.090 435.390 ;
        RECT 2594.710 435.010 2595.010 436.070 ;
        RECT 2642.550 435.690 2642.850 436.070 ;
        RECT 2691.310 436.070 2739.450 436.370 ;
        RECT 2642.550 435.390 2690.690 435.690 ;
        RECT 2593.790 434.710 2595.010 435.010 ;
        RECT 2690.390 435.010 2690.690 435.390 ;
        RECT 2691.310 435.010 2691.610 436.070 ;
        RECT 2739.150 435.690 2739.450 436.070 ;
        RECT 2787.910 436.070 2836.050 436.370 ;
        RECT 2739.150 435.390 2787.290 435.690 ;
        RECT 2690.390 434.710 2691.610 435.010 ;
        RECT 2786.990 435.010 2787.290 435.390 ;
        RECT 2787.910 435.010 2788.210 436.070 ;
        RECT 2835.750 435.690 2836.050 436.070 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2786.990 434.710 2788.210 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 2332.725 434.695 2333.055 434.710 ;
        RECT 2366.510 434.700 2366.890 434.710 ;
      LAYER via3 ;
        RECT 1190.780 2796.340 1191.100 2796.660 ;
        RECT 1190.780 455.780 1191.100 456.100 ;
        RECT 1497.140 437.420 1497.460 437.740 ;
        RECT 1345.340 436.060 1345.660 436.380 ;
        RECT 1497.140 436.060 1497.460 436.380 ;
        RECT 2269.940 437.420 2270.260 437.740 ;
        RECT 1834.780 436.740 1835.100 437.060 ;
        RECT 1587.300 436.060 1587.620 436.380 ;
        RECT 1345.340 434.700 1345.660 435.020 ;
        RECT 1587.300 434.700 1587.620 435.020 ;
        RECT 1834.780 434.700 1835.100 435.020 ;
        RECT 2269.940 436.060 2270.260 436.380 ;
        RECT 2366.540 436.060 2366.860 436.380 ;
        RECT 2366.540 434.700 2366.860 435.020 ;
      LAYER met4 ;
        RECT 1190.775 2796.335 1191.105 2796.665 ;
        RECT 1190.790 456.105 1191.090 2796.335 ;
        RECT 1190.775 455.775 1191.105 456.105 ;
        RECT 1497.135 437.415 1497.465 437.745 ;
        RECT 2269.935 437.415 2270.265 437.745 ;
        RECT 1497.150 436.385 1497.450 437.415 ;
        RECT 1834.775 436.735 1835.105 437.065 ;
        RECT 1345.335 436.055 1345.665 436.385 ;
        RECT 1497.135 436.055 1497.465 436.385 ;
        RECT 1587.295 436.055 1587.625 436.385 ;
        RECT 1345.350 435.025 1345.650 436.055 ;
        RECT 1587.310 435.025 1587.610 436.055 ;
        RECT 1834.790 435.025 1835.090 436.735 ;
        RECT 2269.950 436.385 2270.250 437.415 ;
        RECT 2269.935 436.055 2270.265 436.385 ;
        RECT 2366.535 436.055 2366.865 436.385 ;
        RECT 2366.550 435.025 2366.850 436.055 ;
        RECT 1345.335 434.695 1345.665 435.025 ;
        RECT 1587.295 434.695 1587.625 435.025 ;
        RECT 1834.775 434.695 1835.105 435.025 ;
        RECT 2366.535 434.695 2366.865 435.025 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3501.220 1014.230 3501.280 ;
        RECT 1739.330 3501.220 1739.650 3501.280 ;
        RECT 1013.910 3501.080 1739.650 3501.220 ;
        RECT 1013.910 3501.020 1014.230 3501.080 ;
        RECT 1739.330 3501.020 1739.650 3501.080 ;
      LAYER via ;
        RECT 1013.940 3501.020 1014.200 3501.280 ;
        RECT 1739.360 3501.020 1739.620 3501.280 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3501.310 1014.140 3517.600 ;
        RECT 1013.940 3500.990 1014.200 3501.310 ;
        RECT 1739.360 3500.990 1739.620 3501.310 ;
        RECT 1739.420 2799.970 1739.560 3500.990 ;
        RECT 1742.045 2799.970 1742.325 2800.000 ;
        RECT 1739.420 2799.830 1742.325 2799.970 ;
        RECT 1742.045 2796.000 1742.325 2799.830 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3503.600 689.470 3503.660 ;
        RECT 1766.470 3503.600 1766.790 3503.660 ;
        RECT 689.150 3503.460 1766.790 3503.600 ;
        RECT 689.150 3503.400 689.470 3503.460 ;
        RECT 1766.470 3503.400 1766.790 3503.460 ;
      LAYER via ;
        RECT 689.180 3503.400 689.440 3503.660 ;
        RECT 1766.500 3503.400 1766.760 3503.660 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.690 689.380 3517.600 ;
        RECT 689.180 3503.370 689.440 3503.690 ;
        RECT 1766.500 3503.370 1766.760 3503.690 ;
        RECT 1766.560 2800.650 1766.700 3503.370 ;
        RECT 1766.560 2800.510 1769.460 2800.650 ;
        RECT 1769.320 2799.970 1769.460 2800.510 ;
        RECT 1771.025 2799.970 1771.305 2800.000 ;
        RECT 1769.320 2799.830 1771.305 2799.970 ;
        RECT 1771.025 2796.000 1771.305 2799.830 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.240 365.170 3502.300 ;
        RECT 1794.070 3502.240 1794.390 3502.300 ;
        RECT 364.850 3502.100 1794.390 3502.240 ;
        RECT 364.850 3502.040 365.170 3502.100 ;
        RECT 1794.070 3502.040 1794.390 3502.100 ;
      LAYER via ;
        RECT 364.880 3502.040 365.140 3502.300 ;
        RECT 1794.100 3502.040 1794.360 3502.300 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 1794.100 3502.010 1794.360 3502.330 ;
        RECT 1794.160 2800.650 1794.300 3502.010 ;
        RECT 1794.160 2800.510 1798.900 2800.650 ;
        RECT 1798.760 2799.970 1798.900 2800.510 ;
        RECT 1800.005 2799.970 1800.285 2800.000 ;
        RECT 1798.760 2799.830 1800.285 2799.970 ;
        RECT 1800.005 2796.000 1800.285 2799.830 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 1828.590 3501.475 1828.870 3501.845 ;
        RECT 1828.660 2799.970 1828.800 3501.475 ;
        RECT 1828.985 2799.970 1829.265 2800.000 ;
        RECT 1828.660 2799.830 1829.265 2799.970 ;
        RECT 1828.985 2796.000 1829.265 2799.830 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 1828.590 3501.520 1828.870 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 1828.565 3501.810 1828.895 3501.825 ;
        RECT 40.545 3501.510 1828.895 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 1828.565 3501.495 1828.895 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1856.170 3263.900 1856.490 3263.960 ;
        RECT 15.250 3263.760 1856.490 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1856.170 3263.700 1856.490 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1856.200 3263.700 1856.460 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1856.200 3263.670 1856.460 3263.990 ;
        RECT 1856.260 2799.970 1856.400 3263.670 ;
        RECT 1857.965 2799.970 1858.245 2800.000 ;
        RECT 1856.260 2799.830 1858.245 2799.970 ;
        RECT 1857.965 2796.000 1858.245 2799.830 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 1883.770 2974.220 1884.090 2974.280 ;
        RECT 16.170 2974.080 1884.090 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 1883.770 2974.020 1884.090 2974.080 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 1883.800 2974.020 1884.060 2974.280 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 1883.800 2973.990 1884.060 2974.310 ;
        RECT 1883.860 2800.650 1884.000 2973.990 ;
        RECT 1883.860 2800.510 1885.380 2800.650 ;
        RECT 1885.240 2799.970 1885.380 2800.510 ;
        RECT 1886.945 2799.970 1887.225 2800.000 ;
        RECT 1885.240 2799.830 1887.225 2799.970 ;
        RECT 1886.945 2796.000 1887.225 2799.830 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1915.465 2796.570 1915.745 2800.000 ;
        RECT 1915.990 2796.570 1916.270 2796.685 ;
        RECT 1915.465 2796.430 1916.270 2796.570 ;
        RECT 1915.465 2796.000 1915.745 2796.430 ;
        RECT 1915.990 2796.315 1916.270 2796.430 ;
        RECT 14.810 2790.875 15.090 2791.245 ;
        RECT 14.880 2693.325 15.020 2790.875 ;
        RECT 14.810 2692.955 15.090 2693.325 ;
      LAYER via2 ;
        RECT 1915.990 2796.360 1916.270 2796.640 ;
        RECT 14.810 2790.920 15.090 2791.200 ;
        RECT 14.810 2693.000 15.090 2693.280 ;
      LAYER met3 ;
        RECT 1915.965 2796.660 1916.295 2796.665 ;
        RECT 1915.710 2796.650 1916.295 2796.660 ;
        RECT 1915.510 2796.350 1916.295 2796.650 ;
        RECT 1915.710 2796.340 1916.295 2796.350 ;
        RECT 1915.965 2796.335 1916.295 2796.340 ;
        RECT 14.785 2791.210 15.115 2791.225 ;
        RECT 1915.710 2791.210 1916.090 2791.220 ;
        RECT 14.785 2790.910 1916.090 2791.210 ;
        RECT 14.785 2790.895 15.115 2790.910 ;
        RECT 1915.710 2790.900 1916.090 2790.910 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 14.785 2693.290 15.115 2693.305 ;
        RECT -4.800 2692.990 15.115 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 14.785 2692.975 15.115 2692.990 ;
      LAYER via3 ;
        RECT 1915.740 2796.340 1916.060 2796.660 ;
        RECT 1915.740 2790.900 1916.060 2791.220 ;
      LAYER met4 ;
        RECT 1915.735 2796.335 1916.065 2796.665 ;
        RECT 1915.750 2791.225 1916.050 2796.335 ;
        RECT 1915.735 2790.895 1916.065 2791.225 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 32.730 2812.040 33.050 2812.100 ;
        RECT 1944.490 2812.040 1944.810 2812.100 ;
        RECT 32.730 2811.900 1944.810 2812.040 ;
        RECT 32.730 2811.840 33.050 2811.900 ;
        RECT 1944.490 2811.840 1944.810 2811.900 ;
        RECT 15.250 2405.740 15.570 2405.800 ;
        RECT 32.730 2405.740 33.050 2405.800 ;
        RECT 15.250 2405.600 33.050 2405.740 ;
        RECT 15.250 2405.540 15.570 2405.600 ;
        RECT 32.730 2405.540 33.050 2405.600 ;
      LAYER via ;
        RECT 32.760 2811.840 33.020 2812.100 ;
        RECT 1944.520 2811.840 1944.780 2812.100 ;
        RECT 15.280 2405.540 15.540 2405.800 ;
        RECT 32.760 2405.540 33.020 2405.800 ;
      LAYER met2 ;
        RECT 32.760 2811.810 33.020 2812.130 ;
        RECT 1944.520 2811.810 1944.780 2812.130 ;
        RECT 32.820 2405.830 32.960 2811.810 ;
        RECT 1944.580 2800.000 1944.720 2811.810 ;
        RECT 1944.445 2796.000 1944.725 2800.000 ;
        RECT 15.280 2405.685 15.540 2405.830 ;
        RECT 15.270 2405.315 15.550 2405.685 ;
        RECT 32.760 2405.510 33.020 2405.830 ;
      LAYER via2 ;
        RECT 15.270 2405.360 15.550 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.245 2405.650 15.575 2405.665 ;
        RECT -4.800 2405.350 15.575 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.245 2405.335 15.575 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 27.210 2810.680 27.530 2810.740 ;
        RECT 1973.470 2810.680 1973.790 2810.740 ;
        RECT 27.210 2810.540 1973.790 2810.680 ;
        RECT 27.210 2810.480 27.530 2810.540 ;
        RECT 1973.470 2810.480 1973.790 2810.540 ;
        RECT 13.870 2123.540 14.190 2123.600 ;
        RECT 27.210 2123.540 27.530 2123.600 ;
        RECT 13.870 2123.400 27.530 2123.540 ;
        RECT 13.870 2123.340 14.190 2123.400 ;
        RECT 27.210 2123.340 27.530 2123.400 ;
      LAYER via ;
        RECT 27.240 2810.480 27.500 2810.740 ;
        RECT 1973.500 2810.480 1973.760 2810.740 ;
        RECT 13.900 2123.340 14.160 2123.600 ;
        RECT 27.240 2123.340 27.500 2123.600 ;
      LAYER met2 ;
        RECT 27.240 2810.450 27.500 2810.770 ;
        RECT 1973.500 2810.450 1973.760 2810.770 ;
        RECT 27.300 2123.630 27.440 2810.450 ;
        RECT 1973.560 2800.000 1973.700 2810.450 ;
        RECT 1973.425 2796.000 1973.705 2800.000 ;
        RECT 13.900 2123.310 14.160 2123.630 ;
        RECT 27.240 2123.310 27.500 2123.630 ;
        RECT 13.960 2118.725 14.100 2123.310 ;
        RECT 13.890 2118.355 14.170 2118.725 ;
      LAYER via2 ;
        RECT 13.890 2118.400 14.170 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 13.865 2118.690 14.195 2118.705 ;
        RECT -4.800 2118.390 14.195 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 13.865 2118.375 14.195 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 2809.660 27.070 2809.720 ;
        RECT 2002.450 2809.660 2002.770 2809.720 ;
        RECT 26.750 2809.520 2002.770 2809.660 ;
        RECT 26.750 2809.460 27.070 2809.520 ;
        RECT 2002.450 2809.460 2002.770 2809.520 ;
        RECT 13.870 1834.880 14.190 1834.940 ;
        RECT 26.750 1834.880 27.070 1834.940 ;
        RECT 13.870 1834.740 27.070 1834.880 ;
        RECT 13.870 1834.680 14.190 1834.740 ;
        RECT 26.750 1834.680 27.070 1834.740 ;
      LAYER via ;
        RECT 26.780 2809.460 27.040 2809.720 ;
        RECT 2002.480 2809.460 2002.740 2809.720 ;
        RECT 13.900 1834.680 14.160 1834.940 ;
        RECT 26.780 1834.680 27.040 1834.940 ;
      LAYER met2 ;
        RECT 26.780 2809.430 27.040 2809.750 ;
        RECT 2002.480 2809.430 2002.740 2809.750 ;
        RECT 26.840 1834.970 26.980 2809.430 ;
        RECT 2002.540 2800.000 2002.680 2809.430 ;
        RECT 2002.405 2796.000 2002.685 2800.000 ;
        RECT 13.900 1834.650 14.160 1834.970 ;
        RECT 26.780 1834.650 27.040 1834.970 ;
        RECT 13.960 1831.085 14.100 1834.650 ;
        RECT 13.890 1830.715 14.170 1831.085 ;
      LAYER via2 ;
        RECT 13.890 1830.760 14.170 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 13.865 1831.050 14.195 1831.065 ;
        RECT -4.800 1830.750 14.195 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 13.865 1830.735 14.195 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.570 670.720 1345.890 670.780 ;
        RECT 1376.850 670.720 1377.170 670.780 ;
        RECT 1345.570 670.580 1377.170 670.720 ;
        RECT 1345.570 670.520 1345.890 670.580 ;
        RECT 1376.850 670.520 1377.170 670.580 ;
        RECT 1787.170 670.380 1787.490 670.440 ;
        RECT 1805.570 670.380 1805.890 670.440 ;
        RECT 1787.170 670.240 1805.890 670.380 ;
        RECT 1787.170 670.180 1787.490 670.240 ;
        RECT 1805.570 670.180 1805.890 670.240 ;
        RECT 1992.330 670.380 1992.650 670.440 ;
        RECT 1995.090 670.380 1995.410 670.440 ;
        RECT 1992.330 670.240 1995.410 670.380 ;
        RECT 1992.330 670.180 1992.650 670.240 ;
        RECT 1995.090 670.180 1995.410 670.240 ;
        RECT 2089.390 670.380 2089.710 670.440 ;
        RECT 2091.690 670.380 2092.010 670.440 ;
        RECT 2089.390 670.240 2092.010 670.380 ;
        RECT 2089.390 670.180 2089.710 670.240 ;
        RECT 2091.690 670.180 2092.010 670.240 ;
        RECT 1587.530 670.040 1587.850 670.100 ;
        RECT 1634.450 670.040 1634.770 670.100 ;
        RECT 1587.530 669.900 1634.770 670.040 ;
        RECT 1587.530 669.840 1587.850 669.900 ;
        RECT 1634.450 669.840 1634.770 669.900 ;
        RECT 1255.870 669.700 1256.190 669.760 ;
        RECT 1303.710 669.700 1304.030 669.760 ;
        RECT 1255.870 669.560 1304.030 669.700 ;
        RECT 1255.870 669.500 1256.190 669.560 ;
        RECT 1303.710 669.500 1304.030 669.560 ;
        RECT 1636.290 669.700 1636.610 669.760 ;
        RECT 1683.210 669.700 1683.530 669.760 ;
        RECT 1636.290 669.560 1683.530 669.700 ;
        RECT 1636.290 669.500 1636.610 669.560 ;
        RECT 1683.210 669.500 1683.530 669.560 ;
      LAYER via ;
        RECT 1345.600 670.520 1345.860 670.780 ;
        RECT 1376.880 670.520 1377.140 670.780 ;
        RECT 1787.200 670.180 1787.460 670.440 ;
        RECT 1805.600 670.180 1805.860 670.440 ;
        RECT 1992.360 670.180 1992.620 670.440 ;
        RECT 1995.120 670.180 1995.380 670.440 ;
        RECT 2089.420 670.180 2089.680 670.440 ;
        RECT 2091.720 670.180 2091.980 670.440 ;
        RECT 1587.560 669.840 1587.820 670.100 ;
        RECT 1634.480 669.840 1634.740 670.100 ;
        RECT 1255.900 669.500 1256.160 669.760 ;
        RECT 1303.740 669.500 1304.000 669.760 ;
        RECT 1636.320 669.500 1636.580 669.760 ;
        RECT 1683.240 669.500 1683.500 669.760 ;
      LAYER met2 ;
        RECT 1219.090 2811.955 1219.370 2812.325 ;
        RECT 1219.160 2799.970 1219.300 2811.955 ;
        RECT 1220.865 2799.970 1221.145 2800.000 ;
        RECT 1219.160 2799.830 1221.145 2799.970 ;
        RECT 1220.865 2796.000 1221.145 2799.830 ;
        RECT 2304.230 672.675 2304.510 673.045 ;
        RECT 2236.150 671.315 2236.430 671.685 ;
        RECT 1303.730 670.635 1304.010 671.005 ;
        RECT 1345.590 670.635 1345.870 671.005 ;
        RECT 1303.800 669.790 1303.940 670.635 ;
        RECT 1345.600 670.490 1345.860 670.635 ;
        RECT 1376.880 670.490 1377.140 670.810 ;
        RECT 1683.230 670.635 1683.510 671.005 ;
        RECT 1376.940 670.325 1377.080 670.490 ;
        RECT 1376.870 669.955 1377.150 670.325 ;
        RECT 1413.670 670.210 1413.950 670.325 ;
        RECT 1414.590 670.210 1414.870 670.325 ;
        RECT 1413.670 670.070 1414.870 670.210 ;
        RECT 1413.670 669.955 1413.950 670.070 ;
        RECT 1414.590 669.955 1414.870 670.070 ;
        RECT 1545.230 669.955 1545.510 670.325 ;
        RECT 1587.550 669.955 1587.830 670.325 ;
        RECT 1255.900 669.645 1256.160 669.790 ;
        RECT 1255.890 669.275 1256.170 669.645 ;
        RECT 1303.740 669.470 1304.000 669.790 ;
        RECT 1545.300 668.965 1545.440 669.955 ;
        RECT 1587.560 669.810 1587.820 669.955 ;
        RECT 1634.480 669.810 1634.740 670.130 ;
        RECT 1634.540 669.530 1634.680 669.810 ;
        RECT 1683.300 669.790 1683.440 670.635 ;
        RECT 1787.200 670.325 1787.460 670.470 ;
        RECT 1805.600 670.325 1805.860 670.470 ;
        RECT 1992.360 670.325 1992.620 670.470 ;
        RECT 1995.120 670.325 1995.380 670.470 ;
        RECT 2089.420 670.325 2089.680 670.470 ;
        RECT 2091.720 670.325 2091.980 670.470 ;
        RECT 1787.190 669.955 1787.470 670.325 ;
        RECT 1805.590 669.955 1805.870 670.325 ;
        RECT 1992.350 669.955 1992.630 670.325 ;
        RECT 1995.110 669.955 1995.390 670.325 ;
        RECT 2089.410 669.955 2089.690 670.325 ;
        RECT 2091.710 669.955 2091.990 670.325 ;
        RECT 2235.690 670.210 2235.970 670.325 ;
        RECT 2236.220 670.210 2236.360 671.315 ;
        RECT 2304.300 671.005 2304.440 672.675 ;
        RECT 2304.230 670.635 2304.510 671.005 ;
        RECT 2235.690 670.070 2236.360 670.210 ;
        RECT 2235.690 669.955 2235.970 670.070 ;
        RECT 1636.320 669.645 1636.580 669.790 ;
        RECT 1634.930 669.530 1635.210 669.645 ;
        RECT 1634.540 669.390 1635.210 669.530 ;
        RECT 1634.930 669.275 1635.210 669.390 ;
        RECT 1636.310 669.275 1636.590 669.645 ;
        RECT 1683.240 669.470 1683.500 669.790 ;
        RECT 1545.230 668.595 1545.510 668.965 ;
      LAYER via2 ;
        RECT 1219.090 2812.000 1219.370 2812.280 ;
        RECT 2304.230 672.720 2304.510 673.000 ;
        RECT 2236.150 671.360 2236.430 671.640 ;
        RECT 1303.730 670.680 1304.010 670.960 ;
        RECT 1345.590 670.680 1345.870 670.960 ;
        RECT 1683.230 670.680 1683.510 670.960 ;
        RECT 1376.870 670.000 1377.150 670.280 ;
        RECT 1413.670 670.000 1413.950 670.280 ;
        RECT 1414.590 670.000 1414.870 670.280 ;
        RECT 1545.230 670.000 1545.510 670.280 ;
        RECT 1587.550 670.000 1587.830 670.280 ;
        RECT 1255.890 669.320 1256.170 669.600 ;
        RECT 1787.190 670.000 1787.470 670.280 ;
        RECT 1805.590 670.000 1805.870 670.280 ;
        RECT 1992.350 670.000 1992.630 670.280 ;
        RECT 1995.110 670.000 1995.390 670.280 ;
        RECT 2089.410 670.000 2089.690 670.280 ;
        RECT 2091.710 670.000 2091.990 670.280 ;
        RECT 2235.690 670.000 2235.970 670.280 ;
        RECT 2304.230 670.680 2304.510 670.960 ;
        RECT 1634.930 669.320 1635.210 669.600 ;
        RECT 1636.310 669.320 1636.590 669.600 ;
        RECT 1545.230 668.640 1545.510 668.920 ;
      LAYER met3 ;
        RECT 1189.830 2812.290 1190.210 2812.300 ;
        RECT 1219.065 2812.290 1219.395 2812.305 ;
        RECT 1189.830 2811.990 1219.395 2812.290 ;
        RECT 1189.830 2811.980 1190.210 2811.990 ;
        RECT 1219.065 2811.975 1219.395 2811.990 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2916.710 674.070 2924.800 674.370 ;
        RECT 2269.910 673.010 2270.290 673.020 ;
        RECT 2304.205 673.010 2304.535 673.025 ;
        RECT 2269.910 672.710 2304.535 673.010 ;
        RECT 2269.910 672.700 2270.290 672.710 ;
        RECT 2304.205 672.695 2304.535 672.710 ;
        RECT 2236.125 671.650 2236.455 671.665 ;
        RECT 2269.910 671.650 2270.290 671.660 ;
        RECT 1883.550 671.350 1931.690 671.650 ;
        RECT 1303.705 670.970 1304.035 670.985 ;
        RECT 1345.565 670.970 1345.895 670.985 ;
        RECT 1303.705 670.670 1345.895 670.970 ;
        RECT 1303.705 670.655 1304.035 670.670 ;
        RECT 1345.565 670.655 1345.895 670.670 ;
        RECT 1683.205 670.970 1683.535 670.985 ;
        RECT 1683.205 670.670 1702.610 670.970 ;
        RECT 1683.205 670.655 1683.535 670.670 ;
        RECT 1376.845 670.290 1377.175 670.305 ;
        RECT 1413.645 670.290 1413.975 670.305 ;
        RECT 1376.845 669.990 1413.975 670.290 ;
        RECT 1376.845 669.975 1377.175 669.990 ;
        RECT 1413.645 669.975 1413.975 669.990 ;
        RECT 1414.565 670.290 1414.895 670.305 ;
        RECT 1545.205 670.290 1545.535 670.305 ;
        RECT 1587.525 670.290 1587.855 670.305 ;
        RECT 1414.565 669.990 1418.330 670.290 ;
        RECT 1414.565 669.975 1414.895 669.990 ;
        RECT 1189.830 669.610 1190.210 669.620 ;
        RECT 1255.865 669.610 1256.195 669.625 ;
        RECT 1189.830 669.310 1256.195 669.610 ;
        RECT 1418.030 669.610 1418.330 669.990 ;
        RECT 1545.205 669.990 1587.855 670.290 ;
        RECT 1545.205 669.975 1545.535 669.990 ;
        RECT 1587.525 669.975 1587.855 669.990 ;
        RECT 1634.905 669.610 1635.235 669.625 ;
        RECT 1636.285 669.610 1636.615 669.625 ;
        RECT 1418.030 669.310 1449.610 669.610 ;
        RECT 1189.830 669.300 1190.210 669.310 ;
        RECT 1255.865 669.295 1256.195 669.310 ;
        RECT 1449.310 668.930 1449.610 669.310 ;
        RECT 1634.905 669.310 1636.615 669.610 ;
        RECT 1702.310 669.610 1702.610 670.670 ;
        RECT 1787.165 670.290 1787.495 670.305 ;
        RECT 1752.910 669.990 1787.495 670.290 ;
        RECT 1752.910 669.610 1753.210 669.990 ;
        RECT 1787.165 669.975 1787.495 669.990 ;
        RECT 1805.565 670.290 1805.895 670.305 ;
        RECT 1883.550 670.290 1883.850 671.350 ;
        RECT 1805.565 669.990 1835.090 670.290 ;
        RECT 1805.565 669.975 1805.895 669.990 ;
        RECT 1702.310 669.310 1753.210 669.610 ;
        RECT 1834.790 669.610 1835.090 669.990 ;
        RECT 1849.510 669.990 1883.850 670.290 ;
        RECT 1849.510 669.610 1849.810 669.990 ;
        RECT 1834.790 669.310 1849.810 669.610 ;
        RECT 1931.390 669.610 1931.690 671.350 ;
        RECT 2236.125 671.350 2270.290 671.650 ;
        RECT 2236.125 671.335 2236.455 671.350 ;
        RECT 2269.910 671.340 2270.290 671.350 ;
        RECT 2304.205 670.970 2304.535 670.985 ;
        RECT 2304.205 670.670 2353.050 670.970 ;
        RECT 2304.205 670.655 2304.535 670.670 ;
        RECT 1992.325 670.290 1992.655 670.305 ;
        RECT 1946.110 669.990 1992.655 670.290 ;
        RECT 1946.110 669.610 1946.410 669.990 ;
        RECT 1992.325 669.975 1992.655 669.990 ;
        RECT 1995.085 670.290 1995.415 670.305 ;
        RECT 2089.385 670.290 2089.715 670.305 ;
        RECT 1995.085 669.990 2028.290 670.290 ;
        RECT 1995.085 669.975 1995.415 669.990 ;
        RECT 1931.390 669.310 1946.410 669.610 ;
        RECT 2027.990 669.610 2028.290 669.990 ;
        RECT 2042.710 669.990 2089.715 670.290 ;
        RECT 2042.710 669.610 2043.010 669.990 ;
        RECT 2089.385 669.975 2089.715 669.990 ;
        RECT 2091.685 670.290 2092.015 670.305 ;
        RECT 2235.665 670.290 2235.995 670.305 ;
        RECT 2091.685 669.990 2124.890 670.290 ;
        RECT 2091.685 669.975 2092.015 669.990 ;
        RECT 2027.990 669.310 2043.010 669.610 ;
        RECT 2124.590 669.610 2124.890 669.990 ;
        RECT 2139.310 669.990 2235.995 670.290 ;
        RECT 2352.750 670.290 2353.050 670.670 ;
        RECT 2401.510 670.670 2449.650 670.970 ;
        RECT 2352.750 669.990 2400.890 670.290 ;
        RECT 2139.310 669.610 2139.610 669.990 ;
        RECT 2235.665 669.975 2235.995 669.990 ;
        RECT 2124.590 669.310 2139.610 669.610 ;
        RECT 2400.590 669.610 2400.890 669.990 ;
        RECT 2401.510 669.610 2401.810 670.670 ;
        RECT 2449.350 670.290 2449.650 670.670 ;
        RECT 2498.110 670.670 2546.250 670.970 ;
        RECT 2449.350 669.990 2497.490 670.290 ;
        RECT 2400.590 669.310 2401.810 669.610 ;
        RECT 2497.190 669.610 2497.490 669.990 ;
        RECT 2498.110 669.610 2498.410 670.670 ;
        RECT 2545.950 670.290 2546.250 670.670 ;
        RECT 2594.710 670.670 2642.850 670.970 ;
        RECT 2545.950 669.990 2594.090 670.290 ;
        RECT 2497.190 669.310 2498.410 669.610 ;
        RECT 2593.790 669.610 2594.090 669.990 ;
        RECT 2594.710 669.610 2595.010 670.670 ;
        RECT 2642.550 670.290 2642.850 670.670 ;
        RECT 2691.310 670.670 2739.450 670.970 ;
        RECT 2642.550 669.990 2690.690 670.290 ;
        RECT 2593.790 669.310 2595.010 669.610 ;
        RECT 2690.390 669.610 2690.690 669.990 ;
        RECT 2691.310 669.610 2691.610 670.670 ;
        RECT 2739.150 670.290 2739.450 670.670 ;
        RECT 2787.910 670.670 2836.050 670.970 ;
        RECT 2739.150 669.990 2787.290 670.290 ;
        RECT 2690.390 669.310 2691.610 669.610 ;
        RECT 2786.990 669.610 2787.290 669.990 ;
        RECT 2787.910 669.610 2788.210 670.670 ;
        RECT 2835.750 670.290 2836.050 670.670 ;
        RECT 2916.710 670.290 2917.010 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
        RECT 2835.750 669.990 2883.890 670.290 ;
        RECT 2786.990 669.310 2788.210 669.610 ;
        RECT 2883.590 669.610 2883.890 669.990 ;
        RECT 2884.510 669.990 2917.010 670.290 ;
        RECT 2884.510 669.610 2884.810 669.990 ;
        RECT 2883.590 669.310 2884.810 669.610 ;
        RECT 1634.905 669.295 1635.235 669.310 ;
        RECT 1636.285 669.295 1636.615 669.310 ;
        RECT 1545.205 668.930 1545.535 668.945 ;
        RECT 1449.310 668.630 1545.535 668.930 ;
        RECT 1545.205 668.615 1545.535 668.630 ;
      LAYER via3 ;
        RECT 1189.860 2811.980 1190.180 2812.300 ;
        RECT 2269.940 672.700 2270.260 673.020 ;
        RECT 1189.860 669.300 1190.180 669.620 ;
        RECT 2269.940 671.340 2270.260 671.660 ;
      LAYER met4 ;
        RECT 1189.855 2811.975 1190.185 2812.305 ;
        RECT 1189.870 669.625 1190.170 2811.975 ;
        RECT 2269.935 672.695 2270.265 673.025 ;
        RECT 2269.950 671.665 2270.250 672.695 ;
        RECT 2269.935 671.335 2270.265 671.665 ;
        RECT 1189.855 669.295 1190.185 669.625 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1243.910 2798.100 1244.230 2798.160 ;
        RECT 1200.760 2797.960 1244.230 2798.100 ;
        RECT 1200.760 2797.480 1200.900 2797.960 ;
        RECT 1243.910 2797.900 1244.230 2797.960 ;
        RECT 1200.670 2797.220 1200.990 2797.480 ;
      LAYER via ;
        RECT 1243.940 2797.900 1244.200 2798.160 ;
        RECT 1200.700 2797.220 1200.960 2797.480 ;
      LAYER met2 ;
        RECT 1457.830 2799.035 1458.110 2799.405 ;
        RECT 1483.130 2799.035 1483.410 2799.405 ;
        RECT 1521.310 2799.035 1521.590 2799.405 ;
        RECT 1243.940 2797.870 1244.200 2798.190 ;
        RECT 1200.700 2797.365 1200.960 2797.510 ;
        RECT 1200.690 2796.995 1200.970 2797.365 ;
        RECT 1244.000 2796.685 1244.140 2797.870 ;
        RECT 1263.250 2797.675 1263.530 2798.045 ;
        RECT 1386.530 2797.675 1386.810 2798.045 ;
        RECT 1243.930 2796.315 1244.210 2796.685 ;
        RECT 1262.790 2796.570 1263.070 2796.685 ;
        RECT 1263.320 2796.570 1263.460 2797.675 ;
        RECT 1386.600 2796.685 1386.740 2797.675 ;
        RECT 1457.900 2796.685 1458.040 2799.035 ;
        RECT 1483.200 2798.045 1483.340 2799.035 ;
        RECT 1483.130 2797.675 1483.410 2798.045 ;
        RECT 1521.380 2797.365 1521.520 2799.035 ;
        RECT 1970.270 2797.675 1970.550 2798.045 ;
        RECT 2029.610 2797.930 2029.890 2798.045 ;
        RECT 2031.385 2797.930 2031.665 2800.000 ;
        RECT 2029.610 2797.790 2031.665 2797.930 ;
        RECT 2029.610 2797.675 2029.890 2797.790 ;
        RECT 1521.310 2796.995 1521.590 2797.365 ;
        RECT 1806.580 2797.110 1807.640 2797.250 ;
        RECT 1806.580 2796.685 1806.720 2797.110 ;
        RECT 1807.500 2796.685 1807.640 2797.110 ;
        RECT 1970.340 2796.685 1970.480 2797.675 ;
        RECT 1262.790 2796.430 1263.460 2796.570 ;
        RECT 1262.790 2796.315 1263.070 2796.430 ;
        RECT 1386.530 2796.315 1386.810 2796.685 ;
        RECT 1457.830 2796.315 1458.110 2796.685 ;
        RECT 1806.510 2796.315 1806.790 2796.685 ;
        RECT 1807.430 2796.315 1807.710 2796.685 ;
        RECT 1970.270 2796.315 1970.550 2796.685 ;
        RECT 2031.385 2796.000 2031.665 2797.790 ;
      LAYER via2 ;
        RECT 1457.830 2799.080 1458.110 2799.360 ;
        RECT 1483.130 2799.080 1483.410 2799.360 ;
        RECT 1521.310 2799.080 1521.590 2799.360 ;
        RECT 1200.690 2797.040 1200.970 2797.320 ;
        RECT 1263.250 2797.720 1263.530 2798.000 ;
        RECT 1386.530 2797.720 1386.810 2798.000 ;
        RECT 1243.930 2796.360 1244.210 2796.640 ;
        RECT 1262.790 2796.360 1263.070 2796.640 ;
        RECT 1483.130 2797.720 1483.410 2798.000 ;
        RECT 1970.270 2797.720 1970.550 2798.000 ;
        RECT 2029.610 2797.720 2029.890 2798.000 ;
        RECT 1521.310 2797.040 1521.590 2797.320 ;
        RECT 1386.530 2796.360 1386.810 2796.640 ;
        RECT 1457.830 2796.360 1458.110 2796.640 ;
        RECT 1806.510 2796.360 1806.790 2796.640 ;
        RECT 1807.430 2796.360 1807.710 2796.640 ;
        RECT 1970.270 2796.360 1970.550 2796.640 ;
      LAYER met3 ;
        RECT 1457.805 2799.370 1458.135 2799.385 ;
        RECT 1483.105 2799.370 1483.435 2799.385 ;
        RECT 1457.805 2799.070 1483.435 2799.370 ;
        RECT 1457.805 2799.055 1458.135 2799.070 ;
        RECT 1483.105 2799.055 1483.435 2799.070 ;
        RECT 1497.110 2799.370 1497.490 2799.380 ;
        RECT 1521.285 2799.370 1521.615 2799.385 ;
        RECT 1497.110 2799.070 1521.615 2799.370 ;
        RECT 1497.110 2799.060 1497.490 2799.070 ;
        RECT 1521.285 2799.055 1521.615 2799.070 ;
        RECT 1263.225 2798.010 1263.555 2798.025 ;
        RECT 1386.505 2798.010 1386.835 2798.025 ;
        RECT 1263.225 2797.710 1386.835 2798.010 ;
        RECT 1263.225 2797.695 1263.555 2797.710 ;
        RECT 1386.505 2797.695 1386.835 2797.710 ;
        RECT 1483.105 2798.010 1483.435 2798.025 ;
        RECT 1497.110 2798.010 1497.490 2798.020 ;
        RECT 1483.105 2797.710 1497.490 2798.010 ;
        RECT 1483.105 2797.695 1483.435 2797.710 ;
        RECT 1497.110 2797.700 1497.490 2797.710 ;
        RECT 1970.245 2798.010 1970.575 2798.025 ;
        RECT 2029.585 2798.010 2029.915 2798.025 ;
        RECT 1970.245 2797.710 2029.915 2798.010 ;
        RECT 1970.245 2797.695 1970.575 2797.710 ;
        RECT 2029.585 2797.695 2029.915 2797.710 ;
        RECT 1183.390 2797.330 1183.770 2797.340 ;
        RECT 1200.665 2797.330 1200.995 2797.345 ;
        RECT 1183.390 2797.030 1200.995 2797.330 ;
        RECT 1183.390 2797.020 1183.770 2797.030 ;
        RECT 1200.665 2797.015 1200.995 2797.030 ;
        RECT 1521.285 2797.330 1521.615 2797.345 ;
        RECT 1538.510 2797.330 1538.890 2797.340 ;
        RECT 1521.285 2797.030 1538.890 2797.330 ;
        RECT 1521.285 2797.015 1521.615 2797.030 ;
        RECT 1538.510 2797.020 1538.890 2797.030 ;
        RECT 1608.470 2797.030 1680.530 2797.330 ;
        RECT 1243.905 2796.650 1244.235 2796.665 ;
        RECT 1262.765 2796.650 1263.095 2796.665 ;
        RECT 1243.905 2796.350 1263.095 2796.650 ;
        RECT 1243.905 2796.335 1244.235 2796.350 ;
        RECT 1262.765 2796.335 1263.095 2796.350 ;
        RECT 1386.505 2796.650 1386.835 2796.665 ;
        RECT 1457.805 2796.650 1458.135 2796.665 ;
        RECT 1386.505 2796.350 1458.135 2796.650 ;
        RECT 1386.505 2796.335 1386.835 2796.350 ;
        RECT 1457.805 2796.335 1458.135 2796.350 ;
        RECT 1539.430 2796.650 1539.810 2796.660 ;
        RECT 1608.470 2796.650 1608.770 2797.030 ;
        RECT 1539.430 2796.350 1608.770 2796.650 ;
        RECT 1680.230 2796.650 1680.530 2797.030 ;
        RECT 1850.430 2797.030 1916.970 2797.330 ;
        RECT 1806.485 2796.650 1806.815 2796.665 ;
        RECT 1680.230 2796.350 1806.815 2796.650 ;
        RECT 1539.430 2796.340 1539.810 2796.350 ;
        RECT 1806.485 2796.335 1806.815 2796.350 ;
        RECT 1807.405 2796.650 1807.735 2796.665 ;
        RECT 1850.430 2796.650 1850.730 2797.030 ;
        RECT 1807.405 2796.350 1850.730 2796.650 ;
        RECT 1916.670 2796.650 1916.970 2797.030 ;
        RECT 1970.245 2796.650 1970.575 2796.665 ;
        RECT 1916.670 2796.350 1921.570 2796.650 ;
        RECT 1807.405 2796.335 1807.735 2796.350 ;
        RECT 1921.270 2795.970 1921.570 2796.350 ;
        RECT 1970.030 2796.335 1970.575 2796.650 ;
        RECT 1970.030 2795.970 1970.330 2796.335 ;
        RECT 1921.270 2795.670 1970.330 2795.970 ;
        RECT 1183.390 1545.450 1183.770 1545.460 ;
        RECT 3.070 1545.150 1183.770 1545.450 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 3.070 1544.090 3.370 1545.150 ;
        RECT 1183.390 1545.140 1183.770 1545.150 ;
        RECT -4.800 1543.790 3.370 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
      LAYER via3 ;
        RECT 1497.140 2799.060 1497.460 2799.380 ;
        RECT 1497.140 2797.700 1497.460 2798.020 ;
        RECT 1183.420 2797.020 1183.740 2797.340 ;
        RECT 1538.540 2797.020 1538.860 2797.340 ;
        RECT 1539.460 2796.340 1539.780 2796.660 ;
        RECT 1183.420 1545.140 1183.740 1545.460 ;
      LAYER met4 ;
        RECT 1497.135 2799.055 1497.465 2799.385 ;
        RECT 1497.150 2798.025 1497.450 2799.055 ;
        RECT 1497.135 2797.695 1497.465 2798.025 ;
        RECT 1183.415 2797.015 1183.745 2797.345 ;
        RECT 1538.535 2797.015 1538.865 2797.345 ;
        RECT 1183.430 1545.465 1183.730 2797.015 ;
        RECT 1538.550 2796.650 1538.850 2797.015 ;
        RECT 1539.455 2796.650 1539.785 2796.665 ;
        RECT 1538.550 2796.350 1539.785 2796.650 ;
        RECT 1539.455 2796.335 1539.785 2796.350 ;
        RECT 1183.415 1545.135 1183.745 1545.465 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1449.070 2815.100 1449.390 2815.160 ;
        RECT 2060.410 2815.100 2060.730 2815.160 ;
        RECT 1449.070 2814.960 1524.740 2815.100 ;
        RECT 1449.070 2814.900 1449.390 2814.960 ;
        RECT 1524.600 2814.760 1524.740 2814.960 ;
        RECT 1535.180 2814.960 2060.730 2815.100 ;
        RECT 1535.180 2814.760 1535.320 2814.960 ;
        RECT 2060.410 2814.900 2060.730 2814.960 ;
        RECT 1524.600 2814.620 1535.320 2814.760 ;
        RECT 20.310 2804.900 20.630 2804.960 ;
        RECT 1449.070 2804.900 1449.390 2804.960 ;
        RECT 20.310 2804.760 1449.390 2804.900 ;
        RECT 20.310 2804.700 20.630 2804.760 ;
        RECT 1449.070 2804.700 1449.390 2804.760 ;
      LAYER via ;
        RECT 1449.100 2814.900 1449.360 2815.160 ;
        RECT 2060.440 2814.900 2060.700 2815.160 ;
        RECT 20.340 2804.700 20.600 2804.960 ;
        RECT 1449.100 2804.700 1449.360 2804.960 ;
      LAYER met2 ;
        RECT 1449.100 2814.870 1449.360 2815.190 ;
        RECT 2060.440 2814.870 2060.700 2815.190 ;
        RECT 1449.160 2804.990 1449.300 2814.870 ;
        RECT 20.340 2804.670 20.600 2804.990 ;
        RECT 1449.100 2804.670 1449.360 2804.990 ;
        RECT 20.400 1328.565 20.540 2804.670 ;
        RECT 2060.500 2800.000 2060.640 2814.870 ;
        RECT 2060.365 2796.000 2060.645 2800.000 ;
        RECT 20.330 1328.195 20.610 1328.565 ;
      LAYER via2 ;
        RECT 20.330 1328.240 20.610 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 20.305 1328.530 20.635 1328.545 ;
        RECT -4.800 1328.230 20.635 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 20.305 1328.215 20.635 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1976.765 2805.085 1976.935 2810.695 ;
        RECT 1861.305 2798.625 1862.395 2798.795 ;
      LAYER mcon ;
        RECT 1976.765 2810.525 1976.935 2810.695 ;
        RECT 1862.225 2798.625 1862.395 2798.795 ;
      LAYER met1 ;
        RECT 1976.705 2810.680 1976.995 2810.725 ;
        RECT 2089.390 2810.680 2089.710 2810.740 ;
        RECT 1976.705 2810.540 2089.710 2810.680 ;
        RECT 1976.705 2810.495 1976.995 2810.540 ;
        RECT 2089.390 2810.480 2089.710 2810.540 ;
        RECT 1953.230 2805.240 1953.550 2805.300 ;
        RECT 1976.705 2805.240 1976.995 2805.285 ;
        RECT 1953.230 2805.100 1976.995 2805.240 ;
        RECT 1953.230 2805.040 1953.550 2805.100 ;
        RECT 1976.705 2805.055 1976.995 2805.100 ;
        RECT 19.390 2798.780 19.710 2798.840 ;
        RECT 1861.245 2798.780 1861.535 2798.825 ;
        RECT 19.390 2798.640 1861.535 2798.780 ;
        RECT 19.390 2798.580 19.710 2798.640 ;
        RECT 1861.245 2798.595 1861.535 2798.640 ;
        RECT 1862.165 2798.780 1862.455 2798.825 ;
        RECT 1952.770 2798.780 1953.090 2798.840 ;
        RECT 1862.165 2798.640 1953.090 2798.780 ;
        RECT 1862.165 2798.595 1862.455 2798.640 ;
        RECT 1952.770 2798.580 1953.090 2798.640 ;
      LAYER via ;
        RECT 2089.420 2810.480 2089.680 2810.740 ;
        RECT 1953.260 2805.040 1953.520 2805.300 ;
        RECT 19.420 2798.580 19.680 2798.840 ;
        RECT 1952.800 2798.580 1953.060 2798.840 ;
      LAYER met2 ;
        RECT 2089.420 2810.450 2089.680 2810.770 ;
        RECT 1953.260 2805.010 1953.520 2805.330 ;
        RECT 19.420 2798.550 19.680 2798.870 ;
        RECT 1952.800 2798.610 1953.060 2798.870 ;
        RECT 1953.320 2798.610 1953.460 2805.010 ;
        RECT 2089.480 2800.000 2089.620 2810.450 ;
        RECT 1952.800 2798.550 1953.460 2798.610 ;
        RECT 19.480 1113.005 19.620 2798.550 ;
        RECT 1952.860 2798.470 1953.460 2798.550 ;
        RECT 2089.345 2796.000 2089.625 2800.000 ;
        RECT 19.410 1112.635 19.690 1113.005 ;
      LAYER via2 ;
        RECT 19.410 1112.680 19.690 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 19.385 1112.970 19.715 1112.985 ;
        RECT -4.800 1112.670 19.715 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 19.385 1112.655 19.715 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 899.200 14.190 899.260 ;
        RECT 25.370 899.200 25.690 899.260 ;
        RECT 13.870 899.060 25.690 899.200 ;
        RECT 13.870 899.000 14.190 899.060 ;
        RECT 25.370 899.000 25.690 899.060 ;
      LAYER via ;
        RECT 13.900 899.000 14.160 899.260 ;
        RECT 25.400 899.000 25.660 899.260 ;
      LAYER met2 ;
        RECT 25.390 2810.595 25.670 2810.965 ;
        RECT 2118.390 2810.595 2118.670 2810.965 ;
        RECT 25.460 899.290 25.600 2810.595 ;
        RECT 2118.460 2800.000 2118.600 2810.595 ;
        RECT 2118.325 2796.000 2118.605 2800.000 ;
        RECT 13.900 898.970 14.160 899.290 ;
        RECT 25.400 898.970 25.660 899.290 ;
        RECT 13.960 897.445 14.100 898.970 ;
        RECT 13.890 897.075 14.170 897.445 ;
      LAYER via2 ;
        RECT 25.390 2810.640 25.670 2810.920 ;
        RECT 2118.390 2810.640 2118.670 2810.920 ;
        RECT 13.890 897.120 14.170 897.400 ;
      LAYER met3 ;
        RECT 25.365 2810.930 25.695 2810.945 ;
        RECT 2118.365 2810.930 2118.695 2810.945 ;
        RECT 25.365 2810.630 2118.695 2810.930 ;
        RECT 25.365 2810.615 25.695 2810.630 ;
        RECT 2118.365 2810.615 2118.695 2810.630 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 681.940 14.190 682.000 ;
        RECT 24.450 681.940 24.770 682.000 ;
        RECT 13.870 681.800 24.770 681.940 ;
        RECT 13.870 681.740 14.190 681.800 ;
        RECT 24.450 681.740 24.770 681.800 ;
      LAYER via ;
        RECT 13.900 681.740 14.160 682.000 ;
        RECT 24.480 681.740 24.740 682.000 ;
      LAYER met2 ;
        RECT 24.470 2809.235 24.750 2809.605 ;
        RECT 2147.370 2809.235 2147.650 2809.605 ;
        RECT 24.540 682.030 24.680 2809.235 ;
        RECT 2147.440 2800.000 2147.580 2809.235 ;
        RECT 2147.305 2796.000 2147.585 2800.000 ;
        RECT 13.900 681.885 14.160 682.030 ;
        RECT 13.890 681.515 14.170 681.885 ;
        RECT 24.480 681.710 24.740 682.030 ;
      LAYER via2 ;
        RECT 24.470 2809.280 24.750 2809.560 ;
        RECT 2147.370 2809.280 2147.650 2809.560 ;
        RECT 13.890 681.560 14.170 681.840 ;
      LAYER met3 ;
        RECT 24.445 2809.570 24.775 2809.585 ;
        RECT 2147.345 2809.570 2147.675 2809.585 ;
        RECT 24.445 2809.270 2147.675 2809.570 ;
        RECT 24.445 2809.255 24.775 2809.270 ;
        RECT 2147.345 2809.255 2147.675 2809.270 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 13.865 681.850 14.195 681.865 ;
        RECT -4.800 681.550 14.195 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 13.865 681.535 14.195 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1148.765 2796.245 1148.935 2797.435 ;
        RECT 1183.725 2796.585 1183.895 2797.435 ;
        RECT 1981.365 2796.925 1982.455 2797.095 ;
        RECT 2041.625 2796.925 2042.715 2797.095 ;
        RECT 1981.365 2796.585 1981.535 2796.925 ;
        RECT 48.445 2794.885 48.615 2795.735 ;
        RECT 96.285 2794.885 96.455 2796.075 ;
        RECT 102.265 2795.225 102.435 2796.075 ;
        RECT 207.605 2795.735 207.775 2796.075 ;
        RECT 145.045 2794.545 145.215 2795.395 ;
        RECT 192.885 2794.545 193.055 2795.735 ;
        RECT 206.685 2795.565 207.775 2795.735 ;
        RECT 241.645 2794.885 241.815 2796.075 ;
        RECT 304.205 2795.735 304.375 2796.075 ;
        RECT 289.485 2794.885 289.655 2795.735 ;
        RECT 303.285 2795.565 304.375 2795.735 ;
        RECT 338.245 2794.885 338.415 2796.075 ;
        RECT 400.805 2795.735 400.975 2796.075 ;
        RECT 386.085 2794.885 386.255 2795.735 ;
        RECT 399.885 2795.565 400.975 2795.735 ;
        RECT 434.845 2794.885 435.015 2796.075 ;
        RECT 497.405 2795.735 497.575 2796.075 ;
        RECT 482.685 2794.885 482.855 2795.735 ;
        RECT 496.485 2795.565 497.575 2795.735 ;
        RECT 531.445 2794.885 531.615 2796.075 ;
        RECT 594.005 2795.735 594.175 2796.075 ;
        RECT 579.285 2794.885 579.455 2795.735 ;
        RECT 593.085 2795.565 594.175 2795.735 ;
        RECT 628.045 2794.885 628.215 2796.075 ;
        RECT 690.605 2795.735 690.775 2796.075 ;
        RECT 675.885 2794.885 676.055 2795.735 ;
        RECT 689.685 2795.565 690.775 2795.735 ;
        RECT 724.645 2794.885 724.815 2796.075 ;
        RECT 787.205 2795.735 787.375 2796.075 ;
        RECT 772.485 2794.885 772.655 2795.735 ;
        RECT 786.285 2795.565 787.375 2795.735 ;
        RECT 821.245 2794.885 821.415 2796.075 ;
        RECT 883.805 2795.735 883.975 2796.075 ;
        RECT 869.085 2794.885 869.255 2795.735 ;
        RECT 882.885 2795.565 883.975 2795.735 ;
        RECT 917.845 2794.885 918.015 2796.075 ;
        RECT 980.405 2795.735 980.575 2796.075 ;
        RECT 965.685 2794.885 965.855 2795.735 ;
        RECT 979.485 2795.565 980.575 2795.735 ;
        RECT 1014.445 2794.885 1014.615 2796.075 ;
        RECT 1062.285 2794.885 1062.455 2795.735 ;
      LAYER mcon ;
        RECT 1148.765 2797.265 1148.935 2797.435 ;
        RECT 1183.725 2797.265 1183.895 2797.435 ;
        RECT 1982.285 2796.925 1982.455 2797.095 ;
        RECT 2042.545 2796.925 2042.715 2797.095 ;
        RECT 96.285 2795.905 96.455 2796.075 ;
        RECT 48.445 2795.565 48.615 2795.735 ;
        RECT 102.265 2795.905 102.435 2796.075 ;
        RECT 207.605 2795.905 207.775 2796.075 ;
        RECT 192.885 2795.565 193.055 2795.735 ;
        RECT 241.645 2795.905 241.815 2796.075 ;
        RECT 145.045 2795.225 145.215 2795.395 ;
        RECT 304.205 2795.905 304.375 2796.075 ;
        RECT 289.485 2795.565 289.655 2795.735 ;
        RECT 338.245 2795.905 338.415 2796.075 ;
        RECT 400.805 2795.905 400.975 2796.075 ;
        RECT 386.085 2795.565 386.255 2795.735 ;
        RECT 434.845 2795.905 435.015 2796.075 ;
        RECT 497.405 2795.905 497.575 2796.075 ;
        RECT 482.685 2795.565 482.855 2795.735 ;
        RECT 531.445 2795.905 531.615 2796.075 ;
        RECT 594.005 2795.905 594.175 2796.075 ;
        RECT 579.285 2795.565 579.455 2795.735 ;
        RECT 628.045 2795.905 628.215 2796.075 ;
        RECT 690.605 2795.905 690.775 2796.075 ;
        RECT 675.885 2795.565 676.055 2795.735 ;
        RECT 724.645 2795.905 724.815 2796.075 ;
        RECT 787.205 2795.905 787.375 2796.075 ;
        RECT 772.485 2795.565 772.655 2795.735 ;
        RECT 821.245 2795.905 821.415 2796.075 ;
        RECT 883.805 2795.905 883.975 2796.075 ;
        RECT 869.085 2795.565 869.255 2795.735 ;
        RECT 917.845 2795.905 918.015 2796.075 ;
        RECT 980.405 2795.905 980.575 2796.075 ;
        RECT 965.685 2795.565 965.855 2795.735 ;
        RECT 1014.445 2795.905 1014.615 2796.075 ;
        RECT 1062.285 2795.565 1062.455 2795.735 ;
      LAYER met1 ;
        RECT 1148.705 2797.420 1148.995 2797.465 ;
        RECT 1183.665 2797.420 1183.955 2797.465 ;
        RECT 1148.705 2797.280 1183.955 2797.420 ;
        RECT 1148.705 2797.235 1148.995 2797.280 ;
        RECT 1183.665 2797.235 1183.955 2797.280 ;
        RECT 1982.225 2797.080 1982.515 2797.125 ;
        RECT 2041.565 2797.080 2041.855 2797.125 ;
        RECT 1982.225 2796.940 2041.855 2797.080 ;
        RECT 1982.225 2796.895 1982.515 2796.940 ;
        RECT 2041.565 2796.895 2041.855 2796.940 ;
        RECT 2042.485 2796.895 2042.775 2797.125 ;
        RECT 2174.950 2797.080 2175.270 2797.140 ;
        RECT 2079.820 2796.940 2175.270 2797.080 ;
        RECT 1183.665 2796.555 1183.955 2796.785 ;
        RECT 1148.705 2796.400 1148.995 2796.445 ;
        RECT 1124.400 2796.260 1148.995 2796.400 ;
        RECT 1183.740 2796.400 1183.880 2796.555 ;
        RECT 1849.270 2796.540 1849.590 2796.800 ;
        RECT 1925.630 2796.540 1925.950 2796.800 ;
        RECT 1981.305 2796.555 1981.595 2796.785 ;
        RECT 1849.360 2796.400 1849.500 2796.540 ;
        RECT 1183.740 2796.260 1849.500 2796.400 ;
        RECT 1925.720 2796.400 1925.860 2796.540 ;
        RECT 1981.380 2796.400 1981.520 2796.555 ;
        RECT 1925.720 2796.260 1981.520 2796.400 ;
        RECT 2042.560 2796.400 2042.700 2796.895 ;
        RECT 2079.820 2796.400 2079.960 2796.940 ;
        RECT 2174.950 2796.880 2175.270 2796.940 ;
        RECT 2042.560 2796.260 2079.960 2796.400 ;
        RECT 96.225 2796.060 96.515 2796.105 ;
        RECT 102.205 2796.060 102.495 2796.105 ;
        RECT 96.225 2795.920 102.495 2796.060 ;
        RECT 96.225 2795.875 96.515 2795.920 ;
        RECT 102.205 2795.875 102.495 2795.920 ;
        RECT 207.545 2796.060 207.835 2796.105 ;
        RECT 241.585 2796.060 241.875 2796.105 ;
        RECT 207.545 2795.920 241.875 2796.060 ;
        RECT 207.545 2795.875 207.835 2795.920 ;
        RECT 241.585 2795.875 241.875 2795.920 ;
        RECT 304.145 2796.060 304.435 2796.105 ;
        RECT 338.185 2796.060 338.475 2796.105 ;
        RECT 304.145 2795.920 338.475 2796.060 ;
        RECT 304.145 2795.875 304.435 2795.920 ;
        RECT 338.185 2795.875 338.475 2795.920 ;
        RECT 400.745 2796.060 401.035 2796.105 ;
        RECT 434.785 2796.060 435.075 2796.105 ;
        RECT 400.745 2795.920 435.075 2796.060 ;
        RECT 400.745 2795.875 401.035 2795.920 ;
        RECT 434.785 2795.875 435.075 2795.920 ;
        RECT 497.345 2796.060 497.635 2796.105 ;
        RECT 531.385 2796.060 531.675 2796.105 ;
        RECT 497.345 2795.920 531.675 2796.060 ;
        RECT 497.345 2795.875 497.635 2795.920 ;
        RECT 531.385 2795.875 531.675 2795.920 ;
        RECT 593.945 2796.060 594.235 2796.105 ;
        RECT 627.985 2796.060 628.275 2796.105 ;
        RECT 593.945 2795.920 628.275 2796.060 ;
        RECT 593.945 2795.875 594.235 2795.920 ;
        RECT 627.985 2795.875 628.275 2795.920 ;
        RECT 690.545 2796.060 690.835 2796.105 ;
        RECT 724.585 2796.060 724.875 2796.105 ;
        RECT 690.545 2795.920 724.875 2796.060 ;
        RECT 690.545 2795.875 690.835 2795.920 ;
        RECT 724.585 2795.875 724.875 2795.920 ;
        RECT 787.145 2796.060 787.435 2796.105 ;
        RECT 821.185 2796.060 821.475 2796.105 ;
        RECT 787.145 2795.920 821.475 2796.060 ;
        RECT 787.145 2795.875 787.435 2795.920 ;
        RECT 821.185 2795.875 821.475 2795.920 ;
        RECT 883.745 2796.060 884.035 2796.105 ;
        RECT 917.785 2796.060 918.075 2796.105 ;
        RECT 883.745 2795.920 918.075 2796.060 ;
        RECT 883.745 2795.875 884.035 2795.920 ;
        RECT 917.785 2795.875 918.075 2795.920 ;
        RECT 980.345 2796.060 980.635 2796.105 ;
        RECT 1014.385 2796.060 1014.675 2796.105 ;
        RECT 1124.400 2796.060 1124.540 2796.260 ;
        RECT 1148.705 2796.215 1148.995 2796.260 ;
        RECT 980.345 2795.920 1014.675 2796.060 ;
        RECT 980.345 2795.875 980.635 2795.920 ;
        RECT 1014.385 2795.875 1014.675 2795.920 ;
        RECT 1076.560 2795.920 1124.540 2796.060 ;
        RECT 17.550 2795.720 17.870 2795.780 ;
        RECT 48.385 2795.720 48.675 2795.765 ;
        RECT 17.550 2795.580 48.675 2795.720 ;
        RECT 17.550 2795.520 17.870 2795.580 ;
        RECT 48.385 2795.535 48.675 2795.580 ;
        RECT 192.825 2795.720 193.115 2795.765 ;
        RECT 206.625 2795.720 206.915 2795.765 ;
        RECT 192.825 2795.580 206.915 2795.720 ;
        RECT 192.825 2795.535 193.115 2795.580 ;
        RECT 206.625 2795.535 206.915 2795.580 ;
        RECT 289.425 2795.720 289.715 2795.765 ;
        RECT 303.225 2795.720 303.515 2795.765 ;
        RECT 289.425 2795.580 303.515 2795.720 ;
        RECT 289.425 2795.535 289.715 2795.580 ;
        RECT 303.225 2795.535 303.515 2795.580 ;
        RECT 386.025 2795.720 386.315 2795.765 ;
        RECT 399.825 2795.720 400.115 2795.765 ;
        RECT 386.025 2795.580 400.115 2795.720 ;
        RECT 386.025 2795.535 386.315 2795.580 ;
        RECT 399.825 2795.535 400.115 2795.580 ;
        RECT 482.625 2795.720 482.915 2795.765 ;
        RECT 496.425 2795.720 496.715 2795.765 ;
        RECT 482.625 2795.580 496.715 2795.720 ;
        RECT 482.625 2795.535 482.915 2795.580 ;
        RECT 496.425 2795.535 496.715 2795.580 ;
        RECT 579.225 2795.720 579.515 2795.765 ;
        RECT 593.025 2795.720 593.315 2795.765 ;
        RECT 579.225 2795.580 593.315 2795.720 ;
        RECT 579.225 2795.535 579.515 2795.580 ;
        RECT 593.025 2795.535 593.315 2795.580 ;
        RECT 675.825 2795.720 676.115 2795.765 ;
        RECT 689.625 2795.720 689.915 2795.765 ;
        RECT 675.825 2795.580 689.915 2795.720 ;
        RECT 675.825 2795.535 676.115 2795.580 ;
        RECT 689.625 2795.535 689.915 2795.580 ;
        RECT 772.425 2795.720 772.715 2795.765 ;
        RECT 786.225 2795.720 786.515 2795.765 ;
        RECT 772.425 2795.580 786.515 2795.720 ;
        RECT 772.425 2795.535 772.715 2795.580 ;
        RECT 786.225 2795.535 786.515 2795.580 ;
        RECT 869.025 2795.720 869.315 2795.765 ;
        RECT 882.825 2795.720 883.115 2795.765 ;
        RECT 869.025 2795.580 883.115 2795.720 ;
        RECT 869.025 2795.535 869.315 2795.580 ;
        RECT 882.825 2795.535 883.115 2795.580 ;
        RECT 965.625 2795.720 965.915 2795.765 ;
        RECT 979.425 2795.720 979.715 2795.765 ;
        RECT 965.625 2795.580 979.715 2795.720 ;
        RECT 965.625 2795.535 965.915 2795.580 ;
        RECT 979.425 2795.535 979.715 2795.580 ;
        RECT 1062.225 2795.720 1062.515 2795.765 ;
        RECT 1076.560 2795.720 1076.700 2795.920 ;
        RECT 1062.225 2795.580 1076.700 2795.720 ;
        RECT 1062.225 2795.535 1062.515 2795.580 ;
        RECT 102.205 2795.380 102.495 2795.425 ;
        RECT 144.985 2795.380 145.275 2795.425 ;
        RECT 102.205 2795.240 145.275 2795.380 ;
        RECT 102.205 2795.195 102.495 2795.240 ;
        RECT 144.985 2795.195 145.275 2795.240 ;
        RECT 48.385 2795.040 48.675 2795.085 ;
        RECT 96.225 2795.040 96.515 2795.085 ;
        RECT 48.385 2794.900 96.515 2795.040 ;
        RECT 48.385 2794.855 48.675 2794.900 ;
        RECT 96.225 2794.855 96.515 2794.900 ;
        RECT 241.585 2795.040 241.875 2795.085 ;
        RECT 289.425 2795.040 289.715 2795.085 ;
        RECT 241.585 2794.900 289.715 2795.040 ;
        RECT 241.585 2794.855 241.875 2794.900 ;
        RECT 289.425 2794.855 289.715 2794.900 ;
        RECT 338.185 2795.040 338.475 2795.085 ;
        RECT 386.025 2795.040 386.315 2795.085 ;
        RECT 338.185 2794.900 386.315 2795.040 ;
        RECT 338.185 2794.855 338.475 2794.900 ;
        RECT 386.025 2794.855 386.315 2794.900 ;
        RECT 434.785 2795.040 435.075 2795.085 ;
        RECT 482.625 2795.040 482.915 2795.085 ;
        RECT 434.785 2794.900 482.915 2795.040 ;
        RECT 434.785 2794.855 435.075 2794.900 ;
        RECT 482.625 2794.855 482.915 2794.900 ;
        RECT 531.385 2795.040 531.675 2795.085 ;
        RECT 579.225 2795.040 579.515 2795.085 ;
        RECT 531.385 2794.900 579.515 2795.040 ;
        RECT 531.385 2794.855 531.675 2794.900 ;
        RECT 579.225 2794.855 579.515 2794.900 ;
        RECT 627.985 2795.040 628.275 2795.085 ;
        RECT 675.825 2795.040 676.115 2795.085 ;
        RECT 627.985 2794.900 676.115 2795.040 ;
        RECT 627.985 2794.855 628.275 2794.900 ;
        RECT 675.825 2794.855 676.115 2794.900 ;
        RECT 724.585 2795.040 724.875 2795.085 ;
        RECT 772.425 2795.040 772.715 2795.085 ;
        RECT 724.585 2794.900 772.715 2795.040 ;
        RECT 724.585 2794.855 724.875 2794.900 ;
        RECT 772.425 2794.855 772.715 2794.900 ;
        RECT 821.185 2795.040 821.475 2795.085 ;
        RECT 869.025 2795.040 869.315 2795.085 ;
        RECT 821.185 2794.900 869.315 2795.040 ;
        RECT 821.185 2794.855 821.475 2794.900 ;
        RECT 869.025 2794.855 869.315 2794.900 ;
        RECT 917.785 2795.040 918.075 2795.085 ;
        RECT 965.625 2795.040 965.915 2795.085 ;
        RECT 917.785 2794.900 965.915 2795.040 ;
        RECT 917.785 2794.855 918.075 2794.900 ;
        RECT 965.625 2794.855 965.915 2794.900 ;
        RECT 1014.385 2795.040 1014.675 2795.085 ;
        RECT 1062.225 2795.040 1062.515 2795.085 ;
        RECT 1014.385 2794.900 1062.515 2795.040 ;
        RECT 1014.385 2794.855 1014.675 2794.900 ;
        RECT 1062.225 2794.855 1062.515 2794.900 ;
        RECT 144.985 2794.700 145.275 2794.745 ;
        RECT 192.825 2794.700 193.115 2794.745 ;
        RECT 144.985 2794.560 193.115 2794.700 ;
        RECT 144.985 2794.515 145.275 2794.560 ;
        RECT 192.825 2794.515 193.115 2794.560 ;
      LAYER via ;
        RECT 1849.300 2796.540 1849.560 2796.800 ;
        RECT 1925.660 2796.540 1925.920 2796.800 ;
        RECT 2174.980 2796.880 2175.240 2797.140 ;
        RECT 17.580 2795.520 17.840 2795.780 ;
      LAYER met2 ;
        RECT 1925.650 2799.715 1925.930 2800.085 ;
        RECT 1849.290 2797.675 1849.570 2798.045 ;
        RECT 1849.360 2796.830 1849.500 2797.675 ;
        RECT 1925.720 2796.830 1925.860 2799.715 ;
        RECT 2176.285 2797.250 2176.565 2800.000 ;
        RECT 2175.040 2797.170 2176.565 2797.250 ;
        RECT 2174.980 2797.110 2176.565 2797.170 ;
        RECT 2174.980 2796.850 2175.240 2797.110 ;
        RECT 1849.300 2796.510 1849.560 2796.830 ;
        RECT 1925.660 2796.510 1925.920 2796.830 ;
        RECT 2176.285 2796.000 2176.565 2797.110 ;
        RECT 17.580 2795.490 17.840 2795.810 ;
        RECT 17.640 466.325 17.780 2795.490 ;
        RECT 17.570 465.955 17.850 466.325 ;
      LAYER via2 ;
        RECT 1925.650 2799.760 1925.930 2800.040 ;
        RECT 1849.290 2797.720 1849.570 2798.000 ;
        RECT 17.570 466.000 17.850 466.280 ;
      LAYER met3 ;
        RECT 1925.625 2800.050 1925.955 2800.065 ;
        RECT 1893.670 2799.750 1925.955 2800.050 ;
        RECT 1849.265 2798.010 1849.595 2798.025 ;
        RECT 1893.670 2798.010 1893.970 2799.750 ;
        RECT 1925.625 2799.735 1925.955 2799.750 ;
        RECT 1849.265 2797.710 1893.970 2798.010 ;
        RECT 1849.265 2797.695 1849.595 2797.710 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.545 466.290 17.875 466.305 ;
        RECT -4.800 465.990 17.875 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.545 465.975 17.875 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.790 2813.315 21.070 2813.685 ;
        RECT 2205.330 2813.315 2205.610 2813.685 ;
        RECT 20.330 250.650 20.610 250.765 ;
        RECT 20.860 250.650 21.000 2813.315 ;
        RECT 2205.400 2800.000 2205.540 2813.315 ;
        RECT 2205.265 2796.000 2205.545 2800.000 ;
        RECT 20.330 250.510 21.000 250.650 ;
        RECT 20.330 250.395 20.610 250.510 ;
      LAYER via2 ;
        RECT 20.790 2813.360 21.070 2813.640 ;
        RECT 2205.330 2813.360 2205.610 2813.640 ;
        RECT 20.330 250.440 20.610 250.720 ;
      LAYER met3 ;
        RECT 1786.910 2815.690 1787.290 2815.700 ;
        RECT 1834.750 2815.690 1835.130 2815.700 ;
        RECT 1786.910 2815.390 1835.130 2815.690 ;
        RECT 1786.910 2815.380 1787.290 2815.390 ;
        RECT 1834.750 2815.380 1835.130 2815.390 ;
        RECT 1262.510 2815.010 1262.890 2815.020 ;
        RECT 1268.030 2815.010 1268.410 2815.020 ;
        RECT 1262.510 2814.710 1268.410 2815.010 ;
        RECT 1262.510 2814.700 1262.890 2814.710 ;
        RECT 1268.030 2814.700 1268.410 2814.710 ;
        RECT 1331.510 2815.010 1331.890 2815.020 ;
        RECT 1379.350 2815.010 1379.730 2815.020 ;
        RECT 1331.510 2814.710 1379.730 2815.010 ;
        RECT 1331.510 2814.700 1331.890 2814.710 ;
        RECT 1379.350 2814.700 1379.730 2814.710 ;
        RECT 20.765 2813.650 21.095 2813.665 ;
        RECT 26.030 2813.650 26.410 2813.660 ;
        RECT 20.765 2813.350 26.410 2813.650 ;
        RECT 20.765 2813.335 21.095 2813.350 ;
        RECT 26.030 2813.340 26.410 2813.350 ;
        RECT 627.710 2813.650 628.090 2813.660 ;
        RECT 675.550 2813.650 675.930 2813.660 ;
        RECT 627.710 2813.350 675.930 2813.650 ;
        RECT 627.710 2813.340 628.090 2813.350 ;
        RECT 675.550 2813.340 675.930 2813.350 ;
        RECT 820.910 2813.650 821.290 2813.660 ;
        RECT 836.550 2813.650 836.930 2813.660 ;
        RECT 820.910 2813.350 836.930 2813.650 ;
        RECT 820.910 2813.340 821.290 2813.350 ;
        RECT 836.550 2813.340 836.930 2813.350 ;
        RECT 917.510 2813.650 917.890 2813.660 ;
        RECT 965.350 2813.650 965.730 2813.660 ;
        RECT 917.510 2813.350 965.730 2813.650 ;
        RECT 917.510 2813.340 917.890 2813.350 ;
        RECT 965.350 2813.340 965.730 2813.350 ;
        RECT 1025.150 2813.650 1025.530 2813.660 ;
        RECT 1038.030 2813.650 1038.410 2813.660 ;
        RECT 1025.150 2813.350 1038.410 2813.650 ;
        RECT 1025.150 2813.340 1025.530 2813.350 ;
        RECT 1038.030 2813.340 1038.410 2813.350 ;
        RECT 2121.790 2813.650 2122.170 2813.660 ;
        RECT 2142.030 2813.650 2142.410 2813.660 ;
        RECT 2121.790 2813.350 2142.410 2813.650 ;
        RECT 2121.790 2813.340 2122.170 2813.350 ;
        RECT 2142.030 2813.340 2142.410 2813.350 ;
        RECT 2180.670 2813.650 2181.050 2813.660 ;
        RECT 2205.305 2813.650 2205.635 2813.665 ;
        RECT 2180.670 2813.350 2205.635 2813.650 ;
        RECT 2180.670 2813.340 2181.050 2813.350 ;
        RECT 2205.305 2813.335 2205.635 2813.350 ;
        RECT 1441.910 2808.210 1442.290 2808.220 ;
        RECT 1465.830 2808.210 1466.210 2808.220 ;
        RECT 1441.910 2807.910 1466.210 2808.210 ;
        RECT 1441.910 2807.900 1442.290 2807.910 ;
        RECT 1465.830 2807.900 1466.210 2807.910 ;
        RECT 252.350 2806.850 252.730 2806.860 ;
        RECT 257.870 2806.850 258.250 2806.860 ;
        RECT 252.350 2806.550 258.250 2806.850 ;
        RECT 252.350 2806.540 252.730 2806.550 ;
        RECT 257.870 2806.540 258.250 2806.550 ;
        RECT 428.070 2806.850 428.450 2806.860 ;
        RECT 451.070 2806.850 451.450 2806.860 ;
        RECT 428.070 2806.550 451.450 2806.850 ;
        RECT 428.070 2806.540 428.450 2806.550 ;
        RECT 451.070 2806.540 451.450 2806.550 ;
        RECT 542.150 2806.850 542.530 2806.860 ;
        RECT 548.590 2806.850 548.970 2806.860 ;
        RECT 542.150 2806.550 548.970 2806.850 ;
        RECT 542.150 2806.540 542.530 2806.550 ;
        RECT 548.590 2806.540 548.970 2806.550 ;
        RECT 588.150 2806.850 588.530 2806.860 ;
        RECT 603.790 2806.850 604.170 2806.860 ;
        RECT 588.150 2806.550 604.170 2806.850 ;
        RECT 588.150 2806.540 588.530 2806.550 ;
        RECT 603.790 2806.540 604.170 2806.550 ;
        RECT 678.310 2806.850 678.690 2806.860 ;
        RECT 700.390 2806.850 700.770 2806.860 ;
        RECT 678.310 2806.550 700.770 2806.850 ;
        RECT 678.310 2806.540 678.690 2806.550 ;
        RECT 700.390 2806.540 700.770 2806.550 ;
        RECT 737.190 2806.850 737.570 2806.860 ;
        RECT 772.150 2806.850 772.530 2806.860 ;
        RECT 737.190 2806.550 772.530 2806.850 ;
        RECT 737.190 2806.540 737.570 2806.550 ;
        RECT 772.150 2806.540 772.530 2806.550 ;
        RECT 774.910 2806.850 775.290 2806.860 ;
        RECT 796.990 2806.850 797.370 2806.860 ;
        RECT 774.910 2806.550 797.370 2806.850 ;
        RECT 774.910 2806.540 775.290 2806.550 ;
        RECT 796.990 2806.540 797.370 2806.550 ;
        RECT 880.710 2806.850 881.090 2806.860 ;
        RECT 893.590 2806.850 893.970 2806.860 ;
        RECT 880.710 2806.550 893.970 2806.850 ;
        RECT 880.710 2806.540 881.090 2806.550 ;
        RECT 893.590 2806.540 893.970 2806.550 ;
        RECT 968.110 2806.850 968.490 2806.860 ;
        RECT 983.750 2806.850 984.130 2806.860 ;
        RECT 968.110 2806.550 984.130 2806.850 ;
        RECT 968.110 2806.540 968.490 2806.550 ;
        RECT 983.750 2806.540 984.130 2806.550 ;
        RECT 1118.070 2806.850 1118.450 2806.860 ;
        RECT 1127.270 2806.850 1127.650 2806.860 ;
        RECT 1118.070 2806.550 1127.650 2806.850 ;
        RECT 1118.070 2806.540 1118.450 2806.550 ;
        RECT 1127.270 2806.540 1127.650 2806.550 ;
        RECT 1628.670 2806.850 1629.050 2806.860 ;
        RECT 1675.590 2806.850 1675.970 2806.860 ;
        RECT 1628.670 2806.550 1675.970 2806.850 ;
        RECT 1628.670 2806.540 1629.050 2806.550 ;
        RECT 1675.590 2806.540 1675.970 2806.550 ;
        RECT 1966.310 2806.850 1966.690 2806.860 ;
        RECT 2031.630 2806.850 2032.010 2806.860 ;
        RECT 1966.310 2806.550 2032.010 2806.850 ;
        RECT 1966.310 2806.540 1966.690 2806.550 ;
        RECT 2031.630 2806.540 2032.010 2806.550 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 20.305 250.730 20.635 250.745 ;
        RECT -4.800 250.430 20.635 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 20.305 250.415 20.635 250.430 ;
      LAYER via3 ;
        RECT 1786.940 2815.380 1787.260 2815.700 ;
        RECT 1834.780 2815.380 1835.100 2815.700 ;
        RECT 1262.540 2814.700 1262.860 2815.020 ;
        RECT 1268.060 2814.700 1268.380 2815.020 ;
        RECT 1331.540 2814.700 1331.860 2815.020 ;
        RECT 1379.380 2814.700 1379.700 2815.020 ;
        RECT 26.060 2813.340 26.380 2813.660 ;
        RECT 627.740 2813.340 628.060 2813.660 ;
        RECT 675.580 2813.340 675.900 2813.660 ;
        RECT 820.940 2813.340 821.260 2813.660 ;
        RECT 836.580 2813.340 836.900 2813.660 ;
        RECT 917.540 2813.340 917.860 2813.660 ;
        RECT 965.380 2813.340 965.700 2813.660 ;
        RECT 1025.180 2813.340 1025.500 2813.660 ;
        RECT 1038.060 2813.340 1038.380 2813.660 ;
        RECT 2121.820 2813.340 2122.140 2813.660 ;
        RECT 2142.060 2813.340 2142.380 2813.660 ;
        RECT 2180.700 2813.340 2181.020 2813.660 ;
        RECT 1441.940 2807.900 1442.260 2808.220 ;
        RECT 1465.860 2807.900 1466.180 2808.220 ;
        RECT 252.380 2806.540 252.700 2806.860 ;
        RECT 257.900 2806.540 258.220 2806.860 ;
        RECT 428.100 2806.540 428.420 2806.860 ;
        RECT 451.100 2806.540 451.420 2806.860 ;
        RECT 542.180 2806.540 542.500 2806.860 ;
        RECT 548.620 2806.540 548.940 2806.860 ;
        RECT 588.180 2806.540 588.500 2806.860 ;
        RECT 603.820 2806.540 604.140 2806.860 ;
        RECT 678.340 2806.540 678.660 2806.860 ;
        RECT 700.420 2806.540 700.740 2806.860 ;
        RECT 737.220 2806.540 737.540 2806.860 ;
        RECT 772.180 2806.540 772.500 2806.860 ;
        RECT 774.940 2806.540 775.260 2806.860 ;
        RECT 797.020 2806.540 797.340 2806.860 ;
        RECT 880.740 2806.540 881.060 2806.860 ;
        RECT 893.620 2806.540 893.940 2806.860 ;
        RECT 968.140 2806.540 968.460 2806.860 ;
        RECT 983.780 2806.540 984.100 2806.860 ;
        RECT 1118.100 2806.540 1118.420 2806.860 ;
        RECT 1127.300 2806.540 1127.620 2806.860 ;
        RECT 1628.700 2806.540 1629.020 2806.860 ;
        RECT 1675.620 2806.540 1675.940 2806.860 ;
        RECT 1966.340 2806.540 1966.660 2806.860 ;
        RECT 2031.660 2806.540 2031.980 2806.860 ;
      LAYER met4 ;
        RECT 1786.935 2815.375 1787.265 2815.705 ;
        RECT 1834.775 2815.375 1835.105 2815.705 ;
        RECT 1262.535 2814.695 1262.865 2815.025 ;
        RECT 1268.055 2814.695 1268.385 2815.025 ;
        RECT 1331.535 2814.695 1331.865 2815.025 ;
        RECT 1379.375 2814.695 1379.705 2815.025 ;
        RECT 25.630 2812.910 26.810 2814.090 ;
        RECT 603.390 2812.910 604.570 2814.090 ;
        RECT 627.310 2812.910 628.490 2814.090 ;
        RECT 675.575 2813.335 675.905 2813.665 ;
        RECT 251.950 2806.110 253.130 2807.290 ;
        RECT 257.470 2806.110 258.650 2807.290 ;
        RECT 427.670 2806.110 428.850 2807.290 ;
        RECT 450.670 2806.110 451.850 2807.290 ;
        RECT 541.750 2806.110 542.930 2807.290 ;
        RECT 548.190 2806.110 549.370 2807.290 ;
        RECT 587.750 2806.110 588.930 2807.290 ;
        RECT 603.830 2806.865 604.130 2812.910 ;
        RECT 675.590 2807.290 675.890 2813.335 ;
        RECT 699.990 2812.910 701.170 2814.090 ;
        RECT 796.590 2812.910 797.770 2814.090 ;
        RECT 820.510 2812.910 821.690 2814.090 ;
        RECT 836.150 2812.910 837.330 2814.090 ;
        RECT 893.190 2812.910 894.370 2814.090 ;
        RECT 917.110 2812.910 918.290 2814.090 ;
        RECT 965.375 2813.335 965.705 2813.665 ;
        RECT 603.815 2806.535 604.145 2806.865 ;
        RECT 675.150 2806.110 676.330 2807.290 ;
        RECT 677.910 2806.110 679.090 2807.290 ;
        RECT 700.430 2806.865 700.730 2812.910 ;
        RECT 700.415 2806.535 700.745 2806.865 ;
        RECT 736.790 2806.110 737.970 2807.290 ;
        RECT 771.750 2806.110 772.930 2807.290 ;
        RECT 774.510 2806.110 775.690 2807.290 ;
        RECT 797.030 2806.865 797.330 2812.910 ;
        RECT 797.015 2806.535 797.345 2806.865 ;
        RECT 880.310 2806.110 881.490 2807.290 ;
        RECT 893.630 2806.865 893.930 2812.910 ;
        RECT 965.390 2807.290 965.690 2813.335 ;
        RECT 983.350 2812.910 984.530 2814.090 ;
        RECT 1024.750 2812.910 1025.930 2814.090 ;
        RECT 1038.055 2813.335 1038.385 2813.665 ;
        RECT 893.615 2806.535 893.945 2806.865 ;
        RECT 964.950 2806.110 966.130 2807.290 ;
        RECT 967.710 2806.110 968.890 2807.290 ;
        RECT 983.790 2806.865 984.090 2812.910 ;
        RECT 1038.070 2807.290 1038.370 2813.335 ;
        RECT 1262.550 2810.690 1262.850 2814.695 ;
        RECT 1268.070 2814.090 1268.370 2814.695 ;
        RECT 1267.630 2812.910 1268.810 2814.090 ;
        RECT 1331.550 2810.690 1331.850 2814.695 ;
        RECT 1379.390 2814.090 1379.690 2814.695 ;
        RECT 1786.950 2814.090 1787.250 2815.375 ;
        RECT 1378.950 2812.910 1380.130 2814.090 ;
        RECT 1465.430 2812.910 1466.610 2814.090 ;
        RECT 1675.190 2812.910 1676.370 2814.090 ;
        RECT 1683.470 2813.650 1684.650 2814.090 ;
        RECT 1683.470 2813.350 1686.970 2813.650 ;
        RECT 1683.470 2812.910 1684.650 2813.350 ;
        RECT 1126.870 2809.510 1128.050 2810.690 ;
        RECT 1262.110 2809.510 1263.290 2810.690 ;
        RECT 1331.110 2809.510 1332.290 2810.690 ;
        RECT 1441.510 2809.510 1442.690 2810.690 ;
        RECT 983.775 2806.535 984.105 2806.865 ;
        RECT 1037.630 2806.110 1038.810 2807.290 ;
        RECT 1117.670 2806.110 1118.850 2807.290 ;
        RECT 1127.310 2806.865 1127.610 2809.510 ;
        RECT 1441.950 2808.225 1442.250 2809.510 ;
        RECT 1465.870 2808.225 1466.170 2812.910 ;
        RECT 1441.935 2807.895 1442.265 2808.225 ;
        RECT 1465.855 2807.895 1466.185 2808.225 ;
        RECT 1127.295 2806.535 1127.625 2806.865 ;
        RECT 1592.390 2806.850 1593.570 2807.290 ;
        RECT 1596.070 2806.850 1597.250 2807.290 ;
        RECT 1592.390 2806.550 1597.250 2806.850 ;
        RECT 1592.390 2806.110 1593.570 2806.550 ;
        RECT 1596.070 2806.110 1597.250 2806.550 ;
        RECT 1628.270 2806.110 1629.450 2807.290 ;
        RECT 1675.630 2806.865 1675.930 2812.910 ;
        RECT 1686.670 2810.690 1686.970 2813.350 ;
        RECT 1786.510 2812.910 1787.690 2814.090 ;
        RECT 1834.790 2810.690 1835.090 2815.375 ;
        RECT 1851.830 2813.650 1853.010 2814.090 ;
        RECT 1846.750 2813.350 1853.010 2813.650 ;
        RECT 1846.750 2810.690 1847.050 2813.350 ;
        RECT 1851.830 2812.910 1853.010 2813.350 ;
        RECT 1965.910 2812.910 1967.090 2814.090 ;
        RECT 2121.390 2812.910 2122.570 2814.090 ;
        RECT 2141.630 2812.910 2142.810 2814.090 ;
        RECT 2180.270 2812.910 2181.450 2814.090 ;
        RECT 1686.230 2809.510 1687.410 2810.690 ;
        RECT 1834.350 2809.510 1835.530 2810.690 ;
        RECT 1846.310 2809.510 1847.490 2810.690 ;
        RECT 1966.350 2806.865 1966.650 2812.910 ;
        RECT 2031.230 2809.510 2032.410 2810.690 ;
        RECT 2031.670 2806.865 2031.970 2809.510 ;
        RECT 1675.615 2806.535 1675.945 2806.865 ;
        RECT 1966.335 2806.535 1966.665 2806.865 ;
        RECT 2031.655 2806.535 2031.985 2806.865 ;
      LAYER met5 ;
        RECT 1168.980 2814.300 1177.020 2814.980 ;
        RECT 25.420 2812.700 90.500 2814.300 ;
        RECT 88.900 2807.500 90.500 2812.700 ;
        RECT 155.140 2812.700 186.180 2814.300 ;
        RECT 155.140 2807.500 156.740 2812.700 ;
        RECT 88.900 2805.900 156.740 2807.500 ;
        RECT 184.580 2807.500 186.180 2812.700 ;
        RECT 377.780 2810.900 380.300 2814.300 ;
        RECT 603.180 2812.700 628.700 2814.300 ;
        RECT 699.780 2812.700 725.300 2814.300 ;
        RECT 796.380 2812.700 821.900 2814.300 ;
        RECT 835.940 2812.700 869.740 2814.300 ;
        RECT 892.980 2812.700 918.500 2814.300 ;
        RECT 983.140 2812.700 1026.140 2814.300 ;
        RECT 1054.900 2812.700 1104.340 2814.300 ;
        RECT 330.860 2809.300 380.300 2810.900 ;
        RECT 330.860 2807.500 332.460 2809.300 ;
        RECT 184.580 2805.900 253.340 2807.500 ;
        RECT 257.260 2805.900 332.460 2807.500 ;
        RECT 378.700 2807.500 380.300 2809.300 ;
        RECT 723.700 2807.500 725.300 2812.700 ;
        RECT 868.140 2807.500 869.740 2812.700 ;
        RECT 1054.900 2807.500 1056.500 2812.700 ;
        RECT 378.700 2805.900 429.060 2807.500 ;
        RECT 450.460 2805.900 543.140 2807.500 ;
        RECT 547.980 2805.900 589.140 2807.500 ;
        RECT 674.940 2805.900 679.300 2807.500 ;
        RECT 723.700 2805.900 738.180 2807.500 ;
        RECT 771.540 2805.900 775.900 2807.500 ;
        RECT 868.140 2805.900 881.700 2807.500 ;
        RECT 964.740 2805.900 969.100 2807.500 ;
        RECT 1037.420 2805.900 1056.500 2807.500 ;
        RECT 1102.740 2807.500 1104.340 2812.700 ;
        RECT 1168.980 2813.380 1222.100 2814.300 ;
        RECT 1168.980 2810.900 1170.580 2813.380 ;
        RECT 1175.420 2812.700 1222.100 2813.380 ;
        RECT 1267.420 2812.700 1319.620 2814.300 ;
        RECT 1378.740 2812.700 1425.420 2814.300 ;
        RECT 1465.220 2812.700 1499.020 2814.300 ;
        RECT 1126.660 2809.300 1170.580 2810.900 ;
        RECT 1220.500 2810.900 1222.100 2812.700 ;
        RECT 1318.020 2810.900 1319.620 2812.700 ;
        RECT 1423.820 2810.900 1425.420 2812.700 ;
        RECT 1220.500 2809.300 1263.500 2810.900 ;
        RECT 1318.020 2809.300 1332.500 2810.900 ;
        RECT 1423.820 2809.300 1442.900 2810.900 ;
        RECT 1497.420 2807.500 1499.020 2812.700 ;
        RECT 1585.740 2810.900 1588.260 2814.300 ;
        RECT 1674.980 2812.700 1684.860 2814.300 ;
        RECT 1747.660 2812.700 1787.900 2814.300 ;
        RECT 1851.620 2812.700 1884.500 2814.300 ;
        RECT 1747.660 2810.900 1749.260 2812.700 ;
        RECT 1882.900 2810.900 1884.500 2812.700 ;
        RECT 1896.700 2812.700 1932.340 2814.300 ;
        RECT 1896.700 2810.900 1898.300 2812.700 ;
        RECT 1537.900 2809.300 1588.260 2810.900 ;
        RECT 1686.020 2809.300 1749.260 2810.900 ;
        RECT 1834.140 2809.300 1847.700 2810.900 ;
        RECT 1882.900 2809.300 1898.300 2810.900 ;
        RECT 1537.900 2807.500 1539.500 2809.300 ;
        RECT 1102.740 2805.900 1119.060 2807.500 ;
        RECT 1497.420 2805.900 1539.500 2807.500 ;
        RECT 1586.660 2807.500 1588.260 2809.300 ;
        RECT 1930.740 2807.500 1932.340 2812.700 ;
        RECT 1941.780 2812.700 1967.300 2814.300 ;
        RECT 2055.860 2812.700 2122.780 2814.300 ;
        RECT 2141.420 2812.700 2181.660 2814.300 ;
        RECT 1941.780 2807.500 1943.380 2812.700 ;
        RECT 2055.860 2810.900 2057.460 2812.700 ;
        RECT 2031.020 2809.300 2057.460 2810.900 ;
        RECT 1586.660 2805.900 1593.780 2807.500 ;
        RECT 1595.860 2805.900 1629.660 2807.500 ;
        RECT 1930.740 2805.900 1943.380 2807.500 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2232.930 2796.570 2233.210 2796.685 ;
        RECT 2234.245 2796.570 2234.525 2800.000 ;
        RECT 2232.930 2796.430 2234.525 2796.570 ;
        RECT 2232.930 2796.315 2233.210 2796.430 ;
        RECT 2234.245 2796.000 2234.525 2796.430 ;
        RECT 20.330 40.955 20.610 41.325 ;
        RECT 20.400 35.885 20.540 40.955 ;
        RECT 20.330 35.515 20.610 35.885 ;
      LAYER via2 ;
        RECT 2232.930 2796.360 2233.210 2796.640 ;
        RECT 20.330 41.000 20.610 41.280 ;
        RECT 20.330 35.560 20.610 35.840 ;
      LAYER met3 ;
        RECT 2228.510 2796.650 2228.890 2796.660 ;
        RECT 2232.905 2796.650 2233.235 2796.665 ;
        RECT 2228.510 2796.350 2233.235 2796.650 ;
        RECT 2228.510 2796.340 2228.890 2796.350 ;
        RECT 2232.905 2796.335 2233.235 2796.350 ;
        RECT 20.305 41.290 20.635 41.305 ;
        RECT 2228.510 41.290 2228.890 41.300 ;
        RECT 20.305 40.990 2228.890 41.290 ;
        RECT 20.305 40.975 20.635 40.990 ;
        RECT 2228.510 40.980 2228.890 40.990 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 20.305 35.850 20.635 35.865 ;
        RECT -4.800 35.550 20.635 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 20.305 35.535 20.635 35.550 ;
      LAYER via3 ;
        RECT 2228.540 2796.340 2228.860 2796.660 ;
        RECT 2228.540 40.980 2228.860 41.300 ;
      LAYER met4 ;
        RECT 2228.535 2796.335 2228.865 2796.665 ;
        RECT 2228.550 41.305 2228.850 2796.335 ;
        RECT 2228.535 40.975 2228.865 41.305 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1545.210 905.320 1545.530 905.380 ;
        RECT 1560.390 905.320 1560.710 905.380 ;
        RECT 1545.210 905.180 1560.710 905.320 ;
        RECT 1545.210 905.120 1545.530 905.180 ;
        RECT 1560.390 905.120 1560.710 905.180 ;
        RECT 1992.330 904.980 1992.650 905.040 ;
        RECT 1995.090 904.980 1995.410 905.040 ;
        RECT 1992.330 904.840 1995.410 904.980 ;
        RECT 1992.330 904.780 1992.650 904.840 ;
        RECT 1995.090 904.780 1995.410 904.840 ;
        RECT 2089.390 904.980 2089.710 905.040 ;
        RECT 2091.690 904.980 2092.010 905.040 ;
        RECT 2089.390 904.840 2092.010 904.980 ;
        RECT 2089.390 904.780 2089.710 904.840 ;
        RECT 2091.690 904.780 2092.010 904.840 ;
        RECT 2272.010 904.640 2272.330 904.700 ;
        RECT 2291.790 904.640 2292.110 904.700 ;
        RECT 2272.010 904.500 2292.110 904.640 ;
        RECT 2272.010 904.440 2272.330 904.500 ;
        RECT 2291.790 904.440 2292.110 904.500 ;
        RECT 1352.470 904.300 1352.790 904.360 ;
        RECT 1376.850 904.300 1377.170 904.360 ;
        RECT 1352.470 904.160 1377.170 904.300 ;
        RECT 1352.470 904.100 1352.790 904.160 ;
        RECT 1376.850 904.100 1377.170 904.160 ;
      LAYER via ;
        RECT 1545.240 905.120 1545.500 905.380 ;
        RECT 1560.420 905.120 1560.680 905.380 ;
        RECT 1992.360 904.780 1992.620 905.040 ;
        RECT 1995.120 904.780 1995.380 905.040 ;
        RECT 2089.420 904.780 2089.680 905.040 ;
        RECT 2091.720 904.780 2091.980 905.040 ;
        RECT 2272.040 904.440 2272.300 904.700 ;
        RECT 2291.820 904.440 2292.080 904.700 ;
        RECT 1352.500 904.100 1352.760 904.360 ;
        RECT 1376.880 904.100 1377.140 904.360 ;
      LAYER met2 ;
        RECT 1249.910 2814.675 1250.190 2815.045 ;
        RECT 1249.980 2800.000 1250.120 2814.675 ;
        RECT 1249.845 2796.000 1250.125 2800.000 ;
        RECT 1810.650 907.275 1810.930 907.645 ;
        RECT 1634.930 906.595 1635.210 906.965 ;
        RECT 1635.000 905.605 1635.140 906.595 ;
        RECT 1376.870 905.235 1377.150 905.605 ;
        RECT 1545.230 905.235 1545.510 905.605 ;
        RECT 1560.410 905.235 1560.690 905.605 ;
        RECT 1634.930 905.235 1635.210 905.605 ;
        RECT 1376.940 904.390 1377.080 905.235 ;
        RECT 1545.240 905.090 1545.500 905.235 ;
        RECT 1560.420 905.090 1560.680 905.235 ;
        RECT 1352.500 904.245 1352.760 904.390 ;
        RECT 1352.490 903.875 1352.770 904.245 ;
        RECT 1376.880 904.070 1377.140 904.390 ;
        RECT 1810.720 904.245 1810.860 907.275 ;
        RECT 1992.360 904.925 1992.620 905.070 ;
        RECT 1995.120 904.925 1995.380 905.070 ;
        RECT 2089.420 904.925 2089.680 905.070 ;
        RECT 2091.720 904.925 2091.980 905.070 ;
        RECT 1992.350 904.555 1992.630 904.925 ;
        RECT 1995.110 904.555 1995.390 904.925 ;
        RECT 2089.410 904.555 2089.690 904.925 ;
        RECT 2091.710 904.555 2091.990 904.925 ;
        RECT 2272.030 904.555 2272.310 904.925 ;
        RECT 2291.810 904.555 2292.090 904.925 ;
        RECT 2272.040 904.410 2272.300 904.555 ;
        RECT 2291.820 904.410 2292.080 904.555 ;
        RECT 1810.650 903.875 1810.930 904.245 ;
      LAYER via2 ;
        RECT 1249.910 2814.720 1250.190 2815.000 ;
        RECT 1810.650 907.320 1810.930 907.600 ;
        RECT 1634.930 906.640 1635.210 906.920 ;
        RECT 1376.870 905.280 1377.150 905.560 ;
        RECT 1545.230 905.280 1545.510 905.560 ;
        RECT 1560.410 905.280 1560.690 905.560 ;
        RECT 1634.930 905.280 1635.210 905.560 ;
        RECT 1352.490 903.920 1352.770 904.200 ;
        RECT 1992.350 904.600 1992.630 904.880 ;
        RECT 1995.110 904.600 1995.390 904.880 ;
        RECT 2089.410 904.600 2089.690 904.880 ;
        RECT 2091.710 904.600 2091.990 904.880 ;
        RECT 2272.030 904.600 2272.310 904.880 ;
        RECT 2291.810 904.600 2292.090 904.880 ;
        RECT 1810.650 903.920 1810.930 904.200 ;
      LAYER met3 ;
        RECT 1188.910 2815.010 1189.290 2815.020 ;
        RECT 1249.885 2815.010 1250.215 2815.025 ;
        RECT 1188.910 2814.710 1250.215 2815.010 ;
        RECT 1188.910 2814.700 1189.290 2814.710 ;
        RECT 1249.885 2814.695 1250.215 2814.710 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2916.710 909.350 2924.800 909.650 ;
        RECT 1786.910 907.610 1787.290 907.620 ;
        RECT 1810.625 907.610 1810.955 907.625 ;
        RECT 1786.910 907.310 1810.955 907.610 ;
        RECT 1786.910 907.300 1787.290 907.310 ;
        RECT 1810.625 907.295 1810.955 907.310 ;
        RECT 1634.905 906.930 1635.235 906.945 ;
        RECT 1587.310 906.630 1635.235 906.930 ;
        RECT 1496.190 906.250 1496.570 906.260 ;
        RECT 1462.190 905.950 1496.570 906.250 ;
        RECT 1188.910 905.570 1189.290 905.580 ;
        RECT 1207.310 905.570 1207.690 905.580 ;
        RECT 1376.845 905.570 1377.175 905.585 ;
        RECT 1188.910 905.270 1207.690 905.570 ;
        RECT 1188.910 905.260 1189.290 905.270 ;
        RECT 1207.310 905.260 1207.690 905.270 ;
        RECT 1272.670 905.270 1304.250 905.570 ;
        RECT 1207.310 904.210 1207.690 904.220 ;
        RECT 1272.670 904.210 1272.970 905.270 ;
        RECT 1303.950 904.890 1304.250 905.270 ;
        RECT 1376.845 905.270 1424.770 905.570 ;
        RECT 1376.845 905.255 1377.175 905.270 ;
        RECT 1424.470 904.890 1424.770 905.270 ;
        RECT 1462.190 904.890 1462.490 905.950 ;
        RECT 1496.190 905.940 1496.570 905.950 ;
        RECT 1497.110 905.570 1497.490 905.580 ;
        RECT 1545.205 905.570 1545.535 905.585 ;
        RECT 1497.110 905.270 1545.535 905.570 ;
        RECT 1497.110 905.260 1497.490 905.270 ;
        RECT 1545.205 905.255 1545.535 905.270 ;
        RECT 1560.385 905.570 1560.715 905.585 ;
        RECT 1587.310 905.570 1587.610 906.630 ;
        RECT 1634.905 906.615 1635.235 906.630 ;
        RECT 1786.910 906.250 1787.290 906.260 ;
        RECT 1752.910 905.950 1787.290 906.250 ;
        RECT 1560.385 905.270 1587.610 905.570 ;
        RECT 1634.905 905.570 1635.235 905.585 ;
        RECT 1634.905 905.270 1655.690 905.570 ;
        RECT 1560.385 905.255 1560.715 905.270 ;
        RECT 1634.905 905.255 1635.235 905.270 ;
        RECT 1303.950 904.590 1305.170 904.890 ;
        RECT 1424.470 904.590 1462.490 904.890 ;
        RECT 1655.390 904.890 1655.690 905.270 ;
        RECT 1752.910 904.890 1753.210 905.950 ;
        RECT 1786.910 905.940 1787.290 905.950 ;
        RECT 1883.550 905.950 1931.690 906.250 ;
        RECT 1883.550 904.890 1883.850 905.950 ;
        RECT 1655.390 904.590 1657.530 904.890 ;
        RECT 1207.310 903.910 1272.970 904.210 ;
        RECT 1304.870 904.210 1305.170 904.590 ;
        RECT 1352.465 904.210 1352.795 904.225 ;
        RECT 1304.870 903.910 1352.795 904.210 ;
        RECT 1657.230 904.210 1657.530 904.590 ;
        RECT 1714.270 904.590 1753.210 904.890 ;
        RECT 1849.510 904.590 1883.850 904.890 ;
        RECT 1714.270 904.210 1714.570 904.590 ;
        RECT 1657.230 904.040 1703.530 904.210 ;
        RECT 1704.150 904.040 1714.570 904.210 ;
        RECT 1657.230 903.910 1714.570 904.040 ;
        RECT 1810.625 904.210 1810.955 904.225 ;
        RECT 1849.510 904.210 1849.810 904.590 ;
        RECT 1810.625 903.910 1849.810 904.210 ;
        RECT 1931.390 904.210 1931.690 905.950 ;
        RECT 2138.390 905.270 2187.450 905.570 ;
        RECT 1992.325 904.890 1992.655 904.905 ;
        RECT 1946.110 904.590 1992.655 904.890 ;
        RECT 1946.110 904.210 1946.410 904.590 ;
        RECT 1992.325 904.575 1992.655 904.590 ;
        RECT 1995.085 904.890 1995.415 904.905 ;
        RECT 2089.385 904.890 2089.715 904.905 ;
        RECT 1995.085 904.590 2028.290 904.890 ;
        RECT 1995.085 904.575 1995.415 904.590 ;
        RECT 1931.390 903.910 1946.410 904.210 ;
        RECT 2027.990 904.210 2028.290 904.590 ;
        RECT 2042.710 904.590 2089.715 904.890 ;
        RECT 2042.710 904.210 2043.010 904.590 ;
        RECT 2089.385 904.575 2089.715 904.590 ;
        RECT 2091.685 904.890 2092.015 904.905 ;
        RECT 2091.685 904.590 2124.890 904.890 ;
        RECT 2091.685 904.575 2092.015 904.590 ;
        RECT 2027.990 903.910 2043.010 904.210 ;
        RECT 2124.590 904.210 2124.890 904.590 ;
        RECT 2138.390 904.210 2138.690 905.270 ;
        RECT 2124.590 903.910 2138.690 904.210 ;
        RECT 2187.150 904.210 2187.450 905.270 ;
        RECT 2380.350 905.270 2428.490 905.570 ;
        RECT 2272.005 904.890 2272.335 904.905 ;
        RECT 2235.910 904.590 2272.335 904.890 ;
        RECT 2235.910 904.210 2236.210 904.590 ;
        RECT 2272.005 904.575 2272.335 904.590 ;
        RECT 2291.785 904.890 2292.115 904.905 ;
        RECT 2291.785 904.590 2331.890 904.890 ;
        RECT 2291.785 904.575 2292.115 904.590 ;
        RECT 2187.150 903.910 2236.210 904.210 ;
        RECT 2331.590 904.210 2331.890 904.590 ;
        RECT 2380.350 904.210 2380.650 905.270 ;
        RECT 2331.590 903.910 2380.650 904.210 ;
        RECT 2428.190 904.210 2428.490 905.270 ;
        RECT 2476.950 905.270 2525.090 905.570 ;
        RECT 2476.950 904.210 2477.250 905.270 ;
        RECT 2428.190 903.910 2477.250 904.210 ;
        RECT 2524.790 904.210 2525.090 905.270 ;
        RECT 2573.550 905.270 2621.690 905.570 ;
        RECT 2573.550 904.210 2573.850 905.270 ;
        RECT 2524.790 903.910 2573.850 904.210 ;
        RECT 2621.390 904.210 2621.690 905.270 ;
        RECT 2642.550 905.270 2739.450 905.570 ;
        RECT 2642.550 904.210 2642.850 905.270 ;
        RECT 2739.150 904.890 2739.450 905.270 ;
        RECT 2787.910 905.270 2836.050 905.570 ;
        RECT 2739.150 904.590 2787.290 904.890 ;
        RECT 2621.390 903.910 2642.850 904.210 ;
        RECT 2786.990 904.210 2787.290 904.590 ;
        RECT 2787.910 904.210 2788.210 905.270 ;
        RECT 2835.750 904.890 2836.050 905.270 ;
        RECT 2916.710 904.890 2917.010 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 2835.750 904.590 2917.010 904.890 ;
        RECT 2786.990 903.910 2788.210 904.210 ;
        RECT 1207.310 903.900 1207.690 903.910 ;
        RECT 1352.465 903.895 1352.795 903.910 ;
        RECT 1703.230 903.740 1704.450 903.910 ;
        RECT 1810.625 903.895 1810.955 903.910 ;
      LAYER via3 ;
        RECT 1188.940 2814.700 1189.260 2815.020 ;
        RECT 1786.940 907.300 1787.260 907.620 ;
        RECT 1188.940 905.260 1189.260 905.580 ;
        RECT 1207.340 905.260 1207.660 905.580 ;
        RECT 1207.340 903.900 1207.660 904.220 ;
        RECT 1496.220 905.940 1496.540 906.260 ;
        RECT 1497.140 905.260 1497.460 905.580 ;
        RECT 1786.940 905.940 1787.260 906.260 ;
      LAYER met4 ;
        RECT 1188.935 2814.695 1189.265 2815.025 ;
        RECT 1188.950 905.585 1189.250 2814.695 ;
        RECT 1786.935 907.295 1787.265 907.625 ;
        RECT 1786.950 906.265 1787.250 907.295 ;
        RECT 1496.215 906.250 1496.545 906.265 ;
        RECT 1496.215 905.950 1497.450 906.250 ;
        RECT 1496.215 905.935 1496.545 905.950 ;
        RECT 1497.150 905.585 1497.450 905.950 ;
        RECT 1786.935 905.935 1787.265 906.265 ;
        RECT 1188.935 905.255 1189.265 905.585 ;
        RECT 1207.335 905.255 1207.665 905.585 ;
        RECT 1497.135 905.255 1497.465 905.585 ;
        RECT 1207.350 904.225 1207.650 905.255 ;
        RECT 1207.335 903.895 1207.665 904.225 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1439.025 2801.005 1439.195 2803.215 ;
        RECT 1860.845 2801.005 1861.475 2801.175 ;
      LAYER mcon ;
        RECT 1439.025 2803.045 1439.195 2803.215 ;
        RECT 1861.305 2801.005 1861.475 2801.175 ;
      LAYER met1 ;
        RECT 1278.870 2814.420 1279.190 2814.480 ;
        RECT 1434.810 2814.420 1435.130 2814.480 ;
        RECT 1278.870 2814.280 1435.130 2814.420 ;
        RECT 1278.870 2814.220 1279.190 2814.280 ;
        RECT 1434.810 2814.220 1435.130 2814.280 ;
        RECT 1434.810 2803.200 1435.130 2803.260 ;
        RECT 1438.965 2803.200 1439.255 2803.245 ;
        RECT 1434.810 2803.060 1439.255 2803.200 ;
        RECT 1434.810 2803.000 1435.130 2803.060 ;
        RECT 1438.965 2803.015 1439.255 2803.060 ;
        RECT 1438.965 2801.160 1439.255 2801.205 ;
        RECT 1860.785 2801.160 1861.075 2801.205 ;
        RECT 1438.965 2801.020 1861.075 2801.160 ;
        RECT 1438.965 2800.975 1439.255 2801.020 ;
        RECT 1860.785 2800.975 1861.075 2801.020 ;
        RECT 1861.245 2801.160 1861.535 2801.205 ;
        RECT 2001.070 2801.160 2001.390 2801.220 ;
        RECT 1861.245 2801.020 2001.390 2801.160 ;
        RECT 1861.245 2800.975 1861.535 2801.020 ;
        RECT 2001.070 2800.960 2001.390 2801.020 ;
        RECT 2002.910 2801.160 2003.230 2801.220 ;
        RECT 2898.990 2801.160 2899.310 2801.220 ;
        RECT 2002.910 2801.020 2899.310 2801.160 ;
        RECT 2002.910 2800.960 2003.230 2801.020 ;
        RECT 2898.990 2800.960 2899.310 2801.020 ;
        RECT 2898.990 2763.420 2899.310 2763.480 ;
        RECT 2904.050 2763.420 2904.370 2763.480 ;
        RECT 2898.990 2763.280 2904.370 2763.420 ;
        RECT 2898.990 2763.220 2899.310 2763.280 ;
        RECT 2904.050 2763.220 2904.370 2763.280 ;
      LAYER via ;
        RECT 1278.900 2814.220 1279.160 2814.480 ;
        RECT 1434.840 2814.220 1435.100 2814.480 ;
        RECT 1434.840 2803.000 1435.100 2803.260 ;
        RECT 2001.100 2800.960 2001.360 2801.220 ;
        RECT 2002.940 2800.960 2003.200 2801.220 ;
        RECT 2899.020 2800.960 2899.280 2801.220 ;
        RECT 2899.020 2763.220 2899.280 2763.480 ;
        RECT 2904.080 2763.220 2904.340 2763.480 ;
      LAYER met2 ;
        RECT 1278.900 2814.190 1279.160 2814.510 ;
        RECT 1434.840 2814.190 1435.100 2814.510 ;
        RECT 1278.960 2800.000 1279.100 2814.190 ;
        RECT 1434.900 2803.290 1435.040 2814.190 ;
        RECT 1434.840 2802.970 1435.100 2803.290 ;
        RECT 2001.090 2801.075 2001.370 2801.445 ;
        RECT 2002.930 2801.075 2003.210 2801.445 ;
        RECT 2001.100 2800.930 2001.360 2801.075 ;
        RECT 2002.940 2800.930 2003.200 2801.075 ;
        RECT 2899.020 2800.930 2899.280 2801.250 ;
        RECT 1278.825 2796.000 1279.105 2800.000 ;
        RECT 2899.080 2763.510 2899.220 2800.930 ;
        RECT 2899.020 2763.190 2899.280 2763.510 ;
        RECT 2904.080 2763.190 2904.340 2763.510 ;
        RECT 2904.140 1144.285 2904.280 2763.190 ;
        RECT 2904.070 1143.915 2904.350 1144.285 ;
      LAYER via2 ;
        RECT 2001.090 2801.120 2001.370 2801.400 ;
        RECT 2002.930 2801.120 2003.210 2801.400 ;
        RECT 2904.070 1143.960 2904.350 1144.240 ;
      LAYER met3 ;
        RECT 2001.065 2801.410 2001.395 2801.425 ;
        RECT 2002.905 2801.410 2003.235 2801.425 ;
        RECT 2001.065 2801.110 2003.235 2801.410 ;
        RECT 2001.065 2801.095 2001.395 2801.110 ;
        RECT 2002.905 2801.095 2003.235 2801.110 ;
        RECT 2904.045 1144.250 2904.375 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2904.045 1143.950 2924.800 1144.250 ;
        RECT 2904.045 1143.935 2904.375 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2001.605 2800.665 2002.695 2800.835 ;
      LAYER mcon ;
        RECT 2002.525 2800.665 2002.695 2800.835 ;
      LAYER met1 ;
        RECT 1307.850 2813.060 1308.170 2813.120 ;
        RECT 1393.870 2813.060 1394.190 2813.120 ;
        RECT 1307.850 2812.920 1394.190 2813.060 ;
        RECT 1307.850 2812.860 1308.170 2812.920 ;
        RECT 1393.870 2812.860 1394.190 2812.920 ;
        RECT 1393.870 2800.820 1394.190 2800.880 ;
        RECT 2001.545 2800.820 2001.835 2800.865 ;
        RECT 1393.870 2800.680 2001.835 2800.820 ;
        RECT 1393.870 2800.620 1394.190 2800.680 ;
        RECT 2001.545 2800.635 2001.835 2800.680 ;
        RECT 2002.465 2800.820 2002.755 2800.865 ;
        RECT 2900.370 2800.820 2900.690 2800.880 ;
        RECT 2002.465 2800.680 2900.690 2800.820 ;
        RECT 2002.465 2800.635 2002.755 2800.680 ;
        RECT 2900.370 2800.620 2900.690 2800.680 ;
      LAYER via ;
        RECT 1307.880 2812.860 1308.140 2813.120 ;
        RECT 1393.900 2812.860 1394.160 2813.120 ;
        RECT 1393.900 2800.620 1394.160 2800.880 ;
        RECT 2900.400 2800.620 2900.660 2800.880 ;
      LAYER met2 ;
        RECT 1307.880 2812.830 1308.140 2813.150 ;
        RECT 1393.900 2812.830 1394.160 2813.150 ;
        RECT 1307.940 2800.000 1308.080 2812.830 ;
        RECT 1393.960 2800.910 1394.100 2812.830 ;
        RECT 1393.900 2800.590 1394.160 2800.910 ;
        RECT 2900.400 2800.590 2900.660 2800.910 ;
        RECT 1307.805 2796.000 1308.085 2800.000 ;
        RECT 2900.460 1378.885 2900.600 2800.590 ;
        RECT 2900.390 1378.515 2900.670 1378.885 ;
      LAYER via2 ;
        RECT 2900.390 1378.560 2900.670 1378.840 ;
      LAYER met3 ;
        RECT 2900.365 1378.850 2900.695 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.365 1378.550 2924.800 1378.850 ;
        RECT 2900.365 1378.535 2900.695 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1860.845 2799.645 1863.775 2799.815 ;
      LAYER mcon ;
        RECT 1863.605 2799.645 1863.775 2799.815 ;
      LAYER met1 ;
        RECT 1338.210 2799.800 1338.530 2799.860 ;
        RECT 1860.785 2799.800 1861.075 2799.845 ;
        RECT 1338.210 2799.660 1861.075 2799.800 ;
        RECT 1338.210 2799.600 1338.530 2799.660 ;
        RECT 1860.785 2799.615 1861.075 2799.660 ;
        RECT 1863.545 2799.800 1863.835 2799.845 ;
        RECT 2001.070 2799.800 2001.390 2799.860 ;
        RECT 1863.545 2799.660 2001.390 2799.800 ;
        RECT 1863.545 2799.615 1863.835 2799.660 ;
        RECT 2001.070 2799.600 2001.390 2799.660 ;
        RECT 2002.910 2799.800 2003.230 2799.860 ;
        RECT 2887.950 2799.800 2888.270 2799.860 ;
        RECT 2002.910 2799.660 2888.270 2799.800 ;
        RECT 2002.910 2799.600 2003.230 2799.660 ;
        RECT 2887.950 2799.600 2888.270 2799.660 ;
        RECT 2887.950 1614.560 2888.270 1614.620 ;
        RECT 2899.450 1614.560 2899.770 1614.620 ;
        RECT 2887.950 1614.420 2899.770 1614.560 ;
        RECT 2887.950 1614.360 2888.270 1614.420 ;
        RECT 2899.450 1614.360 2899.770 1614.420 ;
      LAYER via ;
        RECT 1338.240 2799.600 1338.500 2799.860 ;
        RECT 2001.100 2799.600 2001.360 2799.860 ;
        RECT 2002.940 2799.600 2003.200 2799.860 ;
        RECT 2887.980 2799.600 2888.240 2799.860 ;
        RECT 2887.980 1614.360 2888.240 1614.620 ;
        RECT 2899.480 1614.360 2899.740 1614.620 ;
      LAYER met2 ;
        RECT 1336.785 2799.970 1337.065 2800.000 ;
        RECT 1336.785 2799.890 1338.440 2799.970 ;
        RECT 1336.785 2799.830 1338.500 2799.890 ;
        RECT 1336.785 2796.000 1337.065 2799.830 ;
        RECT 1338.240 2799.570 1338.500 2799.830 ;
        RECT 2001.090 2799.715 2001.370 2800.085 ;
        RECT 2002.930 2799.715 2003.210 2800.085 ;
        RECT 2001.100 2799.570 2001.360 2799.715 ;
        RECT 2002.940 2799.570 2003.200 2799.715 ;
        RECT 2887.980 2799.570 2888.240 2799.890 ;
        RECT 2888.040 1614.650 2888.180 2799.570 ;
        RECT 2887.980 1614.330 2888.240 1614.650 ;
        RECT 2899.480 1614.330 2899.740 1614.650 ;
        RECT 2899.540 1613.485 2899.680 1614.330 ;
        RECT 2899.470 1613.115 2899.750 1613.485 ;
      LAYER via2 ;
        RECT 2001.090 2799.760 2001.370 2800.040 ;
        RECT 2002.930 2799.760 2003.210 2800.040 ;
        RECT 2899.470 1613.160 2899.750 1613.440 ;
      LAYER met3 ;
        RECT 2001.065 2800.050 2001.395 2800.065 ;
        RECT 2002.905 2800.050 2003.235 2800.065 ;
        RECT 2001.065 2799.750 2003.235 2800.050 ;
        RECT 2001.065 2799.735 2001.395 2799.750 ;
        RECT 2002.905 2799.735 2003.235 2799.750 ;
        RECT 2899.445 1613.450 2899.775 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2899.445 1613.150 2924.800 1613.450 ;
        RECT 2899.445 1613.135 2899.775 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1365.810 2812.720 1366.130 2812.780 ;
        RECT 2253.150 2812.720 2253.470 2812.780 ;
        RECT 1365.810 2812.580 2253.470 2812.720 ;
        RECT 1365.810 2812.520 1366.130 2812.580 ;
        RECT 2253.150 2812.520 2253.470 2812.580 ;
        RECT 2253.150 1849.160 2253.470 1849.220 ;
        RECT 2898.990 1849.160 2899.310 1849.220 ;
        RECT 2253.150 1849.020 2899.310 1849.160 ;
        RECT 2253.150 1848.960 2253.470 1849.020 ;
        RECT 2898.990 1848.960 2899.310 1849.020 ;
      LAYER via ;
        RECT 1365.840 2812.520 1366.100 2812.780 ;
        RECT 2253.180 2812.520 2253.440 2812.780 ;
        RECT 2253.180 1848.960 2253.440 1849.220 ;
        RECT 2899.020 1848.960 2899.280 1849.220 ;
      LAYER met2 ;
        RECT 1365.840 2812.490 1366.100 2812.810 ;
        RECT 2253.180 2812.490 2253.440 2812.810 ;
        RECT 1365.900 2800.000 1366.040 2812.490 ;
        RECT 1365.765 2796.000 1366.045 2800.000 ;
        RECT 2253.240 1849.250 2253.380 2812.490 ;
        RECT 2253.180 1848.930 2253.440 1849.250 ;
        RECT 2899.020 1848.930 2899.280 1849.250 ;
        RECT 2899.080 1848.085 2899.220 1848.930 ;
        RECT 2899.010 1847.715 2899.290 1848.085 ;
      LAYER via2 ;
        RECT 2899.010 1847.760 2899.290 1848.040 ;
      LAYER met3 ;
        RECT 2898.985 1848.050 2899.315 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2898.985 1847.750 2924.800 1848.050 ;
        RECT 2898.985 1847.735 2899.315 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1394.790 2813.400 1395.110 2813.460 ;
        RECT 2254.990 2813.400 2255.310 2813.460 ;
        RECT 1394.790 2813.260 2255.310 2813.400 ;
        RECT 1394.790 2813.200 1395.110 2813.260 ;
        RECT 2254.990 2813.200 2255.310 2813.260 ;
        RECT 2254.070 2083.760 2254.390 2083.820 ;
        RECT 2898.990 2083.760 2899.310 2083.820 ;
        RECT 2254.070 2083.620 2899.310 2083.760 ;
        RECT 2254.070 2083.560 2254.390 2083.620 ;
        RECT 2898.990 2083.560 2899.310 2083.620 ;
      LAYER via ;
        RECT 1394.820 2813.200 1395.080 2813.460 ;
        RECT 2255.020 2813.200 2255.280 2813.460 ;
        RECT 2254.100 2083.560 2254.360 2083.820 ;
        RECT 2899.020 2083.560 2899.280 2083.820 ;
      LAYER met2 ;
        RECT 1394.820 2813.170 1395.080 2813.490 ;
        RECT 2255.020 2813.170 2255.280 2813.490 ;
        RECT 1394.880 2800.000 1395.020 2813.170 ;
        RECT 1394.745 2796.000 1395.025 2800.000 ;
        RECT 2255.080 2787.050 2255.220 2813.170 ;
        RECT 2254.160 2786.910 2255.220 2787.050 ;
        RECT 2254.160 2083.850 2254.300 2786.910 ;
        RECT 2254.100 2083.530 2254.360 2083.850 ;
        RECT 2899.020 2083.530 2899.280 2083.850 ;
        RECT 2899.080 2082.685 2899.220 2083.530 ;
        RECT 2899.010 2082.315 2899.290 2082.685 ;
      LAYER via2 ;
        RECT 2899.010 2082.360 2899.290 2082.640 ;
      LAYER met3 ;
        RECT 2898.985 2082.650 2899.315 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2898.985 2082.350 2924.800 2082.650 ;
        RECT 2898.985 2082.335 2899.315 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1423.770 2814.080 1424.090 2814.140 ;
        RECT 2255.450 2814.080 2255.770 2814.140 ;
        RECT 1423.770 2813.940 2255.770 2814.080 ;
        RECT 1423.770 2813.880 1424.090 2813.940 ;
        RECT 2255.450 2813.880 2255.770 2813.940 ;
        RECT 2254.990 2318.360 2255.310 2318.420 ;
        RECT 2898.990 2318.360 2899.310 2318.420 ;
        RECT 2254.990 2318.220 2899.310 2318.360 ;
        RECT 2254.990 2318.160 2255.310 2318.220 ;
        RECT 2898.990 2318.160 2899.310 2318.220 ;
      LAYER via ;
        RECT 1423.800 2813.880 1424.060 2814.140 ;
        RECT 2255.480 2813.880 2255.740 2814.140 ;
        RECT 2255.020 2318.160 2255.280 2318.420 ;
        RECT 2899.020 2318.160 2899.280 2318.420 ;
      LAYER met2 ;
        RECT 1423.800 2813.850 1424.060 2814.170 ;
        RECT 2255.480 2813.850 2255.740 2814.170 ;
        RECT 1423.860 2800.000 1424.000 2813.850 ;
        RECT 1423.725 2796.000 1424.005 2800.000 ;
        RECT 2255.540 2786.370 2255.680 2813.850 ;
        RECT 2255.080 2786.230 2255.680 2786.370 ;
        RECT 2255.080 2318.450 2255.220 2786.230 ;
        RECT 2255.020 2318.130 2255.280 2318.450 ;
        RECT 2899.020 2318.130 2899.280 2318.450 ;
        RECT 2899.080 2317.285 2899.220 2318.130 ;
        RECT 2899.010 2316.915 2899.290 2317.285 ;
      LAYER via2 ;
        RECT 2899.010 2316.960 2899.290 2317.240 ;
      LAYER met3 ;
        RECT 2898.985 2317.250 2899.315 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2898.985 2316.950 2924.800 2317.250 ;
        RECT 2898.985 2316.935 2899.315 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 146.100 1352.790 146.160 ;
        RECT 1369.950 146.100 1370.270 146.160 ;
        RECT 1352.470 145.960 1370.270 146.100 ;
        RECT 1352.470 145.900 1352.790 145.960 ;
        RECT 1369.950 145.900 1370.270 145.960 ;
        RECT 1992.330 146.100 1992.650 146.160 ;
        RECT 1995.090 146.100 1995.410 146.160 ;
        RECT 1992.330 145.960 1995.410 146.100 ;
        RECT 1992.330 145.900 1992.650 145.960 ;
        RECT 1995.090 145.900 1995.410 145.960 ;
        RECT 2380.110 146.100 2380.430 146.160 ;
        RECT 2414.610 146.100 2414.930 146.160 ;
        RECT 2380.110 145.960 2414.930 146.100 ;
        RECT 2380.110 145.900 2380.430 145.960 ;
        RECT 2414.610 145.900 2414.930 145.960 ;
        RECT 2089.390 145.760 2089.710 145.820 ;
        RECT 2090.770 145.760 2091.090 145.820 ;
        RECT 2089.390 145.620 2091.090 145.760 ;
        RECT 2089.390 145.560 2089.710 145.620 ;
        RECT 2090.770 145.560 2091.090 145.620 ;
        RECT 2221.870 145.420 2222.190 145.480 ;
        RECT 2246.250 145.420 2246.570 145.480 ;
        RECT 2221.870 145.280 2246.570 145.420 ;
        RECT 2221.870 145.220 2222.190 145.280 ;
        RECT 2246.250 145.220 2246.570 145.280 ;
      LAYER via ;
        RECT 1352.500 145.900 1352.760 146.160 ;
        RECT 1369.980 145.900 1370.240 146.160 ;
        RECT 1992.360 145.900 1992.620 146.160 ;
        RECT 1995.120 145.900 1995.380 146.160 ;
        RECT 2380.140 145.900 2380.400 146.160 ;
        RECT 2414.640 145.900 2414.900 146.160 ;
        RECT 2089.420 145.560 2089.680 145.820 ;
        RECT 2090.800 145.560 2091.060 145.820 ;
        RECT 2221.900 145.220 2222.160 145.480 ;
        RECT 2246.280 145.220 2246.540 145.480 ;
      LAYER met2 ;
        RECT 1172.565 2796.570 1172.845 2800.000 ;
        RECT 1173.090 2796.570 1173.370 2796.685 ;
        RECT 1172.565 2796.430 1173.370 2796.570 ;
        RECT 1172.565 2796.000 1172.845 2796.430 ;
        RECT 1173.090 2796.315 1173.370 2796.430 ;
        RECT 1193.330 162.675 1193.610 163.045 ;
        RECT 1193.400 146.045 1193.540 162.675 ;
        RECT 1459.210 147.715 1459.490 148.085 ;
        RECT 1628.030 147.715 1628.310 148.085 ;
        RECT 1248.530 146.355 1248.810 146.725 ;
        RECT 1369.970 146.355 1370.250 146.725 ;
        RECT 1424.710 146.355 1424.990 146.725 ;
        RECT 1193.330 145.675 1193.610 146.045 ;
        RECT 1248.600 144.685 1248.740 146.355 ;
        RECT 1370.040 146.190 1370.180 146.355 ;
        RECT 1352.500 146.045 1352.760 146.190 ;
        RECT 1352.490 145.675 1352.770 146.045 ;
        RECT 1369.980 145.870 1370.240 146.190 ;
        RECT 1424.780 145.365 1424.920 146.355 ;
        RECT 1459.280 145.365 1459.420 147.715 ;
        RECT 1531.430 147.035 1531.710 147.405 ;
        RECT 1531.500 146.045 1531.640 147.035 ;
        RECT 1628.100 146.725 1628.240 147.715 ;
        RECT 2359.430 147.035 2359.710 147.405 ;
        RECT 1628.030 146.355 1628.310 146.725 ;
        RECT 2246.270 146.355 2246.550 146.725 ;
        RECT 1992.360 146.045 1992.620 146.190 ;
        RECT 1995.120 146.045 1995.380 146.190 ;
        RECT 1531.430 145.675 1531.710 146.045 ;
        RECT 1579.730 145.675 1580.010 146.045 ;
        RECT 1992.350 145.675 1992.630 146.045 ;
        RECT 1995.110 145.675 1995.390 146.045 ;
        RECT 2089.410 145.675 2089.690 146.045 ;
        RECT 2090.790 145.675 2091.070 146.045 ;
        RECT 1579.800 145.365 1579.940 145.675 ;
        RECT 2089.420 145.530 2089.680 145.675 ;
        RECT 2090.800 145.530 2091.060 145.675 ;
        RECT 2246.340 145.510 2246.480 146.355 ;
        RECT 2221.900 145.365 2222.160 145.510 ;
        RECT 1424.710 144.995 1424.990 145.365 ;
        RECT 1459.210 144.995 1459.490 145.365 ;
        RECT 1579.730 144.995 1580.010 145.365 ;
        RECT 2221.890 144.995 2222.170 145.365 ;
        RECT 2246.280 145.190 2246.540 145.510 ;
        RECT 2359.500 145.365 2359.640 147.035 ;
        RECT 2414.630 146.355 2414.910 146.725 ;
        RECT 2414.700 146.190 2414.840 146.355 ;
        RECT 2380.140 146.045 2380.400 146.190 ;
        RECT 2380.130 145.675 2380.410 146.045 ;
        RECT 2414.640 145.870 2414.900 146.190 ;
        RECT 2359.430 144.995 2359.710 145.365 ;
        RECT 1248.530 144.315 1248.810 144.685 ;
      LAYER via2 ;
        RECT 1173.090 2796.360 1173.370 2796.640 ;
        RECT 1193.330 162.720 1193.610 163.000 ;
        RECT 1459.210 147.760 1459.490 148.040 ;
        RECT 1628.030 147.760 1628.310 148.040 ;
        RECT 1248.530 146.400 1248.810 146.680 ;
        RECT 1369.970 146.400 1370.250 146.680 ;
        RECT 1424.710 146.400 1424.990 146.680 ;
        RECT 1193.330 145.720 1193.610 146.000 ;
        RECT 1352.490 145.720 1352.770 146.000 ;
        RECT 1531.430 147.080 1531.710 147.360 ;
        RECT 2359.430 147.080 2359.710 147.360 ;
        RECT 1628.030 146.400 1628.310 146.680 ;
        RECT 2246.270 146.400 2246.550 146.680 ;
        RECT 1531.430 145.720 1531.710 146.000 ;
        RECT 1579.730 145.720 1580.010 146.000 ;
        RECT 1992.350 145.720 1992.630 146.000 ;
        RECT 1995.110 145.720 1995.390 146.000 ;
        RECT 2089.410 145.720 2089.690 146.000 ;
        RECT 2090.790 145.720 2091.070 146.000 ;
        RECT 1424.710 145.040 1424.990 145.320 ;
        RECT 1459.210 145.040 1459.490 145.320 ;
        RECT 1579.730 145.040 1580.010 145.320 ;
        RECT 2221.890 145.040 2222.170 145.320 ;
        RECT 2414.630 146.400 2414.910 146.680 ;
        RECT 2380.130 145.720 2380.410 146.000 ;
        RECT 2359.430 145.040 2359.710 145.320 ;
        RECT 1248.530 144.360 1248.810 144.640 ;
      LAYER met3 ;
        RECT 1171.430 2796.650 1171.810 2796.660 ;
        RECT 1173.065 2796.650 1173.395 2796.665 ;
        RECT 1171.430 2796.350 1173.395 2796.650 ;
        RECT 1171.430 2796.340 1171.810 2796.350 ;
        RECT 1173.065 2796.335 1173.395 2796.350 ;
        RECT 1172.350 163.010 1172.730 163.020 ;
        RECT 1193.305 163.010 1193.635 163.025 ;
        RECT 1172.350 162.710 1193.635 163.010 ;
        RECT 1172.350 162.700 1172.730 162.710 ;
        RECT 1193.305 162.695 1193.635 162.710 ;
        RECT 1459.185 148.050 1459.515 148.065 ;
        RECT 1579.910 148.050 1580.290 148.060 ;
        RECT 1628.005 148.050 1628.335 148.065 ;
        RECT 1459.185 147.750 1483.650 148.050 ;
        RECT 1459.185 147.735 1459.515 147.750 ;
        RECT 1483.350 147.370 1483.650 147.750 ;
        RECT 1579.910 147.750 1628.335 148.050 ;
        RECT 1579.910 147.740 1580.290 147.750 ;
        RECT 1628.005 147.735 1628.335 147.750 ;
        RECT 1531.405 147.370 1531.735 147.385 ;
        RECT 2311.310 147.370 2311.690 147.380 ;
        RECT 2359.405 147.370 2359.735 147.385 ;
        RECT 1248.750 147.070 1318.970 147.370 ;
        RECT 1483.350 147.070 1531.735 147.370 ;
        RECT 1248.750 146.705 1249.050 147.070 ;
        RECT 1248.505 146.690 1249.050 146.705 ;
        RECT 1248.100 146.390 1249.050 146.690 ;
        RECT 1248.505 146.375 1248.835 146.390 ;
        RECT 1193.305 146.010 1193.635 146.025 ;
        RECT 1318.670 146.010 1318.970 147.070 ;
        RECT 1531.405 147.055 1531.735 147.070 ;
        RECT 1752.910 147.070 1800.130 147.370 ;
        RECT 1369.945 146.690 1370.275 146.705 ;
        RECT 1424.685 146.690 1425.015 146.705 ;
        RECT 1369.945 146.390 1425.015 146.690 ;
        RECT 1369.945 146.375 1370.275 146.390 ;
        RECT 1424.685 146.375 1425.015 146.390 ;
        RECT 1628.005 146.690 1628.335 146.705 ;
        RECT 1628.005 146.390 1635.450 146.690 ;
        RECT 1628.005 146.375 1628.335 146.390 ;
        RECT 1352.465 146.010 1352.795 146.025 ;
        RECT 1193.305 145.710 1201.210 146.010 ;
        RECT 1318.670 145.710 1352.795 146.010 ;
        RECT 1193.305 145.695 1193.635 145.710 ;
        RECT 1200.910 144.650 1201.210 145.710 ;
        RECT 1352.465 145.695 1352.795 145.710 ;
        RECT 1531.405 146.010 1531.735 146.025 ;
        RECT 1579.705 146.020 1580.035 146.025 ;
        RECT 1635.150 146.020 1635.450 146.390 ;
        RECT 1579.705 146.010 1580.290 146.020 ;
        RECT 1531.405 145.710 1532.410 146.010 ;
        RECT 1531.405 145.695 1531.735 145.710 ;
        RECT 1424.685 145.330 1425.015 145.345 ;
        RECT 1459.185 145.330 1459.515 145.345 ;
        RECT 1424.685 145.030 1459.515 145.330 ;
        RECT 1532.110 145.330 1532.410 145.710 ;
        RECT 1579.705 145.710 1580.670 146.010 ;
        RECT 1579.705 145.700 1580.290 145.710 ;
        RECT 1635.110 145.700 1635.490 146.020 ;
        RECT 1636.030 146.010 1636.410 146.020 ;
        RECT 1752.910 146.010 1753.210 147.070 ;
        RECT 1636.030 145.710 1753.210 146.010 ;
        RECT 1799.830 146.010 1800.130 147.070 ;
        RECT 1883.550 147.070 1931.690 147.370 ;
        RECT 1834.750 146.690 1835.130 146.700 ;
        RECT 1801.670 146.390 1835.130 146.690 ;
        RECT 1801.670 146.010 1801.970 146.390 ;
        RECT 1834.750 146.380 1835.130 146.390 ;
        RECT 1883.550 146.010 1883.850 147.070 ;
        RECT 1799.830 145.710 1801.970 146.010 ;
        RECT 1849.510 145.710 1883.850 146.010 ;
        RECT 1636.030 145.700 1636.410 145.710 ;
        RECT 1579.705 145.695 1580.035 145.700 ;
        RECT 1579.705 145.330 1580.035 145.345 ;
        RECT 1532.110 145.030 1580.035 145.330 ;
        RECT 1424.685 145.015 1425.015 145.030 ;
        RECT 1459.185 145.015 1459.515 145.030 ;
        RECT 1579.705 145.015 1580.035 145.030 ;
        RECT 1834.750 145.330 1835.130 145.340 ;
        RECT 1849.510 145.330 1849.810 145.710 ;
        RECT 1834.750 145.030 1849.810 145.330 ;
        RECT 1931.390 145.330 1931.690 147.070 ;
        RECT 2311.310 147.070 2359.735 147.370 ;
        RECT 2311.310 147.060 2311.690 147.070 ;
        RECT 2359.405 147.055 2359.735 147.070 ;
        RECT 2246.245 146.690 2246.575 146.705 ;
        RECT 2414.605 146.690 2414.935 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2138.390 146.390 2187.450 146.690 ;
        RECT 1992.325 146.010 1992.655 146.025 ;
        RECT 1946.110 145.710 1992.655 146.010 ;
        RECT 1946.110 145.330 1946.410 145.710 ;
        RECT 1992.325 145.695 1992.655 145.710 ;
        RECT 1995.085 146.010 1995.415 146.025 ;
        RECT 2089.385 146.010 2089.715 146.025 ;
        RECT 1995.085 145.710 2028.290 146.010 ;
        RECT 1995.085 145.695 1995.415 145.710 ;
        RECT 1931.390 145.030 1946.410 145.330 ;
        RECT 2027.990 145.330 2028.290 145.710 ;
        RECT 2042.710 145.710 2089.715 146.010 ;
        RECT 2042.710 145.330 2043.010 145.710 ;
        RECT 2089.385 145.695 2089.715 145.710 ;
        RECT 2090.765 146.010 2091.095 146.025 ;
        RECT 2090.765 145.710 2124.890 146.010 ;
        RECT 2090.765 145.695 2091.095 145.710 ;
        RECT 2027.990 145.030 2043.010 145.330 ;
        RECT 2124.590 145.330 2124.890 145.710 ;
        RECT 2138.390 145.330 2138.690 146.390 ;
        RECT 2124.590 145.030 2138.690 145.330 ;
        RECT 2187.150 145.330 2187.450 146.390 ;
        RECT 2246.245 146.390 2294.170 146.690 ;
        RECT 2246.245 146.375 2246.575 146.390 ;
        RECT 2293.870 146.010 2294.170 146.390 ;
        RECT 2414.605 146.390 2449.650 146.690 ;
        RECT 2414.605 146.375 2414.935 146.390 ;
        RECT 2311.310 146.010 2311.690 146.020 ;
        RECT 2380.105 146.010 2380.435 146.025 ;
        RECT 2293.870 145.710 2311.690 146.010 ;
        RECT 2311.310 145.700 2311.690 145.710 ;
        RECT 2366.550 145.710 2380.435 146.010 ;
        RECT 2449.350 146.010 2449.650 146.390 ;
        RECT 2498.110 146.390 2546.250 146.690 ;
        RECT 2449.350 145.710 2497.490 146.010 ;
        RECT 2221.865 145.330 2222.195 145.345 ;
        RECT 2187.150 145.030 2222.195 145.330 ;
        RECT 1834.750 145.020 1835.130 145.030 ;
        RECT 2221.865 145.015 2222.195 145.030 ;
        RECT 2359.405 145.330 2359.735 145.345 ;
        RECT 2366.550 145.330 2366.850 145.710 ;
        RECT 2380.105 145.695 2380.435 145.710 ;
        RECT 2359.405 145.030 2366.850 145.330 ;
        RECT 2497.190 145.330 2497.490 145.710 ;
        RECT 2498.110 145.330 2498.410 146.390 ;
        RECT 2545.950 146.010 2546.250 146.390 ;
        RECT 2594.710 146.390 2642.850 146.690 ;
        RECT 2545.950 145.710 2594.090 146.010 ;
        RECT 2497.190 145.030 2498.410 145.330 ;
        RECT 2593.790 145.330 2594.090 145.710 ;
        RECT 2594.710 145.330 2595.010 146.390 ;
        RECT 2642.550 146.010 2642.850 146.390 ;
        RECT 2691.310 146.390 2739.450 146.690 ;
        RECT 2642.550 145.710 2690.690 146.010 ;
        RECT 2593.790 145.030 2595.010 145.330 ;
        RECT 2690.390 145.330 2690.690 145.710 ;
        RECT 2691.310 145.330 2691.610 146.390 ;
        RECT 2739.150 146.010 2739.450 146.390 ;
        RECT 2787.910 146.390 2836.050 146.690 ;
        RECT 2739.150 145.710 2787.290 146.010 ;
        RECT 2690.390 145.030 2691.610 145.330 ;
        RECT 2786.990 145.330 2787.290 145.710 ;
        RECT 2787.910 145.330 2788.210 146.390 ;
        RECT 2835.750 146.010 2836.050 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 146.010 2917.010 146.390 ;
        RECT 2835.750 145.710 2883.890 146.010 ;
        RECT 2786.990 145.030 2788.210 145.330 ;
        RECT 2883.590 145.330 2883.890 145.710 ;
        RECT 2884.510 145.710 2917.010 146.010 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2884.510 145.330 2884.810 145.710 ;
        RECT 2883.590 145.030 2884.810 145.330 ;
        RECT 2359.405 145.015 2359.735 145.030 ;
        RECT 1248.505 144.650 1248.835 144.665 ;
        RECT 1200.910 144.350 1248.835 144.650 ;
        RECT 1248.505 144.335 1248.835 144.350 ;
      LAYER via3 ;
        RECT 1171.460 2796.340 1171.780 2796.660 ;
        RECT 1172.380 162.700 1172.700 163.020 ;
        RECT 1579.940 147.740 1580.260 148.060 ;
        RECT 1579.940 145.700 1580.260 146.020 ;
        RECT 1635.140 145.700 1635.460 146.020 ;
        RECT 1636.060 145.700 1636.380 146.020 ;
        RECT 1834.780 146.380 1835.100 146.700 ;
        RECT 1834.780 145.020 1835.100 145.340 ;
        RECT 2311.340 147.060 2311.660 147.380 ;
        RECT 2311.340 145.700 2311.660 146.020 ;
      LAYER met4 ;
        RECT 1171.455 2796.650 1171.785 2796.665 ;
        RECT 1171.455 2796.350 1172.690 2796.650 ;
        RECT 1171.455 2796.335 1171.785 2796.350 ;
        RECT 1172.390 163.025 1172.690 2796.350 ;
        RECT 1172.375 162.695 1172.705 163.025 ;
        RECT 1579.935 147.735 1580.265 148.065 ;
        RECT 1579.950 146.025 1580.250 147.735 ;
        RECT 2311.335 147.055 2311.665 147.385 ;
        RECT 1834.775 146.375 1835.105 146.705 ;
        RECT 1579.935 145.695 1580.265 146.025 ;
        RECT 1635.135 145.695 1635.465 146.025 ;
        RECT 1636.055 145.695 1636.385 146.025 ;
        RECT 1635.150 144.650 1635.450 145.695 ;
        RECT 1636.070 144.650 1636.370 145.695 ;
        RECT 1834.790 145.345 1835.090 146.375 ;
        RECT 2311.350 146.025 2311.650 147.055 ;
        RECT 2311.335 145.695 2311.665 146.025 ;
        RECT 1834.775 145.015 1835.105 145.345 ;
        RECT 1635.150 144.350 1636.370 144.650 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1462.410 2814.420 1462.730 2814.480 ;
        RECT 2251.770 2814.420 2252.090 2814.480 ;
        RECT 1462.410 2814.280 2252.090 2814.420 ;
        RECT 1462.410 2814.220 1462.730 2814.280 ;
        RECT 2251.770 2814.220 2252.090 2814.280 ;
        RECT 2251.770 2785.860 2252.090 2785.920 ;
        RECT 2255.450 2785.860 2255.770 2785.920 ;
        RECT 2251.770 2785.720 2255.770 2785.860 ;
        RECT 2251.770 2785.660 2252.090 2785.720 ;
        RECT 2255.450 2785.660 2255.770 2785.720 ;
        RECT 2255.450 2497.540 2255.770 2497.600 ;
        RECT 2898.990 2497.540 2899.310 2497.600 ;
        RECT 2255.450 2497.400 2899.310 2497.540 ;
        RECT 2255.450 2497.340 2255.770 2497.400 ;
        RECT 2898.990 2497.340 2899.310 2497.400 ;
      LAYER via ;
        RECT 1462.440 2814.220 1462.700 2814.480 ;
        RECT 2251.800 2814.220 2252.060 2814.480 ;
        RECT 2251.800 2785.660 2252.060 2785.920 ;
        RECT 2255.480 2785.660 2255.740 2785.920 ;
        RECT 2255.480 2497.340 2255.740 2497.600 ;
        RECT 2899.020 2497.340 2899.280 2497.600 ;
      LAYER met2 ;
        RECT 1462.440 2814.190 1462.700 2814.510 ;
        RECT 2251.800 2814.190 2252.060 2814.510 ;
        RECT 1462.500 2800.000 1462.640 2814.190 ;
        RECT 1462.365 2796.000 1462.645 2800.000 ;
        RECT 2251.860 2785.950 2252.000 2814.190 ;
        RECT 2251.800 2785.630 2252.060 2785.950 ;
        RECT 2255.480 2785.630 2255.740 2785.950 ;
        RECT 2255.540 2497.630 2255.680 2785.630 ;
        RECT 2255.480 2497.310 2255.740 2497.630 ;
        RECT 2899.020 2497.310 2899.280 2497.630 ;
        RECT 2899.080 2493.405 2899.220 2497.310 ;
        RECT 2899.010 2493.035 2899.290 2493.405 ;
      LAYER via2 ;
        RECT 2899.010 2493.080 2899.290 2493.360 ;
      LAYER met3 ;
        RECT 2898.985 2493.370 2899.315 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2898.985 2493.070 2924.800 2493.370 ;
        RECT 2898.985 2493.055 2899.315 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1519.985 2814.605 1520.155 2815.455 ;
        RECT 1534.705 2814.775 1534.875 2815.115 ;
        RECT 1534.705 2814.605 1535.795 2814.775 ;
        RECT 1552.185 2814.605 1559.255 2814.775 ;
      LAYER mcon ;
        RECT 1519.985 2815.285 1520.155 2815.455 ;
        RECT 1534.705 2814.945 1534.875 2815.115 ;
        RECT 1535.625 2814.605 1535.795 2814.775 ;
        RECT 1559.085 2814.605 1559.255 2814.775 ;
      LAYER met1 ;
        RECT 1519.925 2815.440 1520.215 2815.485 ;
        RECT 1519.925 2815.300 1525.200 2815.440 ;
        RECT 1519.925 2815.255 1520.215 2815.300 ;
        RECT 1525.060 2815.100 1525.200 2815.300 ;
        RECT 1534.645 2815.100 1534.935 2815.145 ;
        RECT 1525.060 2814.960 1534.935 2815.100 ;
        RECT 1534.645 2814.915 1534.935 2814.960 ;
        RECT 1491.390 2814.760 1491.710 2814.820 ;
        RECT 1519.925 2814.760 1520.215 2814.805 ;
        RECT 1491.390 2814.620 1520.215 2814.760 ;
        RECT 1491.390 2814.560 1491.710 2814.620 ;
        RECT 1519.925 2814.575 1520.215 2814.620 ;
        RECT 1535.565 2814.760 1535.855 2814.805 ;
        RECT 1552.125 2814.760 1552.415 2814.805 ;
        RECT 1535.565 2814.620 1552.415 2814.760 ;
        RECT 1535.565 2814.575 1535.855 2814.620 ;
        RECT 1552.125 2814.575 1552.415 2814.620 ;
        RECT 1559.025 2814.760 1559.315 2814.805 ;
        RECT 2252.230 2814.760 2252.550 2814.820 ;
        RECT 1559.025 2814.620 2252.550 2814.760 ;
        RECT 1559.025 2814.575 1559.315 2814.620 ;
        RECT 2252.230 2814.560 2252.550 2814.620 ;
        RECT 2252.230 2732.140 2252.550 2732.200 ;
        RECT 2898.990 2732.140 2899.310 2732.200 ;
        RECT 2252.230 2732.000 2899.310 2732.140 ;
        RECT 2252.230 2731.940 2252.550 2732.000 ;
        RECT 2898.990 2731.940 2899.310 2732.000 ;
      LAYER via ;
        RECT 1491.420 2814.560 1491.680 2814.820 ;
        RECT 2252.260 2814.560 2252.520 2814.820 ;
        RECT 2252.260 2731.940 2252.520 2732.200 ;
        RECT 2899.020 2731.940 2899.280 2732.200 ;
      LAYER met2 ;
        RECT 1491.420 2814.530 1491.680 2814.850 ;
        RECT 2252.260 2814.530 2252.520 2814.850 ;
        RECT 1491.480 2800.000 1491.620 2814.530 ;
        RECT 1491.345 2796.000 1491.625 2800.000 ;
        RECT 2252.320 2732.230 2252.460 2814.530 ;
        RECT 2252.260 2731.910 2252.520 2732.230 ;
        RECT 2899.020 2731.910 2899.280 2732.230 ;
        RECT 2899.080 2728.005 2899.220 2731.910 ;
        RECT 2899.010 2727.635 2899.290 2728.005 ;
      LAYER via2 ;
        RECT 2899.010 2727.680 2899.290 2727.960 ;
      LAYER met3 ;
        RECT 2898.985 2727.970 2899.315 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2898.985 2727.670 2924.800 2727.970 ;
        RECT 2898.985 2727.655 2899.315 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.510 2960.280 1524.830 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1524.510 2960.140 2901.150 2960.280 ;
        RECT 1524.510 2960.080 1524.830 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 1524.540 2960.080 1524.800 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1524.540 2960.050 1524.800 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1524.600 2801.330 1524.740 2960.050 ;
        RECT 1522.760 2801.190 1524.740 2801.330 ;
        RECT 1520.325 2799.970 1520.605 2800.000 ;
        RECT 1522.760 2799.970 1522.900 2801.190 ;
        RECT 1520.325 2799.830 1522.900 2799.970 ;
        RECT 1520.325 2796.000 1520.605 2799.830 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.110 3194.880 1552.430 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 1552.110 3194.740 2901.150 3194.880 ;
        RECT 1552.110 3194.680 1552.430 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
        RECT 1545.670 2825.640 1545.990 2825.700 ;
        RECT 1552.110 2825.640 1552.430 2825.700 ;
        RECT 1545.670 2825.500 1552.430 2825.640 ;
        RECT 1545.670 2825.440 1545.990 2825.500 ;
        RECT 1552.110 2825.440 1552.430 2825.500 ;
      LAYER via ;
        RECT 1552.140 3194.680 1552.400 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
        RECT 1545.700 2825.440 1545.960 2825.700 ;
        RECT 1552.140 2825.440 1552.400 2825.700 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 1552.140 3194.650 1552.400 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 1552.200 2825.730 1552.340 3194.650 ;
        RECT 1545.700 2825.410 1545.960 2825.730 ;
        RECT 1552.140 2825.410 1552.400 2825.730 ;
        RECT 1545.760 2800.650 1545.900 2825.410 ;
        RECT 1545.760 2800.510 1547.280 2800.650 ;
        RECT 1547.140 2799.970 1547.280 2800.510 ;
        RECT 1548.845 2799.970 1549.125 2800.000 ;
        RECT 1547.140 2799.830 1549.125 2799.970 ;
        RECT 1548.845 2796.000 1549.125 2799.830 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 1579.710 3429.480 1580.030 3429.540 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1579.710 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 2149.740 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 1579.710 3429.280 1580.030 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 1573.270 2825.640 1573.590 2825.700 ;
        RECT 1579.710 2825.640 1580.030 2825.700 ;
        RECT 1573.270 2825.500 1580.030 2825.640 ;
        RECT 1573.270 2825.440 1573.590 2825.500 ;
        RECT 1579.710 2825.440 1580.030 2825.500 ;
      LAYER via ;
        RECT 1579.740 3429.280 1580.000 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 1573.300 2825.440 1573.560 2825.700 ;
        RECT 1579.740 2825.440 1580.000 2825.700 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1579.740 3429.250 1580.000 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1579.800 2825.730 1579.940 3429.250 ;
        RECT 1573.300 2825.410 1573.560 2825.730 ;
        RECT 1579.740 2825.410 1580.000 2825.730 ;
        RECT 1573.360 2800.650 1573.500 2825.410 ;
        RECT 1573.360 2800.510 1576.260 2800.650 ;
        RECT 1576.120 2799.970 1576.260 2800.510 ;
        RECT 1577.825 2799.970 1578.105 2800.000 ;
        RECT 1576.120 2799.830 1578.105 2799.970 ;
        RECT 1577.825 2796.000 1578.105 2799.830 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 3503.260 1607.630 3503.320 ;
        RECT 2717.290 3503.260 2717.610 3503.320 ;
        RECT 1607.310 3503.120 2717.610 3503.260 ;
        RECT 1607.310 3503.060 1607.630 3503.120 ;
        RECT 2717.290 3503.060 2717.610 3503.120 ;
      LAYER via ;
        RECT 1607.340 3503.060 1607.600 3503.320 ;
        RECT 2717.320 3503.060 2717.580 3503.320 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3503.350 2717.520 3517.600 ;
        RECT 1607.340 3503.030 1607.600 3503.350 ;
        RECT 2717.320 3503.030 2717.580 3503.350 ;
        RECT 1606.805 2799.970 1607.085 2800.000 ;
        RECT 1607.400 2799.970 1607.540 3503.030 ;
        RECT 1606.805 2799.830 1607.540 2799.970 ;
        RECT 1606.805 2796.000 1607.085 2799.830 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1641.810 3504.960 1642.130 3505.020 ;
        RECT 2392.530 3504.960 2392.850 3505.020 ;
        RECT 1641.810 3504.820 2392.850 3504.960 ;
        RECT 1641.810 3504.760 1642.130 3504.820 ;
        RECT 2392.530 3504.760 2392.850 3504.820 ;
        RECT 1635.370 2825.640 1635.690 2825.700 ;
        RECT 1641.810 2825.640 1642.130 2825.700 ;
        RECT 1635.370 2825.500 1642.130 2825.640 ;
        RECT 1635.370 2825.440 1635.690 2825.500 ;
        RECT 1641.810 2825.440 1642.130 2825.500 ;
      LAYER via ;
        RECT 1641.840 3504.760 1642.100 3505.020 ;
        RECT 2392.560 3504.760 2392.820 3505.020 ;
        RECT 1635.400 2825.440 1635.660 2825.700 ;
        RECT 1641.840 2825.440 1642.100 2825.700 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3505.050 2392.760 3517.600 ;
        RECT 1641.840 3504.730 1642.100 3505.050 ;
        RECT 2392.560 3504.730 2392.820 3505.050 ;
        RECT 1641.900 2825.730 1642.040 3504.730 ;
        RECT 1635.400 2825.410 1635.660 2825.730 ;
        RECT 1641.840 2825.410 1642.100 2825.730 ;
        RECT 1635.460 2799.970 1635.600 2825.410 ;
        RECT 1635.785 2799.970 1636.065 2800.000 ;
        RECT 1635.460 2799.830 1636.065 2799.970 ;
        RECT 1635.785 2796.000 1636.065 2799.830 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1669.410 3499.860 1669.730 3499.920 ;
        RECT 2068.230 3499.860 2068.550 3499.920 ;
        RECT 1669.410 3499.720 2068.550 3499.860 ;
        RECT 1669.410 3499.660 1669.730 3499.720 ;
        RECT 2068.230 3499.660 2068.550 3499.720 ;
        RECT 1662.970 2825.640 1663.290 2825.700 ;
        RECT 1669.410 2825.640 1669.730 2825.700 ;
        RECT 1662.970 2825.500 1669.730 2825.640 ;
        RECT 1662.970 2825.440 1663.290 2825.500 ;
        RECT 1669.410 2825.440 1669.730 2825.500 ;
      LAYER via ;
        RECT 1669.440 3499.660 1669.700 3499.920 ;
        RECT 2068.260 3499.660 2068.520 3499.920 ;
        RECT 1663.000 2825.440 1663.260 2825.700 ;
        RECT 1669.440 2825.440 1669.700 2825.700 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3499.950 2068.460 3517.600 ;
        RECT 1669.440 3499.630 1669.700 3499.950 ;
        RECT 2068.260 3499.630 2068.520 3499.950 ;
        RECT 1669.500 2825.730 1669.640 3499.630 ;
        RECT 1663.000 2825.410 1663.260 2825.730 ;
        RECT 1669.440 2825.410 1669.700 2825.730 ;
        RECT 1663.060 2799.970 1663.200 2825.410 ;
        RECT 1664.765 2799.970 1665.045 2800.000 ;
        RECT 1663.060 2799.830 1665.045 2799.970 ;
        RECT 1664.765 2796.000 1665.045 2799.830 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1697.010 3498.500 1697.330 3498.560 ;
        RECT 1743.930 3498.500 1744.250 3498.560 ;
        RECT 1697.010 3498.360 1744.250 3498.500 ;
        RECT 1697.010 3498.300 1697.330 3498.360 ;
        RECT 1743.930 3498.300 1744.250 3498.360 ;
      LAYER via ;
        RECT 1697.040 3498.300 1697.300 3498.560 ;
        RECT 1743.960 3498.300 1744.220 3498.560 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3498.590 1744.160 3517.600 ;
        RECT 1697.040 3498.270 1697.300 3498.590 ;
        RECT 1743.960 3498.270 1744.220 3498.590 ;
        RECT 1697.100 2800.650 1697.240 3498.270 ;
        RECT 1695.260 2800.510 1697.240 2800.650 ;
        RECT 1693.745 2799.970 1694.025 2800.000 ;
        RECT 1695.260 2799.970 1695.400 2800.510 ;
        RECT 1693.745 2799.830 1695.400 2799.970 ;
        RECT 1693.745 2796.000 1694.025 2799.830 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3498.840 1419.490 3498.900 ;
        RECT 1718.170 3498.840 1718.490 3498.900 ;
        RECT 1419.170 3498.700 1718.490 3498.840 ;
        RECT 1419.170 3498.640 1419.490 3498.700 ;
        RECT 1718.170 3498.640 1718.490 3498.700 ;
      LAYER via ;
        RECT 1419.200 3498.640 1419.460 3498.900 ;
        RECT 1718.200 3498.640 1718.460 3498.900 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3498.930 1419.400 3517.600 ;
        RECT 1419.200 3498.610 1419.460 3498.930 ;
        RECT 1718.200 3498.610 1718.460 3498.930 ;
        RECT 1718.260 2801.330 1718.400 3498.610 ;
        RECT 1718.260 2801.190 1721.160 2801.330 ;
        RECT 1721.020 2799.970 1721.160 2801.190 ;
        RECT 1722.725 2799.970 1723.005 2800.000 ;
        RECT 1721.020 2799.830 1723.005 2799.970 ;
        RECT 1722.725 2796.000 1723.005 2799.830 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1202.970 2797.420 1203.290 2797.480 ;
        RECT 2901.290 2797.420 2901.610 2797.480 ;
        RECT 1202.970 2797.280 2901.610 2797.420 ;
        RECT 1202.970 2797.220 1203.290 2797.280 ;
        RECT 2901.290 2797.220 2901.610 2797.280 ;
      LAYER via ;
        RECT 1203.000 2797.220 1203.260 2797.480 ;
        RECT 2901.320 2797.220 2901.580 2797.480 ;
      LAYER met2 ;
        RECT 1201.545 2797.250 1201.825 2800.000 ;
        RECT 1203.000 2797.250 1203.260 2797.510 ;
        RECT 1201.545 2797.190 1203.260 2797.250 ;
        RECT 2901.320 2797.190 2901.580 2797.510 ;
        RECT 1201.545 2797.110 1203.200 2797.190 ;
        RECT 1201.545 2796.000 1201.825 2797.110 ;
        RECT 2901.380 381.325 2901.520 2797.190 ;
        RECT 2901.310 380.955 2901.590 381.325 ;
      LAYER via2 ;
        RECT 2901.310 381.000 2901.590 381.280 ;
      LAYER met3 ;
        RECT 2901.285 381.290 2901.615 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2901.285 380.990 2924.800 381.290 ;
        RECT 2901.285 380.975 2901.615 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3500.540 1095.190 3500.600 ;
        RECT 1745.770 3500.540 1746.090 3500.600 ;
        RECT 1094.870 3500.400 1746.090 3500.540 ;
        RECT 1094.870 3500.340 1095.190 3500.400 ;
        RECT 1745.770 3500.340 1746.090 3500.400 ;
      LAYER via ;
        RECT 1094.900 3500.340 1095.160 3500.600 ;
        RECT 1745.800 3500.340 1746.060 3500.600 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3500.630 1095.100 3517.600 ;
        RECT 1094.900 3500.310 1095.160 3500.630 ;
        RECT 1745.800 3500.310 1746.060 3500.630 ;
        RECT 1745.860 2801.330 1746.000 3500.310 ;
        RECT 1745.860 2801.190 1749.680 2801.330 ;
        RECT 1749.540 2799.970 1749.680 2801.190 ;
        RECT 1751.705 2799.970 1751.985 2800.000 ;
        RECT 1749.540 2799.830 1751.985 2799.970 ;
        RECT 1751.705 2796.000 1751.985 2799.830 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3504.280 770.890 3504.340 ;
        RECT 1780.270 3504.280 1780.590 3504.340 ;
        RECT 770.570 3504.140 1780.590 3504.280 ;
        RECT 770.570 3504.080 770.890 3504.140 ;
        RECT 1780.270 3504.080 1780.590 3504.140 ;
      LAYER via ;
        RECT 770.600 3504.080 770.860 3504.340 ;
        RECT 1780.300 3504.080 1780.560 3504.340 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3504.370 770.800 3517.600 ;
        RECT 770.600 3504.050 770.860 3504.370 ;
        RECT 1780.300 3504.050 1780.560 3504.370 ;
        RECT 1780.360 2799.970 1780.500 3504.050 ;
        RECT 1780.685 2799.970 1780.965 2800.000 ;
        RECT 1780.360 2799.830 1780.965 2799.970 ;
        RECT 1780.685 2796.000 1780.965 2799.830 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3502.580 446.130 3502.640 ;
        RECT 1807.870 3502.580 1808.190 3502.640 ;
        RECT 445.810 3502.440 1808.190 3502.580 ;
        RECT 445.810 3502.380 446.130 3502.440 ;
        RECT 1807.870 3502.380 1808.190 3502.440 ;
      LAYER via ;
        RECT 445.840 3502.380 446.100 3502.640 ;
        RECT 1807.900 3502.380 1808.160 3502.640 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3502.670 446.040 3517.600 ;
        RECT 445.840 3502.350 446.100 3502.670 ;
        RECT 1807.900 3502.350 1808.160 3502.670 ;
        RECT 1807.960 2799.970 1808.100 3502.350 ;
        RECT 1809.665 2799.970 1809.945 2800.000 ;
        RECT 1807.960 2799.830 1809.945 2799.970 ;
        RECT 1809.665 2796.000 1809.945 2799.830 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1835.470 3501.560 1835.790 3501.620 ;
        RECT 121.510 3501.420 1835.790 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1835.470 3501.360 1835.790 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1835.500 3501.360 1835.760 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1835.500 3501.330 1835.760 3501.650 ;
        RECT 1835.560 2800.650 1835.700 3501.330 ;
        RECT 1835.560 2800.510 1837.080 2800.650 ;
        RECT 1836.940 2799.970 1837.080 2800.510 ;
        RECT 1838.645 2799.970 1838.925 2800.000 ;
        RECT 1836.940 2799.830 1838.925 2799.970 ;
        RECT 1838.645 2796.000 1838.925 2799.830 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1863.070 3339.720 1863.390 3339.780 ;
        RECT 17.090 3339.580 1863.390 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1863.070 3339.520 1863.390 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1863.100 3339.520 1863.360 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1863.100 3339.490 1863.360 3339.810 ;
        RECT 1863.160 2800.650 1863.300 3339.490 ;
        RECT 1863.160 2800.510 1866.060 2800.650 ;
        RECT 1865.920 2799.970 1866.060 2800.510 ;
        RECT 1867.625 2799.970 1867.905 2800.000 ;
        RECT 1865.920 2799.830 1867.905 2799.970 ;
        RECT 1867.625 2796.000 1867.905 2799.830 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 1890.670 3050.040 1890.990 3050.100 ;
        RECT 17.090 3049.900 1890.990 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 1890.670 3049.840 1890.990 3049.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 1890.700 3049.840 1890.960 3050.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 1890.700 3049.810 1890.960 3050.130 ;
        RECT 1890.760 2800.650 1890.900 3049.810 ;
        RECT 1890.760 2800.510 1894.580 2800.650 ;
        RECT 1894.440 2799.970 1894.580 2800.510 ;
        RECT 1896.145 2799.970 1896.425 2800.000 ;
        RECT 1894.440 2799.830 1896.425 2799.970 ;
        RECT 1896.145 2796.000 1896.425 2799.830 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1173.145 2796.925 1173.315 2797.775 ;
      LAYER mcon ;
        RECT 1173.145 2797.605 1173.315 2797.775 ;
      LAYER met1 ;
        RECT 1173.085 2797.760 1173.375 2797.805 ;
        RECT 1173.085 2797.620 1197.220 2797.760 ;
        RECT 1173.085 2797.575 1173.375 2797.620 ;
        RECT 27.670 2797.080 27.990 2797.140 ;
        RECT 1173.085 2797.080 1173.375 2797.125 ;
        RECT 27.670 2796.940 1173.375 2797.080 ;
        RECT 1197.080 2797.080 1197.220 2797.620 ;
        RECT 1924.250 2797.080 1924.570 2797.140 ;
        RECT 1197.080 2796.940 1924.570 2797.080 ;
        RECT 27.670 2796.880 27.990 2796.940 ;
        RECT 1173.085 2796.895 1173.375 2796.940 ;
        RECT 1924.250 2796.880 1924.570 2796.940 ;
        RECT 13.870 2765.460 14.190 2765.520 ;
        RECT 27.670 2765.460 27.990 2765.520 ;
        RECT 13.870 2765.320 27.990 2765.460 ;
        RECT 13.870 2765.260 14.190 2765.320 ;
        RECT 27.670 2765.260 27.990 2765.320 ;
      LAYER via ;
        RECT 27.700 2796.880 27.960 2797.140 ;
        RECT 1924.280 2796.880 1924.540 2797.140 ;
        RECT 13.900 2765.260 14.160 2765.520 ;
        RECT 27.700 2765.260 27.960 2765.520 ;
      LAYER met2 ;
        RECT 1925.125 2797.250 1925.405 2800.000 ;
        RECT 1924.340 2797.170 1925.405 2797.250 ;
        RECT 27.700 2796.850 27.960 2797.170 ;
        RECT 1924.280 2797.110 1925.405 2797.170 ;
        RECT 1924.280 2796.850 1924.540 2797.110 ;
        RECT 27.760 2765.550 27.900 2796.850 ;
        RECT 1925.125 2796.000 1925.405 2797.110 ;
        RECT 13.900 2765.405 14.160 2765.550 ;
        RECT 13.890 2765.035 14.170 2765.405 ;
        RECT 27.700 2765.230 27.960 2765.550 ;
      LAYER via2 ;
        RECT 13.890 2765.080 14.170 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 13.865 2765.370 14.195 2765.385 ;
        RECT -4.800 2765.070 14.195 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 13.865 2765.055 14.195 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 33.190 2811.360 33.510 2811.420 ;
        RECT 1954.150 2811.360 1954.470 2811.420 ;
        RECT 33.190 2811.220 1954.470 2811.360 ;
        RECT 33.190 2811.160 33.510 2811.220 ;
        RECT 1954.150 2811.160 1954.470 2811.220 ;
        RECT 15.250 2477.820 15.570 2477.880 ;
        RECT 33.190 2477.820 33.510 2477.880 ;
        RECT 15.250 2477.680 33.510 2477.820 ;
        RECT 15.250 2477.620 15.570 2477.680 ;
        RECT 33.190 2477.620 33.510 2477.680 ;
      LAYER via ;
        RECT 33.220 2811.160 33.480 2811.420 ;
        RECT 1954.180 2811.160 1954.440 2811.420 ;
        RECT 15.280 2477.620 15.540 2477.880 ;
        RECT 33.220 2477.620 33.480 2477.880 ;
      LAYER met2 ;
        RECT 33.220 2811.130 33.480 2811.450 ;
        RECT 1954.180 2811.130 1954.440 2811.450 ;
        RECT 33.280 2477.910 33.420 2811.130 ;
        RECT 1954.240 2800.000 1954.380 2811.130 ;
        RECT 1954.105 2796.000 1954.385 2800.000 ;
        RECT 15.280 2477.765 15.540 2477.910 ;
        RECT 15.270 2477.395 15.550 2477.765 ;
        RECT 33.220 2477.590 33.480 2477.910 ;
      LAYER via2 ;
        RECT 15.270 2477.440 15.550 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 15.245 2477.730 15.575 2477.745 ;
        RECT -4.800 2477.430 15.575 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 15.245 2477.415 15.575 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 32.270 2810.340 32.590 2810.400 ;
        RECT 1983.130 2810.340 1983.450 2810.400 ;
        RECT 32.270 2810.200 1983.450 2810.340 ;
        RECT 32.270 2810.140 32.590 2810.200 ;
        RECT 1983.130 2810.140 1983.450 2810.200 ;
        RECT 15.710 2193.580 16.030 2193.640 ;
        RECT 32.270 2193.580 32.590 2193.640 ;
        RECT 15.710 2193.440 32.590 2193.580 ;
        RECT 15.710 2193.380 16.030 2193.440 ;
        RECT 32.270 2193.380 32.590 2193.440 ;
      LAYER via ;
        RECT 32.300 2810.140 32.560 2810.400 ;
        RECT 1983.160 2810.140 1983.420 2810.400 ;
        RECT 15.740 2193.380 16.000 2193.640 ;
        RECT 32.300 2193.380 32.560 2193.640 ;
      LAYER met2 ;
        RECT 32.300 2810.110 32.560 2810.430 ;
        RECT 1983.160 2810.110 1983.420 2810.430 ;
        RECT 32.360 2193.670 32.500 2810.110 ;
        RECT 1983.220 2800.000 1983.360 2810.110 ;
        RECT 1983.085 2796.000 1983.365 2800.000 ;
        RECT 15.740 2193.350 16.000 2193.670 ;
        RECT 32.300 2193.350 32.560 2193.670 ;
        RECT 15.800 2190.125 15.940 2193.350 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
      LAYER via2 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.800 2189.790 16.035 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.810 2809.320 32.130 2809.380 ;
        RECT 2012.110 2809.320 2012.430 2809.380 ;
        RECT 31.810 2809.180 2012.430 2809.320 ;
        RECT 31.810 2809.120 32.130 2809.180 ;
        RECT 2012.110 2809.120 2012.430 2809.180 ;
        RECT 15.710 1903.220 16.030 1903.280 ;
        RECT 31.810 1903.220 32.130 1903.280 ;
        RECT 15.710 1903.080 32.130 1903.220 ;
        RECT 15.710 1903.020 16.030 1903.080 ;
        RECT 31.810 1903.020 32.130 1903.080 ;
      LAYER via ;
        RECT 31.840 2809.120 32.100 2809.380 ;
        RECT 2012.140 2809.120 2012.400 2809.380 ;
        RECT 15.740 1903.020 16.000 1903.280 ;
        RECT 31.840 1903.020 32.100 1903.280 ;
      LAYER met2 ;
        RECT 31.840 2809.090 32.100 2809.410 ;
        RECT 2012.140 2809.090 2012.400 2809.410 ;
        RECT 31.900 1903.310 32.040 2809.090 ;
        RECT 2012.200 2800.000 2012.340 2809.090 ;
        RECT 2012.065 2796.000 2012.345 2800.000 ;
        RECT 15.740 1903.165 16.000 1903.310 ;
        RECT 15.730 1902.795 16.010 1903.165 ;
        RECT 31.840 1902.990 32.100 1903.310 ;
      LAYER via2 ;
        RECT 15.730 1902.840 16.010 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 15.705 1903.130 16.035 1903.145 ;
        RECT -4.800 1902.830 16.035 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 15.705 1902.815 16.035 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1861.305 2797.605 1861.935 2797.775 ;
      LAYER mcon ;
        RECT 1861.765 2797.605 1861.935 2797.775 ;
      LAYER met1 ;
        RECT 1232.410 2797.760 1232.730 2797.820 ;
        RECT 1861.245 2797.760 1861.535 2797.805 ;
        RECT 1232.410 2797.620 1861.535 2797.760 ;
        RECT 1232.410 2797.560 1232.730 2797.620 ;
        RECT 1861.245 2797.575 1861.535 2797.620 ;
        RECT 1861.705 2797.760 1861.995 2797.805 ;
        RECT 2902.210 2797.760 2902.530 2797.820 ;
        RECT 1861.705 2797.620 2902.530 2797.760 ;
        RECT 1861.705 2797.575 1861.995 2797.620 ;
        RECT 2902.210 2797.560 2902.530 2797.620 ;
      LAYER via ;
        RECT 1232.440 2797.560 1232.700 2797.820 ;
        RECT 2902.240 2797.560 2902.500 2797.820 ;
      LAYER met2 ;
        RECT 1230.525 2797.930 1230.805 2800.000 ;
        RECT 1230.525 2797.850 1232.640 2797.930 ;
        RECT 1230.525 2797.790 1232.700 2797.850 ;
        RECT 1230.525 2796.000 1230.805 2797.790 ;
        RECT 1232.440 2797.530 1232.700 2797.790 ;
        RECT 2902.240 2797.530 2902.500 2797.850 ;
        RECT 2902.300 615.925 2902.440 2797.530 ;
        RECT 2902.230 615.555 2902.510 615.925 ;
      LAYER via2 ;
        RECT 2902.230 615.600 2902.510 615.880 ;
      LAYER met3 ;
        RECT 2902.205 615.890 2902.535 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2902.205 615.590 2924.800 615.890 ;
        RECT 2902.205 615.575 2902.535 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2808.980 16.950 2809.040 ;
        RECT 2041.090 2808.980 2041.410 2809.040 ;
        RECT 16.630 2808.840 2041.410 2808.980 ;
        RECT 16.630 2808.780 16.950 2808.840 ;
        RECT 2041.090 2808.780 2041.410 2808.840 ;
      LAYER via ;
        RECT 16.660 2808.780 16.920 2809.040 ;
        RECT 2041.120 2808.780 2041.380 2809.040 ;
      LAYER met2 ;
        RECT 16.660 2808.750 16.920 2809.070 ;
        RECT 2041.120 2808.750 2041.380 2809.070 ;
        RECT 16.720 1615.525 16.860 2808.750 ;
        RECT 2041.180 2800.000 2041.320 2808.750 ;
        RECT 2041.045 2796.000 2041.325 2800.000 ;
        RECT 16.650 1615.155 16.930 1615.525 ;
      LAYER via2 ;
        RECT 16.650 1615.200 16.930 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.625 1615.490 16.955 1615.505 ;
        RECT -4.800 1615.190 16.955 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.625 1615.175 16.955 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.350 2808.640 31.670 2808.700 ;
        RECT 2070.070 2808.640 2070.390 2808.700 ;
        RECT 31.350 2808.500 2070.390 2808.640 ;
        RECT 31.350 2808.440 31.670 2808.500 ;
        RECT 2070.070 2808.440 2070.390 2808.500 ;
        RECT 15.710 1400.700 16.030 1400.760 ;
        RECT 31.350 1400.700 31.670 1400.760 ;
        RECT 15.710 1400.560 31.670 1400.700 ;
        RECT 15.710 1400.500 16.030 1400.560 ;
        RECT 31.350 1400.500 31.670 1400.560 ;
      LAYER via ;
        RECT 31.380 2808.440 31.640 2808.700 ;
        RECT 2070.100 2808.440 2070.360 2808.700 ;
        RECT 15.740 1400.500 16.000 1400.760 ;
        RECT 31.380 1400.500 31.640 1400.760 ;
      LAYER met2 ;
        RECT 31.380 2808.410 31.640 2808.730 ;
        RECT 2070.100 2808.410 2070.360 2808.730 ;
        RECT 31.440 1400.790 31.580 2808.410 ;
        RECT 2070.160 2800.000 2070.300 2808.410 ;
        RECT 2070.025 2796.000 2070.305 2800.000 ;
        RECT 15.740 1400.645 16.000 1400.790 ;
        RECT 15.730 1400.275 16.010 1400.645 ;
        RECT 31.380 1400.470 31.640 1400.790 ;
      LAYER via2 ;
        RECT 15.730 1400.320 16.010 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 15.705 1400.610 16.035 1400.625 ;
        RECT -4.800 1400.310 16.035 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 15.705 1400.295 16.035 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 2812.635 20.150 2813.005 ;
        RECT 19.940 1185.085 20.080 2812.635 ;
        RECT 2099.070 2811.275 2099.350 2811.645 ;
        RECT 2099.140 2800.000 2099.280 2811.275 ;
        RECT 2099.005 2796.000 2099.285 2800.000 ;
        RECT 19.870 1184.715 20.150 1185.085 ;
      LAYER via2 ;
        RECT 19.870 2812.680 20.150 2812.960 ;
        RECT 2099.070 2811.320 2099.350 2811.600 ;
        RECT 19.870 1184.760 20.150 1185.040 ;
      LAYER met3 ;
        RECT 19.845 2812.970 20.175 2812.985 ;
        RECT 19.845 2812.670 28.210 2812.970 ;
        RECT 19.845 2812.655 20.175 2812.670 ;
        RECT 27.910 2811.610 28.210 2812.670 ;
        RECT 2099.045 2811.610 2099.375 2811.625 ;
        RECT 27.910 2811.310 2099.375 2811.610 ;
        RECT 2099.045 2811.295 2099.375 2811.310 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 19.845 1185.050 20.175 1185.065 ;
        RECT -4.800 1184.750 20.175 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 19.845 1184.735 20.175 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 2811.275 19.230 2811.645 ;
        RECT 26.770 2811.275 27.050 2811.645 ;
        RECT 19.020 969.525 19.160 2811.275 ;
        RECT 26.840 2810.285 26.980 2811.275 ;
        RECT 26.770 2809.915 27.050 2810.285 ;
        RECT 2128.050 2809.915 2128.330 2810.285 ;
        RECT 2128.120 2800.000 2128.260 2809.915 ;
        RECT 2127.985 2796.000 2128.265 2800.000 ;
        RECT 18.950 969.155 19.230 969.525 ;
      LAYER via2 ;
        RECT 18.950 2811.320 19.230 2811.600 ;
        RECT 26.770 2811.320 27.050 2811.600 ;
        RECT 26.770 2809.960 27.050 2810.240 ;
        RECT 2128.050 2809.960 2128.330 2810.240 ;
        RECT 18.950 969.200 19.230 969.480 ;
      LAYER met3 ;
        RECT 18.925 2811.610 19.255 2811.625 ;
        RECT 26.745 2811.610 27.075 2811.625 ;
        RECT 18.925 2811.310 27.075 2811.610 ;
        RECT 18.925 2811.295 19.255 2811.310 ;
        RECT 26.745 2811.295 27.075 2811.310 ;
        RECT 26.745 2810.250 27.075 2810.265 ;
        RECT 2128.025 2810.250 2128.355 2810.265 ;
        RECT 26.745 2809.950 2128.355 2810.250 ;
        RECT 26.745 2809.935 27.075 2809.950 ;
        RECT 2128.025 2809.935 2128.355 2809.950 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 18.925 969.490 19.255 969.505 ;
        RECT -4.800 969.190 19.255 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 18.925 969.175 19.255 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1183.265 2796.415 1183.435 2796.755 ;
        RECT 1184.185 2796.415 1184.355 2797.095 ;
        RECT 1926.625 2796.755 1926.795 2797.095 ;
        RECT 2079.345 2796.755 2079.515 2797.095 ;
        RECT 1508.485 2796.585 1509.575 2796.755 ;
        RECT 1605.085 2796.585 1606.175 2796.755 ;
        RECT 1701.685 2796.585 1702.775 2796.755 ;
        RECT 1848.885 2796.585 1850.435 2796.755 ;
        RECT 1926.625 2796.585 1927.715 2796.755 ;
        RECT 2042.085 2796.585 2043.175 2796.755 ;
        RECT 2079.345 2796.585 2080.435 2796.755 ;
        RECT 1183.265 2796.245 1184.355 2796.415 ;
      LAYER mcon ;
        RECT 1184.185 2796.925 1184.355 2797.095 ;
        RECT 1183.265 2796.585 1183.435 2796.755 ;
        RECT 1926.625 2796.925 1926.795 2797.095 ;
        RECT 2079.345 2796.925 2079.515 2797.095 ;
        RECT 1509.405 2796.585 1509.575 2796.755 ;
        RECT 1606.005 2796.585 1606.175 2796.755 ;
        RECT 1702.605 2796.585 1702.775 2796.755 ;
        RECT 1850.265 2796.585 1850.435 2796.755 ;
        RECT 1927.545 2796.585 1927.715 2796.755 ;
        RECT 2043.005 2796.585 2043.175 2796.755 ;
        RECT 2080.265 2796.585 2080.435 2796.755 ;
      LAYER met1 ;
        RECT 1184.125 2797.080 1184.415 2797.125 ;
        RECT 1926.565 2797.080 1926.855 2797.125 ;
        RECT 1184.125 2796.940 1196.760 2797.080 ;
        RECT 1184.125 2796.895 1184.415 2796.940 ;
        RECT 18.470 2796.740 18.790 2796.800 ;
        RECT 1183.205 2796.740 1183.495 2796.785 ;
        RECT 18.470 2796.600 1183.495 2796.740 ;
        RECT 1196.620 2796.740 1196.760 2796.940 ;
        RECT 1924.800 2796.940 1926.855 2797.080 ;
        RECT 1508.425 2796.740 1508.715 2796.785 ;
        RECT 1196.620 2796.600 1508.715 2796.740 ;
        RECT 18.470 2796.540 18.790 2796.600 ;
        RECT 1183.205 2796.555 1183.495 2796.600 ;
        RECT 1508.425 2796.555 1508.715 2796.600 ;
        RECT 1509.345 2796.740 1509.635 2796.785 ;
        RECT 1605.025 2796.740 1605.315 2796.785 ;
        RECT 1509.345 2796.600 1605.315 2796.740 ;
        RECT 1509.345 2796.555 1509.635 2796.600 ;
        RECT 1605.025 2796.555 1605.315 2796.600 ;
        RECT 1605.945 2796.740 1606.235 2796.785 ;
        RECT 1701.625 2796.740 1701.915 2796.785 ;
        RECT 1605.945 2796.600 1701.915 2796.740 ;
        RECT 1605.945 2796.555 1606.235 2796.600 ;
        RECT 1701.625 2796.555 1701.915 2796.600 ;
        RECT 1702.545 2796.740 1702.835 2796.785 ;
        RECT 1848.825 2796.740 1849.115 2796.785 ;
        RECT 1702.545 2796.600 1849.115 2796.740 ;
        RECT 1702.545 2796.555 1702.835 2796.600 ;
        RECT 1848.825 2796.555 1849.115 2796.600 ;
        RECT 1850.205 2796.740 1850.495 2796.785 ;
        RECT 1924.800 2796.740 1924.940 2796.940 ;
        RECT 1926.565 2796.895 1926.855 2796.940 ;
        RECT 1981.750 2796.880 1982.070 2797.140 ;
        RECT 2079.285 2797.080 2079.575 2797.125 ;
        RECT 2078.440 2796.940 2079.575 2797.080 ;
        RECT 1850.205 2796.600 1924.940 2796.740 ;
        RECT 1927.485 2796.740 1927.775 2796.785 ;
        RECT 1980.370 2796.740 1980.690 2796.800 ;
        RECT 1927.485 2796.600 1980.690 2796.740 ;
        RECT 1981.840 2796.740 1981.980 2796.880 ;
        RECT 2042.025 2796.740 2042.315 2796.785 ;
        RECT 1981.840 2796.600 2042.315 2796.740 ;
        RECT 1850.205 2796.555 1850.495 2796.600 ;
        RECT 1927.485 2796.555 1927.775 2796.600 ;
        RECT 1980.370 2796.540 1980.690 2796.600 ;
        RECT 2042.025 2796.555 2042.315 2796.600 ;
        RECT 2042.945 2796.740 2043.235 2796.785 ;
        RECT 2078.440 2796.740 2078.580 2796.940 ;
        RECT 2079.285 2796.895 2079.575 2796.940 ;
        RECT 2042.945 2796.600 2078.580 2796.740 ;
        RECT 2080.205 2796.740 2080.495 2796.785 ;
        RECT 2155.630 2796.740 2155.950 2796.800 ;
        RECT 2080.205 2796.600 2155.950 2796.740 ;
        RECT 2042.945 2796.555 2043.235 2796.600 ;
        RECT 2080.205 2796.555 2080.495 2796.600 ;
        RECT 2155.630 2796.540 2155.950 2796.600 ;
      LAYER via ;
        RECT 18.500 2796.540 18.760 2796.800 ;
        RECT 1981.780 2796.880 1982.040 2797.140 ;
        RECT 1980.400 2796.540 1980.660 2796.800 ;
        RECT 2155.660 2796.540 2155.920 2796.800 ;
      LAYER met2 ;
        RECT 1980.460 2797.170 1981.980 2797.250 ;
        RECT 1980.460 2797.110 1982.040 2797.170 ;
        RECT 1980.460 2796.830 1980.600 2797.110 ;
        RECT 1981.780 2796.850 1982.040 2797.110 ;
        RECT 18.500 2796.510 18.760 2796.830 ;
        RECT 1980.400 2796.510 1980.660 2796.830 ;
        RECT 2155.660 2796.570 2155.920 2796.830 ;
        RECT 2156.965 2796.570 2157.245 2800.000 ;
        RECT 2155.660 2796.510 2157.245 2796.570 ;
        RECT 18.560 753.965 18.700 2796.510 ;
        RECT 2155.720 2796.430 2157.245 2796.510 ;
        RECT 2156.965 2796.000 2157.245 2796.430 ;
        RECT 18.490 753.595 18.770 753.965 ;
      LAYER via2 ;
        RECT 18.490 753.640 18.770 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 18.465 753.930 18.795 753.945 ;
        RECT -4.800 753.630 18.795 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 18.465 753.615 18.795 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.030 2808.555 18.310 2808.925 ;
        RECT 2186.010 2808.555 2186.290 2808.925 ;
        RECT 18.100 538.405 18.240 2808.555 ;
        RECT 2186.080 2800.000 2186.220 2808.555 ;
        RECT 2185.945 2796.000 2186.225 2800.000 ;
        RECT 18.030 538.035 18.310 538.405 ;
      LAYER via2 ;
        RECT 18.030 2808.600 18.310 2808.880 ;
        RECT 2186.010 2808.600 2186.290 2808.880 ;
        RECT 18.030 538.080 18.310 538.360 ;
      LAYER met3 ;
        RECT 18.005 2808.890 18.335 2808.905 ;
        RECT 2185.985 2808.890 2186.315 2808.905 ;
        RECT 18.005 2808.590 2186.315 2808.890 ;
        RECT 18.005 2808.575 18.335 2808.590 ;
        RECT 2185.985 2808.575 2186.315 2808.590 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 18.005 538.370 18.335 538.385 ;
        RECT -4.800 538.070 18.335 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 18.005 538.055 18.335 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2173.130 2796.995 2173.410 2797.365 ;
        RECT 2214.070 2797.250 2214.350 2797.365 ;
        RECT 2214.925 2797.250 2215.205 2800.000 ;
        RECT 2214.070 2797.110 2215.205 2797.250 ;
        RECT 2214.070 2796.995 2214.350 2797.110 ;
        RECT 2173.200 2796.685 2173.340 2796.995 ;
        RECT 2173.130 2796.315 2173.410 2796.685 ;
        RECT 2214.925 2796.000 2215.205 2797.110 ;
        RECT 17.110 2794.955 17.390 2795.325 ;
        RECT 17.180 322.845 17.320 2794.955 ;
        RECT 17.110 322.475 17.390 322.845 ;
      LAYER via2 ;
        RECT 2173.130 2797.040 2173.410 2797.320 ;
        RECT 2214.070 2797.040 2214.350 2797.320 ;
        RECT 2173.130 2796.360 2173.410 2796.640 ;
        RECT 17.110 2795.000 17.390 2795.280 ;
        RECT 17.110 322.520 17.390 322.800 ;
      LAYER met3 ;
        RECT 1110.710 2797.330 1111.090 2797.340 ;
        RECT 1920.310 2797.330 1920.690 2797.340 ;
        RECT 2045.430 2797.330 2045.810 2797.340 ;
        RECT 2173.105 2797.330 2173.435 2797.345 ;
        RECT 2214.045 2797.330 2214.375 2797.345 ;
        RECT 1110.710 2797.030 1182.810 2797.330 ;
        RECT 1110.710 2797.020 1111.090 2797.030 ;
        RECT 1110.710 2795.970 1111.090 2795.980 ;
        RECT 1076.710 2795.670 1111.090 2795.970 ;
        RECT 17.085 2795.290 17.415 2795.305 ;
        RECT 1076.710 2795.290 1077.010 2795.670 ;
        RECT 1110.710 2795.660 1111.090 2795.670 ;
        RECT 17.085 2794.990 1077.010 2795.290 ;
        RECT 1182.510 2795.290 1182.810 2797.030 ;
        RECT 1263.470 2797.030 1458.810 2797.330 ;
        RECT 1262.510 2795.970 1262.890 2795.980 ;
        RECT 1263.470 2795.970 1263.770 2797.030 ;
        RECT 1458.510 2796.650 1458.810 2797.030 ;
        RECT 1920.310 2797.030 1972.170 2797.330 ;
        RECT 1920.310 2797.020 1920.690 2797.030 ;
        RECT 1497.110 2796.650 1497.490 2796.660 ;
        RECT 1458.510 2796.350 1497.490 2796.650 ;
        RECT 1497.110 2796.340 1497.490 2796.350 ;
        RECT 1262.510 2795.670 1263.770 2795.970 ;
        RECT 1559.670 2795.970 1560.050 2795.980 ;
        RECT 1760.230 2795.970 1760.610 2795.980 ;
        RECT 1920.310 2795.970 1920.690 2795.980 ;
        RECT 1559.670 2795.670 1594.050 2795.970 ;
        RECT 1262.510 2795.660 1262.890 2795.670 ;
        RECT 1559.670 2795.660 1560.050 2795.670 ;
        RECT 1593.750 2795.300 1594.050 2795.670 ;
        RECT 1656.310 2795.670 1684.210 2795.970 ;
        RECT 1220.190 2795.290 1220.570 2795.300 ;
        RECT 1182.510 2794.990 1220.570 2795.290 ;
        RECT 17.085 2794.975 17.415 2794.990 ;
        RECT 1220.190 2794.980 1220.570 2794.990 ;
        RECT 1497.110 2795.290 1497.490 2795.300 ;
        RECT 1558.750 2795.290 1559.130 2795.300 ;
        RECT 1497.110 2794.990 1559.130 2795.290 ;
        RECT 1497.110 2794.980 1497.490 2794.990 ;
        RECT 1558.750 2794.980 1559.130 2794.990 ;
        RECT 1593.710 2794.980 1594.090 2795.300 ;
        RECT 1220.190 2793.930 1220.570 2793.940 ;
        RECT 1262.510 2793.930 1262.890 2793.940 ;
        RECT 1220.190 2793.630 1262.890 2793.930 ;
        RECT 1220.190 2793.620 1220.570 2793.630 ;
        RECT 1262.510 2793.620 1262.890 2793.630 ;
        RECT 1593.710 2793.930 1594.090 2793.940 ;
        RECT 1656.310 2793.930 1656.610 2795.670 ;
        RECT 1683.910 2795.290 1684.210 2795.670 ;
        RECT 1760.230 2795.670 1807.490 2795.970 ;
        RECT 1760.230 2795.660 1760.610 2795.670 ;
        RECT 1690.310 2795.290 1690.690 2795.300 ;
        RECT 1759.310 2795.290 1759.690 2795.300 ;
        RECT 1683.910 2794.990 1690.690 2795.290 ;
        RECT 1690.310 2794.980 1690.690 2794.990 ;
        RECT 1758.430 2794.990 1759.690 2795.290 ;
        RECT 1807.190 2795.290 1807.490 2795.670 ;
        RECT 1879.870 2795.670 1920.690 2795.970 ;
        RECT 1879.870 2795.290 1880.170 2795.670 ;
        RECT 1920.310 2795.660 1920.690 2795.670 ;
        RECT 1807.190 2794.990 1880.170 2795.290 ;
        RECT 1971.870 2795.290 1972.170 2797.030 ;
        RECT 2045.430 2797.030 2076.820 2797.330 ;
        RECT 2045.430 2797.020 2045.810 2797.030 ;
        RECT 1980.110 2796.650 1980.490 2796.660 ;
        RECT 1980.110 2796.350 2021.850 2796.650 ;
        RECT 1980.110 2796.340 1980.490 2796.350 ;
        RECT 1980.110 2795.290 1980.490 2795.300 ;
        RECT 1971.870 2794.990 1980.490 2795.290 ;
        RECT 2021.550 2795.290 2021.850 2796.350 ;
        RECT 2076.520 2795.970 2076.820 2797.030 ;
        RECT 2173.105 2797.030 2214.375 2797.330 ;
        RECT 2173.105 2797.015 2173.435 2797.030 ;
        RECT 2214.045 2797.015 2214.375 2797.030 ;
        RECT 2138.390 2796.650 2140.530 2796.820 ;
        RECT 2173.105 2796.650 2173.435 2796.665 ;
        RECT 2138.390 2796.520 2173.435 2796.650 ;
        RECT 2138.390 2795.970 2138.690 2796.520 ;
        RECT 2140.230 2796.350 2173.435 2796.520 ;
        RECT 2173.105 2796.335 2173.435 2796.350 ;
        RECT 2076.520 2795.670 2138.690 2795.970 ;
        RECT 2045.430 2795.290 2045.810 2795.300 ;
        RECT 2021.550 2794.990 2045.810 2795.290 ;
        RECT 1593.710 2793.630 1656.610 2793.930 ;
        RECT 1690.310 2793.930 1690.690 2793.940 ;
        RECT 1758.430 2793.930 1758.730 2794.990 ;
        RECT 1759.310 2794.980 1759.690 2794.990 ;
        RECT 1980.110 2794.980 1980.490 2794.990 ;
        RECT 2045.430 2794.980 2045.810 2794.990 ;
        RECT 1690.310 2793.630 1758.730 2793.930 ;
        RECT 1593.710 2793.620 1594.090 2793.630 ;
        RECT 1690.310 2793.620 1690.690 2793.630 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 17.085 322.810 17.415 322.825 ;
        RECT -4.800 322.510 17.415 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 17.085 322.495 17.415 322.510 ;
      LAYER via3 ;
        RECT 1110.740 2797.020 1111.060 2797.340 ;
        RECT 1110.740 2795.660 1111.060 2795.980 ;
        RECT 1262.540 2795.660 1262.860 2795.980 ;
        RECT 1920.340 2797.020 1920.660 2797.340 ;
        RECT 1497.140 2796.340 1497.460 2796.660 ;
        RECT 1559.700 2795.660 1560.020 2795.980 ;
        RECT 1220.220 2794.980 1220.540 2795.300 ;
        RECT 1497.140 2794.980 1497.460 2795.300 ;
        RECT 1558.780 2794.980 1559.100 2795.300 ;
        RECT 1593.740 2794.980 1594.060 2795.300 ;
        RECT 1220.220 2793.620 1220.540 2793.940 ;
        RECT 1262.540 2793.620 1262.860 2793.940 ;
        RECT 1593.740 2793.620 1594.060 2793.940 ;
        RECT 1760.260 2795.660 1760.580 2795.980 ;
        RECT 1690.340 2794.980 1690.660 2795.300 ;
        RECT 1690.340 2793.620 1690.660 2793.940 ;
        RECT 1759.340 2794.980 1759.660 2795.300 ;
        RECT 1920.340 2795.660 1920.660 2795.980 ;
        RECT 2045.460 2797.020 2045.780 2797.340 ;
        RECT 1980.140 2796.340 1980.460 2796.660 ;
        RECT 1980.140 2794.980 1980.460 2795.300 ;
        RECT 2045.460 2794.980 2045.780 2795.300 ;
      LAYER met4 ;
        RECT 1110.735 2797.015 1111.065 2797.345 ;
        RECT 1920.335 2797.015 1920.665 2797.345 ;
        RECT 2045.455 2797.015 2045.785 2797.345 ;
        RECT 1110.750 2795.985 1111.050 2797.015 ;
        RECT 1497.135 2796.335 1497.465 2796.665 ;
        RECT 1558.790 2796.350 1560.010 2796.650 ;
        RECT 1110.735 2795.655 1111.065 2795.985 ;
        RECT 1262.535 2795.655 1262.865 2795.985 ;
        RECT 1220.215 2794.975 1220.545 2795.305 ;
        RECT 1220.230 2793.945 1220.530 2794.975 ;
        RECT 1262.550 2793.945 1262.850 2795.655 ;
        RECT 1497.150 2795.305 1497.450 2796.335 ;
        RECT 1558.790 2795.305 1559.090 2796.350 ;
        RECT 1559.710 2795.985 1560.010 2796.350 ;
        RECT 1759.350 2796.350 1760.570 2796.650 ;
        RECT 1559.695 2795.655 1560.025 2795.985 ;
        RECT 1759.350 2795.305 1759.650 2796.350 ;
        RECT 1760.270 2795.985 1760.570 2796.350 ;
        RECT 1920.350 2795.985 1920.650 2797.015 ;
        RECT 1980.135 2796.335 1980.465 2796.665 ;
        RECT 1760.255 2795.655 1760.585 2795.985 ;
        RECT 1920.335 2795.655 1920.665 2795.985 ;
        RECT 1980.150 2795.305 1980.450 2796.335 ;
        RECT 2045.470 2795.305 2045.770 2797.015 ;
        RECT 1497.135 2794.975 1497.465 2795.305 ;
        RECT 1558.775 2794.975 1559.105 2795.305 ;
        RECT 1593.735 2794.975 1594.065 2795.305 ;
        RECT 1690.335 2794.975 1690.665 2795.305 ;
        RECT 1759.335 2794.975 1759.665 2795.305 ;
        RECT 1980.135 2794.975 1980.465 2795.305 ;
        RECT 2045.455 2794.975 2045.785 2795.305 ;
        RECT 1593.750 2793.945 1594.050 2794.975 ;
        RECT 1690.350 2793.945 1690.650 2794.975 ;
        RECT 1220.215 2793.615 1220.545 2793.945 ;
        RECT 1262.535 2793.615 1262.865 2793.945 ;
        RECT 1593.735 2793.615 1594.065 2793.945 ;
        RECT 1690.335 2793.615 1690.665 2793.945 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2242.590 2796.570 2242.870 2796.685 ;
        RECT 2243.905 2796.570 2244.185 2800.000 ;
        RECT 2242.590 2796.430 2244.185 2796.570 ;
        RECT 2242.590 2796.315 2242.870 2796.430 ;
        RECT 2243.905 2796.000 2244.185 2796.430 ;
      LAYER via2 ;
        RECT 2242.590 2796.360 2242.870 2796.640 ;
      LAYER met3 ;
        RECT 2242.565 2796.660 2242.895 2796.665 ;
        RECT 2242.310 2796.650 2242.895 2796.660 ;
        RECT 2242.110 2796.350 2242.895 2796.650 ;
        RECT 2242.310 2796.340 2242.895 2796.350 ;
        RECT 2242.565 2796.335 2242.895 2796.340 ;
        RECT 2242.310 109.970 2242.690 109.980 ;
        RECT 3.070 109.670 2242.690 109.970 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 3.070 107.250 3.370 109.670 ;
        RECT 2242.310 109.660 2242.690 109.670 ;
        RECT -4.800 106.950 3.370 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
      LAYER via3 ;
        RECT 2242.340 2796.340 2242.660 2796.660 ;
        RECT 2242.340 109.660 2242.660 109.980 ;
      LAYER met4 ;
        RECT 2242.335 2796.335 2242.665 2796.665 ;
        RECT 2242.350 109.985 2242.650 2796.335 ;
        RECT 2242.335 109.655 2242.665 109.985 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1952.845 2797.945 1953.935 2798.115 ;
      LAYER mcon ;
        RECT 1953.765 2797.945 1953.935 2798.115 ;
      LAYER met1 ;
        RECT 1260.930 2798.100 1261.250 2798.160 ;
        RECT 1952.785 2798.100 1953.075 2798.145 ;
        RECT 1260.930 2797.960 1953.075 2798.100 ;
        RECT 1260.930 2797.900 1261.250 2797.960 ;
        RECT 1952.785 2797.915 1953.075 2797.960 ;
        RECT 1953.705 2798.100 1953.995 2798.145 ;
        RECT 2903.130 2798.100 2903.450 2798.160 ;
        RECT 1953.705 2797.960 2903.450 2798.100 ;
        RECT 1953.705 2797.915 1953.995 2797.960 ;
        RECT 2903.130 2797.900 2903.450 2797.960 ;
      LAYER via ;
        RECT 1260.960 2797.900 1261.220 2798.160 ;
        RECT 2903.160 2797.900 2903.420 2798.160 ;
      LAYER met2 ;
        RECT 1259.505 2797.930 1259.785 2800.000 ;
        RECT 1260.960 2797.930 1261.220 2798.190 ;
        RECT 1259.505 2797.870 1261.220 2797.930 ;
        RECT 2903.160 2797.870 2903.420 2798.190 ;
        RECT 1259.505 2797.790 1261.160 2797.870 ;
        RECT 1259.505 2796.000 1259.785 2797.790 ;
        RECT 2903.220 850.525 2903.360 2797.870 ;
        RECT 2903.150 850.155 2903.430 850.525 ;
      LAYER via2 ;
        RECT 2903.150 850.200 2903.430 850.480 ;
      LAYER met3 ;
        RECT 2903.125 850.490 2903.455 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2903.125 850.190 2924.800 850.490 ;
        RECT 2903.125 850.175 2903.455 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1953.305 2798.285 1954.395 2798.455 ;
      LAYER mcon ;
        RECT 1954.225 2798.285 1954.395 2798.455 ;
      LAYER met1 ;
        RECT 1290.370 2798.440 1290.690 2798.500 ;
        RECT 1953.245 2798.440 1953.535 2798.485 ;
        RECT 1290.370 2798.300 1953.535 2798.440 ;
        RECT 1290.370 2798.240 1290.690 2798.300 ;
        RECT 1953.245 2798.255 1953.535 2798.300 ;
        RECT 1954.165 2798.440 1954.455 2798.485 ;
        RECT 2903.590 2798.440 2903.910 2798.500 ;
        RECT 1954.165 2798.300 2903.910 2798.440 ;
        RECT 1954.165 2798.255 1954.455 2798.300 ;
        RECT 2903.590 2798.240 2903.910 2798.300 ;
      LAYER via ;
        RECT 1290.400 2798.240 1290.660 2798.500 ;
        RECT 2903.620 2798.240 2903.880 2798.500 ;
      LAYER met2 ;
        RECT 1288.485 2798.610 1288.765 2800.000 ;
        RECT 1288.485 2798.530 1290.600 2798.610 ;
        RECT 1288.485 2798.470 1290.660 2798.530 ;
        RECT 1288.485 2796.000 1288.765 2798.470 ;
        RECT 1290.400 2798.210 1290.660 2798.470 ;
        RECT 2903.620 2798.210 2903.880 2798.530 ;
        RECT 2903.680 1085.125 2903.820 2798.210 ;
        RECT 2903.610 1084.755 2903.890 1085.125 ;
      LAYER via2 ;
        RECT 2903.610 1084.800 2903.890 1085.080 ;
      LAYER met3 ;
        RECT 2903.585 1085.090 2903.915 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2903.585 1084.790 2924.800 1085.090 ;
        RECT 2903.585 1084.775 2903.915 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1860.845 2798.965 1862.855 2799.135 ;
        RECT 1953.305 2798.965 1954.395 2799.135 ;
        RECT 2001.145 2798.965 2002.235 2799.135 ;
      LAYER mcon ;
        RECT 1862.685 2798.965 1862.855 2799.135 ;
        RECT 1954.225 2798.965 1954.395 2799.135 ;
        RECT 2002.065 2798.965 2002.235 2799.135 ;
      LAYER met1 ;
        RECT 1317.970 2799.120 1318.290 2799.180 ;
        RECT 1860.785 2799.120 1861.075 2799.165 ;
        RECT 1317.970 2798.980 1861.075 2799.120 ;
        RECT 1317.970 2798.920 1318.290 2798.980 ;
        RECT 1860.785 2798.935 1861.075 2798.980 ;
        RECT 1862.625 2799.120 1862.915 2799.165 ;
        RECT 1953.245 2799.120 1953.535 2799.165 ;
        RECT 1862.625 2798.980 1953.535 2799.120 ;
        RECT 1862.625 2798.935 1862.915 2798.980 ;
        RECT 1953.245 2798.935 1953.535 2798.980 ;
        RECT 1954.165 2799.120 1954.455 2799.165 ;
        RECT 2001.085 2799.120 2001.375 2799.165 ;
        RECT 1954.165 2798.980 2001.375 2799.120 ;
        RECT 1954.165 2798.935 1954.455 2798.980 ;
        RECT 2001.085 2798.935 2001.375 2798.980 ;
        RECT 2002.005 2799.120 2002.295 2799.165 ;
        RECT 2900.830 2799.120 2901.150 2799.180 ;
        RECT 2002.005 2798.980 2901.150 2799.120 ;
        RECT 2002.005 2798.935 2002.295 2798.980 ;
        RECT 2900.830 2798.920 2901.150 2798.980 ;
      LAYER via ;
        RECT 1318.000 2798.920 1318.260 2799.180 ;
        RECT 2900.860 2798.920 2901.120 2799.180 ;
      LAYER met2 ;
        RECT 1317.465 2799.290 1317.745 2800.000 ;
        RECT 1317.465 2799.210 1318.200 2799.290 ;
        RECT 1317.465 2799.150 1318.260 2799.210 ;
        RECT 1317.465 2796.000 1317.745 2799.150 ;
        RECT 1318.000 2798.890 1318.260 2799.150 ;
        RECT 2900.860 2798.890 2901.120 2799.210 ;
        RECT 2900.920 1319.725 2901.060 2798.890 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2001.605 2799.985 2002.695 2800.155 ;
      LAYER mcon ;
        RECT 2002.525 2799.985 2002.695 2800.155 ;
      LAYER met1 ;
        RECT 1348.330 2800.140 1348.650 2800.200 ;
        RECT 2001.545 2800.140 2001.835 2800.185 ;
        RECT 1348.330 2800.000 2001.835 2800.140 ;
        RECT 1348.330 2799.940 1348.650 2800.000 ;
        RECT 2001.545 2799.955 2001.835 2800.000 ;
        RECT 2002.465 2800.140 2002.755 2800.185 ;
        RECT 2899.910 2800.140 2900.230 2800.200 ;
        RECT 2002.465 2800.000 2900.230 2800.140 ;
        RECT 2002.465 2799.955 2002.755 2800.000 ;
        RECT 2899.910 2799.940 2900.230 2800.000 ;
      LAYER via ;
        RECT 1348.360 2799.940 1348.620 2800.200 ;
        RECT 2899.940 2799.940 2900.200 2800.200 ;
      LAYER met2 ;
        RECT 1346.445 2799.970 1346.725 2800.000 ;
        RECT 1348.360 2799.970 1348.620 2800.230 ;
        RECT 1346.445 2799.910 1348.620 2799.970 ;
        RECT 2899.940 2799.910 2900.200 2800.230 ;
        RECT 1346.445 2799.830 1348.560 2799.910 ;
        RECT 1346.445 2796.000 1346.725 2799.830 ;
        RECT 2900.000 1554.325 2900.140 2799.910 ;
        RECT 2899.930 1553.955 2900.210 1554.325 ;
      LAYER via2 ;
        RECT 2899.930 1554.000 2900.210 1554.280 ;
      LAYER met3 ;
        RECT 2899.905 1554.290 2900.235 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2899.905 1553.990 2924.800 1554.290 ;
        RECT 2899.905 1553.975 2900.235 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1375.470 2800.480 1375.790 2800.540 ;
        RECT 2001.070 2800.480 2001.390 2800.540 ;
        RECT 1375.470 2800.340 2001.390 2800.480 ;
        RECT 1375.470 2800.280 1375.790 2800.340 ;
        RECT 2001.070 2800.280 2001.390 2800.340 ;
        RECT 2002.910 2800.480 2003.230 2800.540 ;
        RECT 2899.450 2800.480 2899.770 2800.540 ;
        RECT 2002.910 2800.340 2899.770 2800.480 ;
        RECT 2002.910 2800.280 2003.230 2800.340 ;
        RECT 2899.450 2800.280 2899.770 2800.340 ;
      LAYER via ;
        RECT 1375.500 2800.280 1375.760 2800.540 ;
        RECT 2001.100 2800.280 2001.360 2800.540 ;
        RECT 2002.940 2800.280 2003.200 2800.540 ;
        RECT 2899.480 2800.280 2899.740 2800.540 ;
      LAYER met2 ;
        RECT 1375.500 2800.250 1375.760 2800.570 ;
        RECT 2001.090 2800.395 2001.370 2800.765 ;
        RECT 2002.930 2800.395 2003.210 2800.765 ;
        RECT 2001.100 2800.250 2001.360 2800.395 ;
        RECT 2002.940 2800.250 2003.200 2800.395 ;
        RECT 2899.480 2800.250 2899.740 2800.570 ;
        RECT 1375.560 2800.000 1375.700 2800.250 ;
        RECT 1375.425 2796.000 1375.705 2800.000 ;
        RECT 2899.540 1789.605 2899.680 2800.250 ;
        RECT 2899.470 1789.235 2899.750 1789.605 ;
      LAYER via2 ;
        RECT 2001.090 2800.440 2001.370 2800.720 ;
        RECT 2002.930 2800.440 2003.210 2800.720 ;
        RECT 2899.470 1789.280 2899.750 1789.560 ;
      LAYER met3 ;
        RECT 2001.065 2800.730 2001.395 2800.745 ;
        RECT 2002.905 2800.730 2003.235 2800.745 ;
        RECT 2001.065 2800.430 2003.235 2800.730 ;
        RECT 2001.065 2800.415 2001.395 2800.430 ;
        RECT 2002.905 2800.415 2003.235 2800.430 ;
        RECT 2899.445 1789.570 2899.775 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2899.445 1789.270 2924.800 1789.570 ;
        RECT 2899.445 1789.255 2899.775 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1404.450 2813.740 1404.770 2813.800 ;
        RECT 2253.610 2813.740 2253.930 2813.800 ;
        RECT 1404.450 2813.600 2253.930 2813.740 ;
        RECT 1404.450 2813.540 1404.770 2813.600 ;
        RECT 2253.610 2813.540 2253.930 2813.600 ;
        RECT 2253.610 2028.340 2253.930 2028.400 ;
        RECT 2898.990 2028.340 2899.310 2028.400 ;
        RECT 2253.610 2028.200 2899.310 2028.340 ;
        RECT 2253.610 2028.140 2253.930 2028.200 ;
        RECT 2898.990 2028.140 2899.310 2028.200 ;
      LAYER via ;
        RECT 1404.480 2813.540 1404.740 2813.800 ;
        RECT 2253.640 2813.540 2253.900 2813.800 ;
        RECT 2253.640 2028.140 2253.900 2028.400 ;
        RECT 2899.020 2028.140 2899.280 2028.400 ;
      LAYER met2 ;
        RECT 1404.480 2813.510 1404.740 2813.830 ;
        RECT 2253.640 2813.510 2253.900 2813.830 ;
        RECT 1404.540 2800.000 1404.680 2813.510 ;
        RECT 1404.405 2796.000 1404.685 2800.000 ;
        RECT 2253.700 2028.430 2253.840 2813.510 ;
        RECT 2253.640 2028.110 2253.900 2028.430 ;
        RECT 2899.020 2028.110 2899.280 2028.430 ;
        RECT 2899.080 2024.205 2899.220 2028.110 ;
        RECT 2899.010 2023.835 2899.290 2024.205 ;
      LAYER via2 ;
        RECT 2899.010 2023.880 2899.290 2024.160 ;
      LAYER met3 ;
        RECT 2898.985 2024.170 2899.315 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2898.985 2023.870 2924.800 2024.170 ;
        RECT 2898.985 2023.855 2899.315 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1433.430 2813.060 1433.750 2813.120 ;
        RECT 2314.790 2813.060 2315.110 2813.120 ;
        RECT 1433.430 2812.920 2315.110 2813.060 ;
        RECT 1433.430 2812.860 1433.750 2812.920 ;
        RECT 2314.790 2812.860 2315.110 2812.920 ;
        RECT 2314.790 2262.940 2315.110 2263.000 ;
        RECT 2898.990 2262.940 2899.310 2263.000 ;
        RECT 2314.790 2262.800 2899.310 2262.940 ;
        RECT 2314.790 2262.740 2315.110 2262.800 ;
        RECT 2898.990 2262.740 2899.310 2262.800 ;
      LAYER via ;
        RECT 1433.460 2812.860 1433.720 2813.120 ;
        RECT 2314.820 2812.860 2315.080 2813.120 ;
        RECT 2314.820 2262.740 2315.080 2263.000 ;
        RECT 2899.020 2262.740 2899.280 2263.000 ;
      LAYER met2 ;
        RECT 1433.460 2812.830 1433.720 2813.150 ;
        RECT 2314.820 2812.830 2315.080 2813.150 ;
        RECT 1433.520 2800.000 1433.660 2812.830 ;
        RECT 1433.385 2796.000 1433.665 2800.000 ;
        RECT 2314.880 2263.030 2315.020 2812.830 ;
        RECT 2314.820 2262.710 2315.080 2263.030 ;
        RECT 2899.020 2262.710 2899.280 2263.030 ;
        RECT 2899.080 2258.805 2899.220 2262.710 ;
        RECT 2899.010 2258.435 2899.290 2258.805 ;
      LAYER via2 ;
        RECT 2899.010 2258.480 2899.290 2258.760 ;
      LAYER met3 ;
        RECT 2898.985 2258.770 2899.315 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2898.985 2258.470 2924.800 2258.770 ;
        RECT 2898.985 2258.455 2899.315 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 634.410 59.060 634.730 59.120 ;
        RECT 1387.890 59.060 1388.210 59.120 ;
        RECT 634.410 58.920 1388.210 59.060 ;
        RECT 634.410 58.860 634.730 58.920 ;
        RECT 1387.890 58.860 1388.210 58.920 ;
      LAYER via ;
        RECT 634.440 58.860 634.700 59.120 ;
        RECT 1387.920 58.860 1388.180 59.120 ;
      LAYER met2 ;
        RECT 1387.845 1700.000 1388.125 1704.000 ;
        RECT 1387.980 59.150 1388.120 1700.000 ;
        RECT 634.440 58.830 634.700 59.150 ;
        RECT 1387.920 58.830 1388.180 59.150 ;
        RECT 634.500 17.410 634.640 58.830 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 35.940 2063.030 36.000 ;
        RECT 2417.370 35.940 2417.690 36.000 ;
        RECT 2062.710 35.800 2417.690 35.940 ;
        RECT 2062.710 35.740 2063.030 35.800 ;
        RECT 2417.370 35.740 2417.690 35.800 ;
      LAYER via ;
        RECT 2062.740 35.740 2063.000 36.000 ;
        RECT 2417.400 35.740 2417.660 36.000 ;
      LAYER met2 ;
        RECT 2061.285 1700.410 2061.565 1704.000 ;
        RECT 2061.285 1700.270 2062.940 1700.410 ;
        RECT 2061.285 1700.000 2061.565 1700.270 ;
        RECT 2062.800 36.030 2062.940 1700.270 ;
        RECT 2062.740 35.710 2063.000 36.030 ;
        RECT 2417.400 35.710 2417.660 36.030 ;
        RECT 2417.460 2.400 2417.600 35.710 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2069.150 36.280 2069.470 36.340 ;
        RECT 2434.850 36.280 2435.170 36.340 ;
        RECT 2069.150 36.140 2435.170 36.280 ;
        RECT 2069.150 36.080 2069.470 36.140 ;
        RECT 2434.850 36.080 2435.170 36.140 ;
      LAYER via ;
        RECT 2069.180 36.080 2069.440 36.340 ;
        RECT 2434.880 36.080 2435.140 36.340 ;
      LAYER met2 ;
        RECT 2067.725 1700.410 2068.005 1704.000 ;
        RECT 2067.725 1700.270 2069.380 1700.410 ;
        RECT 2067.725 1700.000 2068.005 1700.270 ;
        RECT 2069.240 36.370 2069.380 1700.270 ;
        RECT 2069.180 36.050 2069.440 36.370 ;
        RECT 2434.880 36.050 2435.140 36.370 ;
        RECT 2434.940 2.400 2435.080 36.050 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2076.050 36.620 2076.370 36.680 ;
        RECT 2452.790 36.620 2453.110 36.680 ;
        RECT 2076.050 36.480 2453.110 36.620 ;
        RECT 2076.050 36.420 2076.370 36.480 ;
        RECT 2452.790 36.420 2453.110 36.480 ;
      LAYER via ;
        RECT 2076.080 36.420 2076.340 36.680 ;
        RECT 2452.820 36.420 2453.080 36.680 ;
      LAYER met2 ;
        RECT 2074.625 1700.410 2074.905 1704.000 ;
        RECT 2074.625 1700.270 2076.280 1700.410 ;
        RECT 2074.625 1700.000 2074.905 1700.270 ;
        RECT 2076.140 36.710 2076.280 1700.270 ;
        RECT 2076.080 36.390 2076.340 36.710 ;
        RECT 2452.820 36.390 2453.080 36.710 ;
        RECT 2452.880 2.400 2453.020 36.390 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2082.490 36.960 2082.810 37.020 ;
        RECT 2470.730 36.960 2471.050 37.020 ;
        RECT 2082.490 36.820 2471.050 36.960 ;
        RECT 2082.490 36.760 2082.810 36.820 ;
        RECT 2470.730 36.760 2471.050 36.820 ;
      LAYER via ;
        RECT 2082.520 36.760 2082.780 37.020 ;
        RECT 2470.760 36.760 2471.020 37.020 ;
      LAYER met2 ;
        RECT 2081.525 1700.410 2081.805 1704.000 ;
        RECT 2081.525 1700.270 2082.720 1700.410 ;
        RECT 2081.525 1700.000 2081.805 1700.270 ;
        RECT 2082.580 37.050 2082.720 1700.270 ;
        RECT 2082.520 36.730 2082.780 37.050 ;
        RECT 2470.760 36.730 2471.020 37.050 ;
        RECT 2470.820 2.400 2470.960 36.730 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2089.850 37.300 2090.170 37.360 ;
        RECT 2488.670 37.300 2488.990 37.360 ;
        RECT 2089.850 37.160 2488.990 37.300 ;
        RECT 2089.850 37.100 2090.170 37.160 ;
        RECT 2488.670 37.100 2488.990 37.160 ;
      LAYER via ;
        RECT 2089.880 37.100 2090.140 37.360 ;
        RECT 2488.700 37.100 2488.960 37.360 ;
      LAYER met2 ;
        RECT 2087.965 1700.410 2088.245 1704.000 ;
        RECT 2087.965 1700.270 2090.080 1700.410 ;
        RECT 2087.965 1700.000 2088.245 1700.270 ;
        RECT 2089.940 37.390 2090.080 1700.270 ;
        RECT 2089.880 37.070 2090.140 37.390 ;
        RECT 2488.700 37.070 2488.960 37.390 ;
        RECT 2488.760 2.400 2488.900 37.070 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2096.750 37.640 2097.070 37.700 ;
        RECT 2506.150 37.640 2506.470 37.700 ;
        RECT 2096.750 37.500 2506.470 37.640 ;
        RECT 2096.750 37.440 2097.070 37.500 ;
        RECT 2506.150 37.440 2506.470 37.500 ;
      LAYER via ;
        RECT 2096.780 37.440 2097.040 37.700 ;
        RECT 2506.180 37.440 2506.440 37.700 ;
      LAYER met2 ;
        RECT 2094.865 1700.410 2095.145 1704.000 ;
        RECT 2094.865 1700.270 2096.980 1700.410 ;
        RECT 2094.865 1700.000 2095.145 1700.270 ;
        RECT 2096.840 37.730 2096.980 1700.270 ;
        RECT 2096.780 37.410 2097.040 37.730 ;
        RECT 2506.180 37.410 2506.440 37.730 ;
        RECT 2506.240 2.400 2506.380 37.410 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2103.650 41.380 2103.970 41.440 ;
        RECT 2524.090 41.380 2524.410 41.440 ;
        RECT 2103.650 41.240 2524.410 41.380 ;
        RECT 2103.650 41.180 2103.970 41.240 ;
        RECT 2524.090 41.180 2524.410 41.240 ;
      LAYER via ;
        RECT 2103.680 41.180 2103.940 41.440 ;
        RECT 2524.120 41.180 2524.380 41.440 ;
      LAYER met2 ;
        RECT 2101.305 1701.090 2101.585 1704.000 ;
        RECT 2101.305 1700.950 2103.420 1701.090 ;
        RECT 2101.305 1700.000 2101.585 1700.950 ;
        RECT 2103.280 1688.850 2103.420 1700.950 ;
        RECT 2103.280 1688.710 2103.880 1688.850 ;
        RECT 2103.740 41.470 2103.880 1688.710 ;
        RECT 2103.680 41.150 2103.940 41.470 ;
        RECT 2524.120 41.150 2524.380 41.470 ;
        RECT 2524.180 2.400 2524.320 41.150 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2110.550 41.040 2110.870 41.100 ;
        RECT 2542.030 41.040 2542.350 41.100 ;
        RECT 2110.550 40.900 2542.350 41.040 ;
        RECT 2110.550 40.840 2110.870 40.900 ;
        RECT 2542.030 40.840 2542.350 40.900 ;
      LAYER via ;
        RECT 2110.580 40.840 2110.840 41.100 ;
        RECT 2542.060 40.840 2542.320 41.100 ;
      LAYER met2 ;
        RECT 2108.205 1700.410 2108.485 1704.000 ;
        RECT 2108.205 1700.270 2109.860 1700.410 ;
        RECT 2108.205 1700.000 2108.485 1700.270 ;
        RECT 2109.720 1688.850 2109.860 1700.270 ;
        RECT 2109.720 1688.710 2110.780 1688.850 ;
        RECT 2110.640 41.130 2110.780 1688.710 ;
        RECT 2110.580 40.810 2110.840 41.130 ;
        RECT 2542.060 40.810 2542.320 41.130 ;
        RECT 2542.120 2.400 2542.260 40.810 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2115.150 1688.680 2115.470 1688.740 ;
        RECT 2117.910 1688.680 2118.230 1688.740 ;
        RECT 2115.150 1688.540 2118.230 1688.680 ;
        RECT 2115.150 1688.480 2115.470 1688.540 ;
        RECT 2117.910 1688.480 2118.230 1688.540 ;
        RECT 2117.910 21.320 2118.230 21.380 ;
        RECT 2559.970 21.320 2560.290 21.380 ;
        RECT 2117.910 21.180 2560.290 21.320 ;
        RECT 2117.910 21.120 2118.230 21.180 ;
        RECT 2559.970 21.120 2560.290 21.180 ;
      LAYER via ;
        RECT 2115.180 1688.480 2115.440 1688.740 ;
        RECT 2117.940 1688.480 2118.200 1688.740 ;
        RECT 2117.940 21.120 2118.200 21.380 ;
        RECT 2560.000 21.120 2560.260 21.380 ;
      LAYER met2 ;
        RECT 2115.105 1700.000 2115.385 1704.000 ;
        RECT 2115.240 1688.770 2115.380 1700.000 ;
        RECT 2115.180 1688.450 2115.440 1688.770 ;
        RECT 2117.940 1688.450 2118.200 1688.770 ;
        RECT 2118.000 21.410 2118.140 1688.450 ;
        RECT 2117.940 21.090 2118.200 21.410 ;
        RECT 2560.000 21.090 2560.260 21.410 ;
        RECT 2560.060 2.400 2560.200 21.090 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2121.590 1688.680 2121.910 1688.740 ;
        RECT 2124.810 1688.680 2125.130 1688.740 ;
        RECT 2121.590 1688.540 2125.130 1688.680 ;
        RECT 2121.590 1688.480 2121.910 1688.540 ;
        RECT 2124.810 1688.480 2125.130 1688.540 ;
        RECT 2124.810 21.660 2125.130 21.720 ;
        RECT 2577.910 21.660 2578.230 21.720 ;
        RECT 2124.810 21.520 2578.230 21.660 ;
        RECT 2124.810 21.460 2125.130 21.520 ;
        RECT 2577.910 21.460 2578.230 21.520 ;
      LAYER via ;
        RECT 2121.620 1688.480 2121.880 1688.740 ;
        RECT 2124.840 1688.480 2125.100 1688.740 ;
        RECT 2124.840 21.460 2125.100 21.720 ;
        RECT 2577.940 21.460 2578.200 21.720 ;
      LAYER met2 ;
        RECT 2121.545 1700.000 2121.825 1704.000 ;
        RECT 2121.680 1688.770 2121.820 1700.000 ;
        RECT 2121.620 1688.450 2121.880 1688.770 ;
        RECT 2124.840 1688.450 2125.100 1688.770 ;
        RECT 2124.900 21.750 2125.040 1688.450 ;
        RECT 2124.840 21.430 2125.100 21.750 ;
        RECT 2577.940 21.430 2578.200 21.750 ;
        RECT 2578.000 2.400 2578.140 21.430 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1450.525 1538.925 1450.695 1579.555 ;
        RECT 1450.525 1364.845 1450.695 1400.715 ;
        RECT 1450.525 1264.205 1450.695 1304.155 ;
        RECT 1450.065 227.885 1450.235 275.655 ;
        RECT 1450.065 131.325 1450.235 179.435 ;
        RECT 1450.525 60.945 1450.695 62.475 ;
      LAYER mcon ;
        RECT 1450.525 1579.385 1450.695 1579.555 ;
        RECT 1450.525 1400.545 1450.695 1400.715 ;
        RECT 1450.525 1303.985 1450.695 1304.155 ;
        RECT 1450.065 275.485 1450.235 275.655 ;
        RECT 1450.065 179.265 1450.235 179.435 ;
        RECT 1450.525 62.305 1450.695 62.475 ;
      LAYER met1 ;
        RECT 1449.990 1642.440 1450.310 1642.500 ;
        RECT 1453.210 1642.440 1453.530 1642.500 ;
        RECT 1449.990 1642.300 1453.530 1642.440 ;
        RECT 1449.990 1642.240 1450.310 1642.300 ;
        RECT 1453.210 1642.240 1453.530 1642.300 ;
        RECT 1449.990 1607.900 1450.310 1608.160 ;
        RECT 1450.080 1607.420 1450.220 1607.900 ;
        RECT 1450.450 1607.420 1450.770 1607.480 ;
        RECT 1450.080 1607.280 1450.770 1607.420 ;
        RECT 1450.450 1607.220 1450.770 1607.280 ;
        RECT 1450.450 1579.540 1450.770 1579.600 ;
        RECT 1450.255 1579.400 1450.770 1579.540 ;
        RECT 1450.450 1579.340 1450.770 1579.400 ;
        RECT 1450.465 1539.080 1450.755 1539.125 ;
        RECT 1451.370 1539.080 1451.690 1539.140 ;
        RECT 1450.465 1538.940 1451.690 1539.080 ;
        RECT 1450.465 1538.895 1450.755 1538.940 ;
        RECT 1451.370 1538.880 1451.690 1538.940 ;
        RECT 1450.450 1497.600 1450.770 1497.660 ;
        RECT 1451.370 1497.600 1451.690 1497.660 ;
        RECT 1450.450 1497.460 1451.690 1497.600 ;
        RECT 1450.450 1497.400 1450.770 1497.460 ;
        RECT 1451.370 1497.400 1451.690 1497.460 ;
        RECT 1450.450 1400.700 1450.770 1400.760 ;
        RECT 1450.255 1400.560 1450.770 1400.700 ;
        RECT 1450.450 1400.500 1450.770 1400.560 ;
        RECT 1450.450 1365.000 1450.770 1365.060 ;
        RECT 1450.255 1364.860 1450.770 1365.000 ;
        RECT 1450.450 1364.800 1450.770 1364.860 ;
        RECT 1450.450 1304.140 1450.770 1304.200 ;
        RECT 1450.255 1304.000 1450.770 1304.140 ;
        RECT 1450.450 1303.940 1450.770 1304.000 ;
        RECT 1450.450 1264.360 1450.770 1264.420 ;
        RECT 1450.255 1264.220 1450.770 1264.360 ;
        RECT 1450.450 1264.160 1450.770 1264.220 ;
        RECT 1450.450 772.720 1450.770 772.780 ;
        RECT 1450.910 772.720 1451.230 772.780 ;
        RECT 1450.450 772.580 1451.230 772.720 ;
        RECT 1450.450 772.520 1450.770 772.580 ;
        RECT 1450.910 772.520 1451.230 772.580 ;
        RECT 1450.450 497.120 1450.770 497.380 ;
        RECT 1450.540 496.700 1450.680 497.120 ;
        RECT 1450.450 496.440 1450.770 496.700 ;
        RECT 1450.450 379.480 1450.770 379.740 ;
        RECT 1450.540 379.000 1450.680 379.480 ;
        RECT 1450.910 379.000 1451.230 379.060 ;
        RECT 1450.540 378.860 1451.230 379.000 ;
        RECT 1450.910 378.800 1451.230 378.860 ;
        RECT 1449.990 354.520 1450.310 354.580 ;
        RECT 1450.910 354.520 1451.230 354.580 ;
        RECT 1449.990 354.380 1451.230 354.520 ;
        RECT 1449.990 354.320 1450.310 354.380 ;
        RECT 1450.910 354.320 1451.230 354.380 ;
        RECT 1450.450 276.660 1450.770 276.720 ;
        RECT 1450.080 276.520 1450.770 276.660 ;
        RECT 1450.080 276.380 1450.220 276.520 ;
        RECT 1450.450 276.460 1450.770 276.520 ;
        RECT 1449.990 276.120 1450.310 276.380 ;
        RECT 1449.990 275.640 1450.310 275.700 ;
        RECT 1449.795 275.500 1450.310 275.640 ;
        RECT 1449.990 275.440 1450.310 275.500 ;
        RECT 1449.990 228.040 1450.310 228.100 ;
        RECT 1449.795 227.900 1450.310 228.040 ;
        RECT 1449.990 227.840 1450.310 227.900 ;
        RECT 1449.990 179.420 1450.310 179.480 ;
        RECT 1449.795 179.280 1450.310 179.420 ;
        RECT 1449.990 179.220 1450.310 179.280 ;
        RECT 1450.005 131.480 1450.295 131.525 ;
        RECT 1450.910 131.480 1451.230 131.540 ;
        RECT 1450.005 131.340 1451.230 131.480 ;
        RECT 1450.005 131.295 1450.295 131.340 ;
        RECT 1450.910 131.280 1451.230 131.340 ;
        RECT 1450.450 62.460 1450.770 62.520 ;
        RECT 1450.255 62.320 1450.770 62.460 ;
        RECT 1450.450 62.260 1450.770 62.320 ;
        RECT 811.510 61.100 811.830 61.160 ;
        RECT 1450.465 61.100 1450.755 61.145 ;
        RECT 811.510 60.960 1450.755 61.100 ;
        RECT 811.510 60.900 811.830 60.960 ;
        RECT 1450.465 60.915 1450.755 60.960 ;
      LAYER via ;
        RECT 1450.020 1642.240 1450.280 1642.500 ;
        RECT 1453.240 1642.240 1453.500 1642.500 ;
        RECT 1450.020 1607.900 1450.280 1608.160 ;
        RECT 1450.480 1607.220 1450.740 1607.480 ;
        RECT 1450.480 1579.340 1450.740 1579.600 ;
        RECT 1451.400 1538.880 1451.660 1539.140 ;
        RECT 1450.480 1497.400 1450.740 1497.660 ;
        RECT 1451.400 1497.400 1451.660 1497.660 ;
        RECT 1450.480 1400.500 1450.740 1400.760 ;
        RECT 1450.480 1364.800 1450.740 1365.060 ;
        RECT 1450.480 1303.940 1450.740 1304.200 ;
        RECT 1450.480 1264.160 1450.740 1264.420 ;
        RECT 1450.480 772.520 1450.740 772.780 ;
        RECT 1450.940 772.520 1451.200 772.780 ;
        RECT 1450.480 497.120 1450.740 497.380 ;
        RECT 1450.480 496.440 1450.740 496.700 ;
        RECT 1450.480 379.480 1450.740 379.740 ;
        RECT 1450.940 378.800 1451.200 379.060 ;
        RECT 1450.020 354.320 1450.280 354.580 ;
        RECT 1450.940 354.320 1451.200 354.580 ;
        RECT 1450.480 276.460 1450.740 276.720 ;
        RECT 1450.020 276.120 1450.280 276.380 ;
        RECT 1450.020 275.440 1450.280 275.700 ;
        RECT 1450.020 227.840 1450.280 228.100 ;
        RECT 1450.020 179.220 1450.280 179.480 ;
        RECT 1450.940 131.280 1451.200 131.540 ;
        RECT 1450.480 62.260 1450.740 62.520 ;
        RECT 811.540 60.900 811.800 61.160 ;
      LAYER met2 ;
        RECT 1455.005 1700.410 1455.285 1704.000 ;
        RECT 1453.300 1700.270 1455.285 1700.410 ;
        RECT 1453.300 1642.530 1453.440 1700.270 ;
        RECT 1455.005 1700.000 1455.285 1700.270 ;
        RECT 1450.020 1642.210 1450.280 1642.530 ;
        RECT 1453.240 1642.210 1453.500 1642.530 ;
        RECT 1450.080 1608.190 1450.220 1642.210 ;
        RECT 1450.020 1607.870 1450.280 1608.190 ;
        RECT 1450.480 1607.190 1450.740 1607.510 ;
        RECT 1450.540 1579.630 1450.680 1607.190 ;
        RECT 1450.480 1579.310 1450.740 1579.630 ;
        RECT 1451.400 1538.850 1451.660 1539.170 ;
        RECT 1451.460 1497.690 1451.600 1538.850 ;
        RECT 1450.480 1497.370 1450.740 1497.690 ;
        RECT 1451.400 1497.370 1451.660 1497.690 ;
        RECT 1450.540 1462.410 1450.680 1497.370 ;
        RECT 1450.080 1462.270 1450.680 1462.410 ;
        RECT 1450.080 1461.050 1450.220 1462.270 ;
        RECT 1450.080 1460.910 1450.680 1461.050 ;
        RECT 1450.540 1400.790 1450.680 1460.910 ;
        RECT 1450.480 1400.470 1450.740 1400.790 ;
        RECT 1450.480 1364.770 1450.740 1365.090 ;
        RECT 1450.540 1304.230 1450.680 1364.770 ;
        RECT 1450.480 1303.910 1450.740 1304.230 ;
        RECT 1450.480 1264.130 1450.740 1264.450 ;
        RECT 1450.540 883.050 1450.680 1264.130 ;
        RECT 1450.080 882.910 1450.680 883.050 ;
        RECT 1450.080 881.690 1450.220 882.910 ;
        RECT 1450.080 881.550 1450.680 881.690 ;
        RECT 1450.540 787.170 1450.680 881.550 ;
        RECT 1450.540 787.030 1451.140 787.170 ;
        RECT 1451.000 786.660 1451.140 787.030 ;
        RECT 1450.540 786.520 1451.140 786.660 ;
        RECT 1450.540 772.810 1450.680 786.520 ;
        RECT 1450.480 772.490 1450.740 772.810 ;
        RECT 1450.940 772.490 1451.200 772.810 ;
        RECT 1451.000 677.125 1451.140 772.490 ;
        RECT 1450.930 676.755 1451.210 677.125 ;
        RECT 1450.470 676.075 1450.750 676.445 ;
        RECT 1450.540 580.450 1450.680 676.075 ;
        RECT 1450.540 580.310 1451.140 580.450 ;
        RECT 1451.000 524.690 1451.140 580.310 ;
        RECT 1450.540 524.550 1451.140 524.690 ;
        RECT 1450.540 497.410 1450.680 524.550 ;
        RECT 1450.480 497.090 1450.740 497.410 ;
        RECT 1450.480 496.410 1450.740 496.730 ;
        RECT 1450.540 379.770 1450.680 496.410 ;
        RECT 1450.480 379.450 1450.740 379.770 ;
        RECT 1450.940 378.770 1451.200 379.090 ;
        RECT 1451.000 354.610 1451.140 378.770 ;
        RECT 1450.020 354.290 1450.280 354.610 ;
        RECT 1450.940 354.290 1451.200 354.610 ;
        RECT 1450.080 283.290 1450.220 354.290 ;
        RECT 1450.080 283.150 1450.680 283.290 ;
        RECT 1450.540 276.750 1450.680 283.150 ;
        RECT 1450.480 276.430 1450.740 276.750 ;
        RECT 1450.020 276.090 1450.280 276.410 ;
        RECT 1450.080 275.730 1450.220 276.090 ;
        RECT 1450.020 275.410 1450.280 275.730 ;
        RECT 1450.020 227.810 1450.280 228.130 ;
        RECT 1450.080 186.050 1450.220 227.810 ;
        RECT 1450.080 185.910 1450.680 186.050 ;
        RECT 1450.540 179.930 1450.680 185.910 ;
        RECT 1450.080 179.790 1450.680 179.930 ;
        RECT 1450.080 179.510 1450.220 179.790 ;
        RECT 1450.020 179.190 1450.280 179.510 ;
        RECT 1450.940 131.250 1451.200 131.570 ;
        RECT 1451.000 130.290 1451.140 131.250 ;
        RECT 1450.540 130.150 1451.140 130.290 ;
        RECT 1450.540 62.550 1450.680 130.150 ;
        RECT 1450.480 62.230 1450.740 62.550 ;
        RECT 811.540 60.870 811.800 61.190 ;
        RECT 811.600 2.400 811.740 60.870 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 1450.930 676.800 1451.210 677.080 ;
        RECT 1450.470 676.120 1450.750 676.400 ;
      LAYER met3 ;
        RECT 1450.905 677.090 1451.235 677.105 ;
        RECT 1450.230 676.790 1451.235 677.090 ;
        RECT 1450.230 676.425 1450.530 676.790 ;
        RECT 1450.905 676.775 1451.235 676.790 ;
        RECT 1450.230 676.110 1450.775 676.425 ;
        RECT 1450.445 676.095 1450.775 676.110 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2128.490 1688.680 2128.810 1688.740 ;
        RECT 2131.710 1688.680 2132.030 1688.740 ;
        RECT 2128.490 1688.540 2132.030 1688.680 ;
        RECT 2128.490 1688.480 2128.810 1688.540 ;
        RECT 2131.710 1688.480 2132.030 1688.540 ;
        RECT 2131.250 22.000 2131.570 22.060 ;
        RECT 2595.390 22.000 2595.710 22.060 ;
        RECT 2131.250 21.860 2595.710 22.000 ;
        RECT 2131.250 21.800 2131.570 21.860 ;
        RECT 2595.390 21.800 2595.710 21.860 ;
      LAYER via ;
        RECT 2128.520 1688.480 2128.780 1688.740 ;
        RECT 2131.740 1688.480 2132.000 1688.740 ;
        RECT 2131.280 21.800 2131.540 22.060 ;
        RECT 2595.420 21.800 2595.680 22.060 ;
      LAYER met2 ;
        RECT 2128.445 1700.000 2128.725 1704.000 ;
        RECT 2128.580 1688.770 2128.720 1700.000 ;
        RECT 2128.520 1688.450 2128.780 1688.770 ;
        RECT 2131.740 1688.450 2132.000 1688.770 ;
        RECT 2131.800 28.290 2131.940 1688.450 ;
        RECT 2131.340 28.150 2131.940 28.290 ;
        RECT 2131.340 22.090 2131.480 28.150 ;
        RECT 2131.280 21.770 2131.540 22.090 ;
        RECT 2595.420 21.770 2595.680 22.090 ;
        RECT 2595.480 2.400 2595.620 21.770 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2135.390 1688.680 2135.710 1688.740 ;
        RECT 2138.610 1688.680 2138.930 1688.740 ;
        RECT 2135.390 1688.540 2138.930 1688.680 ;
        RECT 2135.390 1688.480 2135.710 1688.540 ;
        RECT 2138.610 1688.480 2138.930 1688.540 ;
        RECT 2138.610 22.340 2138.930 22.400 ;
        RECT 2613.330 22.340 2613.650 22.400 ;
        RECT 2138.610 22.200 2613.650 22.340 ;
        RECT 2138.610 22.140 2138.930 22.200 ;
        RECT 2613.330 22.140 2613.650 22.200 ;
      LAYER via ;
        RECT 2135.420 1688.480 2135.680 1688.740 ;
        RECT 2138.640 1688.480 2138.900 1688.740 ;
        RECT 2138.640 22.140 2138.900 22.400 ;
        RECT 2613.360 22.140 2613.620 22.400 ;
      LAYER met2 ;
        RECT 2135.345 1700.000 2135.625 1704.000 ;
        RECT 2135.480 1688.770 2135.620 1700.000 ;
        RECT 2135.420 1688.450 2135.680 1688.770 ;
        RECT 2138.640 1688.450 2138.900 1688.770 ;
        RECT 2138.700 22.430 2138.840 1688.450 ;
        RECT 2138.640 22.110 2138.900 22.430 ;
        RECT 2613.360 22.110 2613.620 22.430 ;
        RECT 2613.420 2.400 2613.560 22.110 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2141.830 1686.980 2142.150 1687.040 ;
        RECT 2145.510 1686.980 2145.830 1687.040 ;
        RECT 2141.830 1686.840 2145.830 1686.980 ;
        RECT 2141.830 1686.780 2142.150 1686.840 ;
        RECT 2145.510 1686.780 2145.830 1686.840 ;
        RECT 2145.510 22.680 2145.830 22.740 ;
        RECT 2631.270 22.680 2631.590 22.740 ;
        RECT 2145.510 22.540 2631.590 22.680 ;
        RECT 2145.510 22.480 2145.830 22.540 ;
        RECT 2631.270 22.480 2631.590 22.540 ;
      LAYER via ;
        RECT 2141.860 1686.780 2142.120 1687.040 ;
        RECT 2145.540 1686.780 2145.800 1687.040 ;
        RECT 2145.540 22.480 2145.800 22.740 ;
        RECT 2631.300 22.480 2631.560 22.740 ;
      LAYER met2 ;
        RECT 2141.785 1700.000 2142.065 1704.000 ;
        RECT 2141.920 1687.070 2142.060 1700.000 ;
        RECT 2141.860 1686.750 2142.120 1687.070 ;
        RECT 2145.540 1686.750 2145.800 1687.070 ;
        RECT 2145.600 22.770 2145.740 1686.750 ;
        RECT 2145.540 22.450 2145.800 22.770 ;
        RECT 2631.300 22.450 2631.560 22.770 ;
        RECT 2631.360 2.400 2631.500 22.450 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2148.730 1686.980 2149.050 1687.040 ;
        RECT 2152.410 1686.980 2152.730 1687.040 ;
        RECT 2148.730 1686.840 2152.730 1686.980 ;
        RECT 2148.730 1686.780 2149.050 1686.840 ;
        RECT 2152.410 1686.780 2152.730 1686.840 ;
        RECT 2152.410 23.020 2152.730 23.080 ;
        RECT 2649.210 23.020 2649.530 23.080 ;
        RECT 2152.410 22.880 2649.530 23.020 ;
        RECT 2152.410 22.820 2152.730 22.880 ;
        RECT 2649.210 22.820 2649.530 22.880 ;
      LAYER via ;
        RECT 2148.760 1686.780 2149.020 1687.040 ;
        RECT 2152.440 1686.780 2152.700 1687.040 ;
        RECT 2152.440 22.820 2152.700 23.080 ;
        RECT 2649.240 22.820 2649.500 23.080 ;
      LAYER met2 ;
        RECT 2148.685 1700.000 2148.965 1704.000 ;
        RECT 2148.820 1687.070 2148.960 1700.000 ;
        RECT 2148.760 1686.750 2149.020 1687.070 ;
        RECT 2152.440 1686.750 2152.700 1687.070 ;
        RECT 2152.500 23.110 2152.640 1686.750 ;
        RECT 2152.440 22.790 2152.700 23.110 ;
        RECT 2649.240 22.790 2649.500 23.110 ;
        RECT 2649.300 2.400 2649.440 22.790 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2155.630 1686.980 2155.950 1687.040 ;
        RECT 2159.310 1686.980 2159.630 1687.040 ;
        RECT 2155.630 1686.840 2159.630 1686.980 ;
        RECT 2155.630 1686.780 2155.950 1686.840 ;
        RECT 2159.310 1686.780 2159.630 1686.840 ;
        RECT 2159.310 23.360 2159.630 23.420 ;
        RECT 2667.150 23.360 2667.470 23.420 ;
        RECT 2159.310 23.220 2667.470 23.360 ;
        RECT 2159.310 23.160 2159.630 23.220 ;
        RECT 2667.150 23.160 2667.470 23.220 ;
      LAYER via ;
        RECT 2155.660 1686.780 2155.920 1687.040 ;
        RECT 2159.340 1686.780 2159.600 1687.040 ;
        RECT 2159.340 23.160 2159.600 23.420 ;
        RECT 2667.180 23.160 2667.440 23.420 ;
      LAYER met2 ;
        RECT 2155.585 1700.000 2155.865 1704.000 ;
        RECT 2155.720 1687.070 2155.860 1700.000 ;
        RECT 2155.660 1686.750 2155.920 1687.070 ;
        RECT 2159.340 1686.750 2159.600 1687.070 ;
        RECT 2159.400 23.450 2159.540 1686.750 ;
        RECT 2159.340 23.130 2159.600 23.450 ;
        RECT 2667.180 23.130 2667.440 23.450 ;
        RECT 2667.240 2.400 2667.380 23.130 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2162.070 1686.980 2162.390 1687.040 ;
        RECT 2166.210 1686.980 2166.530 1687.040 ;
        RECT 2162.070 1686.840 2166.530 1686.980 ;
        RECT 2162.070 1686.780 2162.390 1686.840 ;
        RECT 2166.210 1686.780 2166.530 1686.840 ;
        RECT 2166.210 23.700 2166.530 23.760 ;
        RECT 2684.630 23.700 2684.950 23.760 ;
        RECT 2166.210 23.560 2684.950 23.700 ;
        RECT 2166.210 23.500 2166.530 23.560 ;
        RECT 2684.630 23.500 2684.950 23.560 ;
      LAYER via ;
        RECT 2162.100 1686.780 2162.360 1687.040 ;
        RECT 2166.240 1686.780 2166.500 1687.040 ;
        RECT 2166.240 23.500 2166.500 23.760 ;
        RECT 2684.660 23.500 2684.920 23.760 ;
      LAYER met2 ;
        RECT 2162.025 1700.000 2162.305 1704.000 ;
        RECT 2162.160 1687.070 2162.300 1700.000 ;
        RECT 2162.100 1686.750 2162.360 1687.070 ;
        RECT 2166.240 1686.750 2166.500 1687.070 ;
        RECT 2166.300 23.790 2166.440 1686.750 ;
        RECT 2166.240 23.470 2166.500 23.790 ;
        RECT 2684.660 23.470 2684.920 23.790 ;
        RECT 2684.720 2.400 2684.860 23.470 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2168.970 1686.980 2169.290 1687.040 ;
        RECT 2173.110 1686.980 2173.430 1687.040 ;
        RECT 2168.970 1686.840 2173.430 1686.980 ;
        RECT 2168.970 1686.780 2169.290 1686.840 ;
        RECT 2173.110 1686.780 2173.430 1686.840 ;
        RECT 2173.110 436.600 2173.430 436.860 ;
        RECT 2173.200 435.840 2173.340 436.600 ;
        RECT 2173.110 435.580 2173.430 435.840 ;
        RECT 2173.110 85.040 2173.430 85.300 ;
        RECT 2173.200 84.280 2173.340 85.040 ;
        RECT 2173.110 84.020 2173.430 84.280 ;
        RECT 2173.110 27.440 2173.430 27.500 ;
        RECT 2702.570 27.440 2702.890 27.500 ;
        RECT 2173.110 27.300 2702.890 27.440 ;
        RECT 2173.110 27.240 2173.430 27.300 ;
        RECT 2702.570 27.240 2702.890 27.300 ;
      LAYER via ;
        RECT 2169.000 1686.780 2169.260 1687.040 ;
        RECT 2173.140 1686.780 2173.400 1687.040 ;
        RECT 2173.140 436.600 2173.400 436.860 ;
        RECT 2173.140 435.580 2173.400 435.840 ;
        RECT 2173.140 85.040 2173.400 85.300 ;
        RECT 2173.140 84.020 2173.400 84.280 ;
        RECT 2173.140 27.240 2173.400 27.500 ;
        RECT 2702.600 27.240 2702.860 27.500 ;
      LAYER met2 ;
        RECT 2168.925 1700.000 2169.205 1704.000 ;
        RECT 2169.060 1687.070 2169.200 1700.000 ;
        RECT 2169.000 1686.750 2169.260 1687.070 ;
        RECT 2173.140 1686.750 2173.400 1687.070 ;
        RECT 2173.200 436.890 2173.340 1686.750 ;
        RECT 2173.140 436.570 2173.400 436.890 ;
        RECT 2173.140 435.550 2173.400 435.870 ;
        RECT 2173.200 85.330 2173.340 435.550 ;
        RECT 2173.140 85.010 2173.400 85.330 ;
        RECT 2173.140 83.990 2173.400 84.310 ;
        RECT 2173.200 27.530 2173.340 83.990 ;
        RECT 2173.140 27.210 2173.400 27.530 ;
        RECT 2702.600 27.210 2702.860 27.530 ;
        RECT 2702.660 2.400 2702.800 27.210 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2177.250 1678.140 2177.570 1678.200 ;
        RECT 2180.010 1678.140 2180.330 1678.200 ;
        RECT 2177.250 1678.000 2180.330 1678.140 ;
        RECT 2177.250 1677.940 2177.570 1678.000 ;
        RECT 2180.010 1677.940 2180.330 1678.000 ;
        RECT 2180.010 27.100 2180.330 27.160 ;
        RECT 2720.510 27.100 2720.830 27.160 ;
        RECT 2180.010 26.960 2720.830 27.100 ;
        RECT 2180.010 26.900 2180.330 26.960 ;
        RECT 2720.510 26.900 2720.830 26.960 ;
      LAYER via ;
        RECT 2177.280 1677.940 2177.540 1678.200 ;
        RECT 2180.040 1677.940 2180.300 1678.200 ;
        RECT 2180.040 26.900 2180.300 27.160 ;
        RECT 2720.540 26.900 2720.800 27.160 ;
      LAYER met2 ;
        RECT 2175.365 1700.410 2175.645 1704.000 ;
        RECT 2175.365 1700.270 2177.480 1700.410 ;
        RECT 2175.365 1700.000 2175.645 1700.270 ;
        RECT 2177.340 1678.230 2177.480 1700.270 ;
        RECT 2177.280 1677.910 2177.540 1678.230 ;
        RECT 2180.040 1677.910 2180.300 1678.230 ;
        RECT 2180.100 27.190 2180.240 1677.910 ;
        RECT 2180.040 26.870 2180.300 27.190 ;
        RECT 2720.540 26.870 2720.800 27.190 ;
        RECT 2720.600 2.400 2720.740 26.870 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2182.310 1688.340 2182.630 1688.400 ;
        RECT 2186.910 1688.340 2187.230 1688.400 ;
        RECT 2182.310 1688.200 2187.230 1688.340 ;
        RECT 2182.310 1688.140 2182.630 1688.200 ;
        RECT 2186.910 1688.140 2187.230 1688.200 ;
        RECT 2186.910 26.760 2187.230 26.820 ;
        RECT 2738.450 26.760 2738.770 26.820 ;
        RECT 2186.910 26.620 2738.770 26.760 ;
        RECT 2186.910 26.560 2187.230 26.620 ;
        RECT 2738.450 26.560 2738.770 26.620 ;
      LAYER via ;
        RECT 2182.340 1688.140 2182.600 1688.400 ;
        RECT 2186.940 1688.140 2187.200 1688.400 ;
        RECT 2186.940 26.560 2187.200 26.820 ;
        RECT 2738.480 26.560 2738.740 26.820 ;
      LAYER met2 ;
        RECT 2182.265 1700.000 2182.545 1704.000 ;
        RECT 2182.400 1688.430 2182.540 1700.000 ;
        RECT 2182.340 1688.110 2182.600 1688.430 ;
        RECT 2186.940 1688.110 2187.200 1688.430 ;
        RECT 2187.000 26.850 2187.140 1688.110 ;
        RECT 2186.940 26.530 2187.200 26.850 ;
        RECT 2738.480 26.530 2738.740 26.850 ;
        RECT 2738.540 2.400 2738.680 26.530 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2189.210 1686.980 2189.530 1687.040 ;
        RECT 2193.810 1686.980 2194.130 1687.040 ;
        RECT 2189.210 1686.840 2194.130 1686.980 ;
        RECT 2189.210 1686.780 2189.530 1686.840 ;
        RECT 2193.810 1686.780 2194.130 1686.840 ;
        RECT 2193.810 26.420 2194.130 26.480 ;
        RECT 2755.930 26.420 2756.250 26.480 ;
        RECT 2193.810 26.280 2756.250 26.420 ;
        RECT 2193.810 26.220 2194.130 26.280 ;
        RECT 2755.930 26.220 2756.250 26.280 ;
      LAYER via ;
        RECT 2189.240 1686.780 2189.500 1687.040 ;
        RECT 2193.840 1686.780 2194.100 1687.040 ;
        RECT 2193.840 26.220 2194.100 26.480 ;
        RECT 2755.960 26.220 2756.220 26.480 ;
      LAYER met2 ;
        RECT 2189.165 1700.000 2189.445 1704.000 ;
        RECT 2189.300 1687.070 2189.440 1700.000 ;
        RECT 2189.240 1686.750 2189.500 1687.070 ;
        RECT 2193.840 1686.750 2194.100 1687.070 ;
        RECT 2193.900 26.510 2194.040 1686.750 ;
        RECT 2193.840 26.190 2194.100 26.510 ;
        RECT 2755.960 26.190 2756.220 26.510 ;
        RECT 2756.020 2.400 2756.160 26.190 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1457.425 1442.025 1457.595 1490.475 ;
        RECT 1457.425 1256.385 1457.595 1304.155 ;
        RECT 1457.425 1207.425 1457.595 1255.875 ;
        RECT 1456.965 1014.645 1457.135 1103.895 ;
        RECT 1457.885 607.325 1458.055 621.095 ;
        RECT 1457.425 331.245 1457.595 396.695 ;
      LAYER mcon ;
        RECT 1457.425 1490.305 1457.595 1490.475 ;
        RECT 1457.425 1303.985 1457.595 1304.155 ;
        RECT 1457.425 1255.705 1457.595 1255.875 ;
        RECT 1456.965 1103.725 1457.135 1103.895 ;
        RECT 1457.885 620.925 1458.055 621.095 ;
        RECT 1457.425 396.525 1457.595 396.695 ;
      LAYER met1 ;
        RECT 1457.810 1642.440 1458.130 1642.500 ;
        RECT 1460.570 1642.440 1460.890 1642.500 ;
        RECT 1457.810 1642.300 1460.890 1642.440 ;
        RECT 1457.810 1642.240 1458.130 1642.300 ;
        RECT 1460.570 1642.240 1460.890 1642.300 ;
        RECT 1457.350 1545.880 1457.670 1545.940 ;
        RECT 1457.810 1545.880 1458.130 1545.940 ;
        RECT 1457.350 1545.740 1458.130 1545.880 ;
        RECT 1457.350 1545.680 1457.670 1545.740 ;
        RECT 1457.810 1545.680 1458.130 1545.740 ;
        RECT 1457.350 1497.260 1457.670 1497.320 ;
        RECT 1457.810 1497.260 1458.130 1497.320 ;
        RECT 1457.350 1497.120 1458.130 1497.260 ;
        RECT 1457.350 1497.060 1457.670 1497.120 ;
        RECT 1457.810 1497.060 1458.130 1497.120 ;
        RECT 1457.350 1490.460 1457.670 1490.520 ;
        RECT 1457.155 1490.320 1457.670 1490.460 ;
        RECT 1457.350 1490.260 1457.670 1490.320 ;
        RECT 1457.350 1442.180 1457.670 1442.240 ;
        RECT 1457.155 1442.040 1457.670 1442.180 ;
        RECT 1457.350 1441.980 1457.670 1442.040 ;
        RECT 1457.350 1400.700 1457.670 1400.760 ;
        RECT 1457.810 1400.700 1458.130 1400.760 ;
        RECT 1457.350 1400.560 1458.130 1400.700 ;
        RECT 1457.350 1400.500 1457.670 1400.560 ;
        RECT 1457.810 1400.500 1458.130 1400.560 ;
        RECT 1457.350 1345.620 1457.670 1345.680 ;
        RECT 1458.270 1345.620 1458.590 1345.680 ;
        RECT 1457.350 1345.480 1458.590 1345.620 ;
        RECT 1457.350 1345.420 1457.670 1345.480 ;
        RECT 1458.270 1345.420 1458.590 1345.480 ;
        RECT 1457.350 1317.880 1457.670 1318.140 ;
        RECT 1457.440 1317.400 1457.580 1317.880 ;
        RECT 1457.810 1317.400 1458.130 1317.460 ;
        RECT 1457.440 1317.260 1458.130 1317.400 ;
        RECT 1457.810 1317.200 1458.130 1317.260 ;
        RECT 1457.365 1304.140 1457.655 1304.185 ;
        RECT 1457.810 1304.140 1458.130 1304.200 ;
        RECT 1457.365 1304.000 1458.130 1304.140 ;
        RECT 1457.365 1303.955 1457.655 1304.000 ;
        RECT 1457.810 1303.940 1458.130 1304.000 ;
        RECT 1457.350 1256.540 1457.670 1256.600 ;
        RECT 1457.155 1256.400 1457.670 1256.540 ;
        RECT 1457.350 1256.340 1457.670 1256.400 ;
        RECT 1457.350 1255.860 1457.670 1255.920 ;
        RECT 1457.155 1255.720 1457.670 1255.860 ;
        RECT 1457.350 1255.660 1457.670 1255.720 ;
        RECT 1457.365 1207.580 1457.655 1207.625 ;
        RECT 1457.810 1207.580 1458.130 1207.640 ;
        RECT 1457.365 1207.440 1458.130 1207.580 ;
        RECT 1457.365 1207.395 1457.655 1207.440 ;
        RECT 1457.810 1207.380 1458.130 1207.440 ;
        RECT 1457.810 1152.500 1458.130 1152.560 ;
        RECT 1458.270 1152.500 1458.590 1152.560 ;
        RECT 1457.810 1152.360 1458.590 1152.500 ;
        RECT 1457.810 1152.300 1458.130 1152.360 ;
        RECT 1458.270 1152.300 1458.590 1152.360 ;
        RECT 1456.890 1104.560 1457.210 1104.620 ;
        RECT 1458.730 1104.560 1459.050 1104.620 ;
        RECT 1456.890 1104.420 1459.050 1104.560 ;
        RECT 1456.890 1104.360 1457.210 1104.420 ;
        RECT 1458.730 1104.360 1459.050 1104.420 ;
        RECT 1456.890 1103.880 1457.210 1103.940 ;
        RECT 1456.695 1103.740 1457.210 1103.880 ;
        RECT 1456.890 1103.680 1457.210 1103.740 ;
        RECT 1456.890 1014.800 1457.210 1014.860 ;
        RECT 1456.695 1014.660 1457.210 1014.800 ;
        RECT 1456.890 1014.600 1457.210 1014.660 ;
        RECT 1456.890 1007.320 1457.210 1007.380 ;
        RECT 1458.270 1007.320 1458.590 1007.380 ;
        RECT 1456.890 1007.180 1458.590 1007.320 ;
        RECT 1456.890 1007.120 1457.210 1007.180 ;
        RECT 1458.270 1007.120 1458.590 1007.180 ;
        RECT 1456.890 869.620 1457.210 869.680 ;
        RECT 1457.350 869.620 1457.670 869.680 ;
        RECT 1456.890 869.480 1457.670 869.620 ;
        RECT 1456.890 869.420 1457.210 869.480 ;
        RECT 1457.350 869.420 1457.670 869.480 ;
        RECT 1457.810 621.080 1458.130 621.140 ;
        RECT 1457.615 620.940 1458.130 621.080 ;
        RECT 1457.810 620.880 1458.130 620.940 ;
        RECT 1457.810 607.480 1458.130 607.540 ;
        RECT 1457.615 607.340 1458.130 607.480 ;
        RECT 1457.810 607.280 1458.130 607.340 ;
        RECT 1457.350 421.160 1457.670 421.220 ;
        RECT 1457.810 421.160 1458.130 421.220 ;
        RECT 1457.350 421.020 1458.130 421.160 ;
        RECT 1457.350 420.960 1457.670 421.020 ;
        RECT 1457.810 420.960 1458.130 421.020 ;
        RECT 1457.365 396.680 1457.655 396.725 ;
        RECT 1457.810 396.680 1458.130 396.740 ;
        RECT 1457.365 396.540 1458.130 396.680 ;
        RECT 1457.365 396.495 1457.655 396.540 ;
        RECT 1457.810 396.480 1458.130 396.540 ;
        RECT 1457.365 331.400 1457.655 331.445 ;
        RECT 1457.365 331.260 1458.040 331.400 ;
        RECT 1457.365 331.215 1457.655 331.260 ;
        RECT 1457.350 330.720 1457.670 330.780 ;
        RECT 1457.900 330.720 1458.040 331.260 ;
        RECT 1457.350 330.580 1458.040 330.720 ;
        RECT 1457.350 330.520 1457.670 330.580 ;
        RECT 1457.350 234.840 1457.670 234.900 ;
        RECT 1457.810 234.840 1458.130 234.900 ;
        RECT 1457.350 234.700 1458.130 234.840 ;
        RECT 1457.350 234.640 1457.670 234.700 ;
        RECT 1457.810 234.640 1458.130 234.700 ;
        RECT 829.450 61.440 829.770 61.500 ;
        RECT 1458.270 61.440 1458.590 61.500 ;
        RECT 829.450 61.300 1458.590 61.440 ;
        RECT 829.450 61.240 829.770 61.300 ;
        RECT 1458.270 61.240 1458.590 61.300 ;
      LAYER via ;
        RECT 1457.840 1642.240 1458.100 1642.500 ;
        RECT 1460.600 1642.240 1460.860 1642.500 ;
        RECT 1457.380 1545.680 1457.640 1545.940 ;
        RECT 1457.840 1545.680 1458.100 1545.940 ;
        RECT 1457.380 1497.060 1457.640 1497.320 ;
        RECT 1457.840 1497.060 1458.100 1497.320 ;
        RECT 1457.380 1490.260 1457.640 1490.520 ;
        RECT 1457.380 1441.980 1457.640 1442.240 ;
        RECT 1457.380 1400.500 1457.640 1400.760 ;
        RECT 1457.840 1400.500 1458.100 1400.760 ;
        RECT 1457.380 1345.420 1457.640 1345.680 ;
        RECT 1458.300 1345.420 1458.560 1345.680 ;
        RECT 1457.380 1317.880 1457.640 1318.140 ;
        RECT 1457.840 1317.200 1458.100 1317.460 ;
        RECT 1457.840 1303.940 1458.100 1304.200 ;
        RECT 1457.380 1256.340 1457.640 1256.600 ;
        RECT 1457.380 1255.660 1457.640 1255.920 ;
        RECT 1457.840 1207.380 1458.100 1207.640 ;
        RECT 1457.840 1152.300 1458.100 1152.560 ;
        RECT 1458.300 1152.300 1458.560 1152.560 ;
        RECT 1456.920 1104.360 1457.180 1104.620 ;
        RECT 1458.760 1104.360 1459.020 1104.620 ;
        RECT 1456.920 1103.680 1457.180 1103.940 ;
        RECT 1456.920 1014.600 1457.180 1014.860 ;
        RECT 1456.920 1007.120 1457.180 1007.380 ;
        RECT 1458.300 1007.120 1458.560 1007.380 ;
        RECT 1456.920 869.420 1457.180 869.680 ;
        RECT 1457.380 869.420 1457.640 869.680 ;
        RECT 1457.840 620.880 1458.100 621.140 ;
        RECT 1457.840 607.280 1458.100 607.540 ;
        RECT 1457.380 420.960 1457.640 421.220 ;
        RECT 1457.840 420.960 1458.100 421.220 ;
        RECT 1457.840 396.480 1458.100 396.740 ;
        RECT 1457.380 330.520 1457.640 330.780 ;
        RECT 1457.380 234.640 1457.640 234.900 ;
        RECT 1457.840 234.640 1458.100 234.900 ;
        RECT 829.480 61.240 829.740 61.500 ;
        RECT 1458.300 61.240 1458.560 61.500 ;
      LAYER met2 ;
        RECT 1461.905 1700.410 1462.185 1704.000 ;
        RECT 1460.660 1700.270 1462.185 1700.410 ;
        RECT 1460.660 1642.530 1460.800 1700.270 ;
        RECT 1461.905 1700.000 1462.185 1700.270 ;
        RECT 1457.840 1642.210 1458.100 1642.530 ;
        RECT 1460.600 1642.210 1460.860 1642.530 ;
        RECT 1457.900 1545.970 1458.040 1642.210 ;
        RECT 1457.380 1545.650 1457.640 1545.970 ;
        RECT 1457.840 1545.650 1458.100 1545.970 ;
        RECT 1457.440 1521.570 1457.580 1545.650 ;
        RECT 1457.440 1521.430 1458.040 1521.570 ;
        RECT 1457.900 1497.350 1458.040 1521.430 ;
        RECT 1457.380 1497.030 1457.640 1497.350 ;
        RECT 1457.840 1497.030 1458.100 1497.350 ;
        RECT 1457.440 1490.550 1457.580 1497.030 ;
        RECT 1457.380 1490.230 1457.640 1490.550 ;
        RECT 1457.380 1441.950 1457.640 1442.270 ;
        RECT 1457.440 1425.010 1457.580 1441.950 ;
        RECT 1456.980 1424.870 1457.580 1425.010 ;
        RECT 1456.980 1413.450 1457.120 1424.870 ;
        RECT 1456.980 1413.310 1458.040 1413.450 ;
        RECT 1457.900 1400.790 1458.040 1413.310 ;
        RECT 1457.380 1400.470 1457.640 1400.790 ;
        RECT 1457.840 1400.470 1458.100 1400.790 ;
        RECT 1457.440 1393.845 1457.580 1400.470 ;
        RECT 1457.370 1393.475 1457.650 1393.845 ;
        RECT 1458.290 1393.475 1458.570 1393.845 ;
        RECT 1458.360 1345.710 1458.500 1393.475 ;
        RECT 1457.380 1345.390 1457.640 1345.710 ;
        RECT 1458.300 1345.390 1458.560 1345.710 ;
        RECT 1457.440 1318.170 1457.580 1345.390 ;
        RECT 1457.380 1317.850 1457.640 1318.170 ;
        RECT 1457.840 1317.170 1458.100 1317.490 ;
        RECT 1457.900 1304.230 1458.040 1317.170 ;
        RECT 1457.840 1303.910 1458.100 1304.230 ;
        RECT 1457.380 1256.310 1457.640 1256.630 ;
        RECT 1457.440 1255.950 1457.580 1256.310 ;
        RECT 1457.380 1255.630 1457.640 1255.950 ;
        RECT 1457.840 1207.350 1458.100 1207.670 ;
        RECT 1457.900 1167.970 1458.040 1207.350 ;
        RECT 1457.900 1167.830 1458.500 1167.970 ;
        RECT 1458.360 1152.590 1458.500 1167.830 ;
        RECT 1457.840 1152.445 1458.100 1152.590 ;
        RECT 1457.830 1152.075 1458.110 1152.445 ;
        RECT 1458.300 1152.270 1458.560 1152.590 ;
        RECT 1458.750 1152.075 1459.030 1152.445 ;
        RECT 1458.820 1104.650 1458.960 1152.075 ;
        RECT 1456.920 1104.330 1457.180 1104.650 ;
        RECT 1458.760 1104.330 1459.020 1104.650 ;
        RECT 1456.980 1103.970 1457.120 1104.330 ;
        RECT 1456.920 1103.650 1457.180 1103.970 ;
        RECT 1456.920 1014.570 1457.180 1014.890 ;
        RECT 1456.980 1007.410 1457.120 1014.570 ;
        RECT 1456.920 1007.090 1457.180 1007.410 ;
        RECT 1458.300 1007.090 1458.560 1007.410 ;
        RECT 1458.360 931.330 1458.500 1007.090 ;
        RECT 1457.900 931.190 1458.500 931.330 ;
        RECT 1457.900 917.845 1458.040 931.190 ;
        RECT 1456.910 917.475 1457.190 917.845 ;
        RECT 1457.830 917.475 1458.110 917.845 ;
        RECT 1456.980 869.710 1457.120 917.475 ;
        RECT 1456.920 869.390 1457.180 869.710 ;
        RECT 1457.380 869.565 1457.640 869.710 ;
        RECT 1457.370 869.195 1457.650 869.565 ;
        RECT 1458.750 869.195 1459.030 869.565 ;
        RECT 1458.820 821.285 1458.960 869.195 ;
        RECT 1457.830 820.915 1458.110 821.285 ;
        RECT 1458.750 820.915 1459.030 821.285 ;
        RECT 1457.900 773.685 1458.040 820.915 ;
        RECT 1457.830 773.315 1458.110 773.685 ;
        RECT 1458.290 771.955 1458.570 772.325 ;
        RECT 1458.360 737.530 1458.500 771.955 ;
        RECT 1457.900 737.390 1458.500 737.530 ;
        RECT 1457.900 677.125 1458.040 737.390 ;
        RECT 1457.830 676.755 1458.110 677.125 ;
        RECT 1457.830 675.395 1458.110 675.765 ;
        RECT 1457.900 621.170 1458.040 675.395 ;
        RECT 1457.840 620.850 1458.100 621.170 ;
        RECT 1457.840 607.250 1458.100 607.570 ;
        RECT 1457.900 510.525 1458.040 607.250 ;
        RECT 1457.830 510.155 1458.110 510.525 ;
        RECT 1457.370 509.475 1457.650 509.845 ;
        RECT 1457.440 421.250 1457.580 509.475 ;
        RECT 1457.380 420.930 1457.640 421.250 ;
        RECT 1457.840 420.930 1458.100 421.250 ;
        RECT 1457.900 396.770 1458.040 420.930 ;
        RECT 1457.840 396.450 1458.100 396.770 ;
        RECT 1457.380 330.490 1457.640 330.810 ;
        RECT 1457.440 234.930 1457.580 330.490 ;
        RECT 1457.380 234.610 1457.640 234.930 ;
        RECT 1457.840 234.610 1458.100 234.930 ;
        RECT 1457.900 207.130 1458.040 234.610 ;
        RECT 1457.900 206.990 1458.500 207.130 ;
        RECT 1458.360 206.450 1458.500 206.990 ;
        RECT 1457.900 206.310 1458.500 206.450 ;
        RECT 1457.900 186.050 1458.040 206.310 ;
        RECT 1457.900 185.910 1458.500 186.050 ;
        RECT 1458.360 61.530 1458.500 185.910 ;
        RECT 829.480 61.210 829.740 61.530 ;
        RECT 1458.300 61.210 1458.560 61.530 ;
        RECT 829.540 2.400 829.680 61.210 ;
        RECT 829.330 -4.800 829.890 2.400 ;
      LAYER via2 ;
        RECT 1457.370 1393.520 1457.650 1393.800 ;
        RECT 1458.290 1393.520 1458.570 1393.800 ;
        RECT 1457.830 1152.120 1458.110 1152.400 ;
        RECT 1458.750 1152.120 1459.030 1152.400 ;
        RECT 1456.910 917.520 1457.190 917.800 ;
        RECT 1457.830 917.520 1458.110 917.800 ;
        RECT 1457.370 869.240 1457.650 869.520 ;
        RECT 1458.750 869.240 1459.030 869.520 ;
        RECT 1457.830 820.960 1458.110 821.240 ;
        RECT 1458.750 820.960 1459.030 821.240 ;
        RECT 1457.830 773.360 1458.110 773.640 ;
        RECT 1458.290 772.000 1458.570 772.280 ;
        RECT 1457.830 676.800 1458.110 677.080 ;
        RECT 1457.830 675.440 1458.110 675.720 ;
        RECT 1457.830 510.200 1458.110 510.480 ;
        RECT 1457.370 509.520 1457.650 509.800 ;
      LAYER met3 ;
        RECT 1457.345 1393.810 1457.675 1393.825 ;
        RECT 1458.265 1393.810 1458.595 1393.825 ;
        RECT 1457.345 1393.510 1458.595 1393.810 ;
        RECT 1457.345 1393.495 1457.675 1393.510 ;
        RECT 1458.265 1393.495 1458.595 1393.510 ;
        RECT 1457.805 1152.410 1458.135 1152.425 ;
        RECT 1458.725 1152.410 1459.055 1152.425 ;
        RECT 1457.805 1152.110 1459.055 1152.410 ;
        RECT 1457.805 1152.095 1458.135 1152.110 ;
        RECT 1458.725 1152.095 1459.055 1152.110 ;
        RECT 1456.885 917.810 1457.215 917.825 ;
        RECT 1457.805 917.810 1458.135 917.825 ;
        RECT 1456.885 917.510 1458.135 917.810 ;
        RECT 1456.885 917.495 1457.215 917.510 ;
        RECT 1457.805 917.495 1458.135 917.510 ;
        RECT 1457.345 869.530 1457.675 869.545 ;
        RECT 1458.725 869.530 1459.055 869.545 ;
        RECT 1457.345 869.230 1459.055 869.530 ;
        RECT 1457.345 869.215 1457.675 869.230 ;
        RECT 1458.725 869.215 1459.055 869.230 ;
        RECT 1457.805 821.250 1458.135 821.265 ;
        RECT 1458.725 821.250 1459.055 821.265 ;
        RECT 1457.805 820.950 1459.055 821.250 ;
        RECT 1457.805 820.935 1458.135 820.950 ;
        RECT 1458.725 820.935 1459.055 820.950 ;
        RECT 1457.805 773.650 1458.135 773.665 ;
        RECT 1457.590 773.335 1458.135 773.650 ;
        RECT 1457.590 772.290 1457.890 773.335 ;
        RECT 1458.265 772.290 1458.595 772.305 ;
        RECT 1457.590 771.990 1458.595 772.290 ;
        RECT 1458.265 771.975 1458.595 771.990 ;
        RECT 1457.805 677.090 1458.135 677.105 ;
        RECT 1457.590 676.775 1458.135 677.090 ;
        RECT 1457.590 675.745 1457.890 676.775 ;
        RECT 1457.590 675.430 1458.135 675.745 ;
        RECT 1457.805 675.415 1458.135 675.430 ;
        RECT 1457.805 510.490 1458.135 510.505 ;
        RECT 1457.805 510.190 1458.810 510.490 ;
        RECT 1457.805 510.175 1458.135 510.190 ;
        RECT 1457.345 509.810 1457.675 509.825 ;
        RECT 1458.510 509.810 1458.810 510.190 ;
        RECT 1457.345 509.510 1458.810 509.810 ;
        RECT 1457.345 509.495 1457.675 509.510 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2195.650 1686.980 2195.970 1687.040 ;
        RECT 2200.250 1686.980 2200.570 1687.040 ;
        RECT 2195.650 1686.840 2200.570 1686.980 ;
        RECT 2195.650 1686.780 2195.970 1686.840 ;
        RECT 2200.250 1686.780 2200.570 1686.840 ;
        RECT 2200.250 26.080 2200.570 26.140 ;
        RECT 2773.870 26.080 2774.190 26.140 ;
        RECT 2200.250 25.940 2774.190 26.080 ;
        RECT 2200.250 25.880 2200.570 25.940 ;
        RECT 2773.870 25.880 2774.190 25.940 ;
      LAYER via ;
        RECT 2195.680 1686.780 2195.940 1687.040 ;
        RECT 2200.280 1686.780 2200.540 1687.040 ;
        RECT 2200.280 25.880 2200.540 26.140 ;
        RECT 2773.900 25.880 2774.160 26.140 ;
      LAYER met2 ;
        RECT 2195.605 1700.000 2195.885 1704.000 ;
        RECT 2195.740 1687.070 2195.880 1700.000 ;
        RECT 2195.680 1686.750 2195.940 1687.070 ;
        RECT 2200.280 1686.750 2200.540 1687.070 ;
        RECT 2200.340 26.170 2200.480 1686.750 ;
        RECT 2200.280 25.850 2200.540 26.170 ;
        RECT 2773.900 25.850 2774.160 26.170 ;
        RECT 2773.960 2.400 2774.100 25.850 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2202.550 1686.980 2202.870 1687.040 ;
        RECT 2207.610 1686.980 2207.930 1687.040 ;
        RECT 2202.550 1686.840 2207.930 1686.980 ;
        RECT 2202.550 1686.780 2202.870 1686.840 ;
        RECT 2207.610 1686.780 2207.930 1686.840 ;
        RECT 2207.610 25.740 2207.930 25.800 ;
        RECT 2791.810 25.740 2792.130 25.800 ;
        RECT 2207.610 25.600 2792.130 25.740 ;
        RECT 2207.610 25.540 2207.930 25.600 ;
        RECT 2791.810 25.540 2792.130 25.600 ;
      LAYER via ;
        RECT 2202.580 1686.780 2202.840 1687.040 ;
        RECT 2207.640 1686.780 2207.900 1687.040 ;
        RECT 2207.640 25.540 2207.900 25.800 ;
        RECT 2791.840 25.540 2792.100 25.800 ;
      LAYER met2 ;
        RECT 2202.505 1700.000 2202.785 1704.000 ;
        RECT 2202.640 1687.070 2202.780 1700.000 ;
        RECT 2202.580 1686.750 2202.840 1687.070 ;
        RECT 2207.640 1686.750 2207.900 1687.070 ;
        RECT 2207.700 25.830 2207.840 1686.750 ;
        RECT 2207.640 25.510 2207.900 25.830 ;
        RECT 2791.840 25.510 2792.100 25.830 ;
        RECT 2791.900 2.400 2792.040 25.510 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2209.450 1686.980 2209.770 1687.040 ;
        RECT 2214.050 1686.980 2214.370 1687.040 ;
        RECT 2209.450 1686.840 2214.370 1686.980 ;
        RECT 2209.450 1686.780 2209.770 1686.840 ;
        RECT 2214.050 1686.780 2214.370 1686.840 ;
        RECT 2214.050 25.400 2214.370 25.460 ;
        RECT 2809.750 25.400 2810.070 25.460 ;
        RECT 2214.050 25.260 2810.070 25.400 ;
        RECT 2214.050 25.200 2214.370 25.260 ;
        RECT 2809.750 25.200 2810.070 25.260 ;
      LAYER via ;
        RECT 2209.480 1686.780 2209.740 1687.040 ;
        RECT 2214.080 1686.780 2214.340 1687.040 ;
        RECT 2214.080 25.200 2214.340 25.460 ;
        RECT 2809.780 25.200 2810.040 25.460 ;
      LAYER met2 ;
        RECT 2209.405 1700.000 2209.685 1704.000 ;
        RECT 2209.540 1687.070 2209.680 1700.000 ;
        RECT 2209.480 1686.750 2209.740 1687.070 ;
        RECT 2214.080 1686.750 2214.340 1687.070 ;
        RECT 2214.140 25.490 2214.280 1686.750 ;
        RECT 2214.080 25.170 2214.340 25.490 ;
        RECT 2809.780 25.170 2810.040 25.490 ;
        RECT 2809.840 2.400 2809.980 25.170 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2215.890 1686.980 2216.210 1687.040 ;
        RECT 2221.410 1686.980 2221.730 1687.040 ;
        RECT 2215.890 1686.840 2221.730 1686.980 ;
        RECT 2215.890 1686.780 2216.210 1686.840 ;
        RECT 2221.410 1686.780 2221.730 1686.840 ;
        RECT 2221.410 25.060 2221.730 25.120 ;
        RECT 2827.690 25.060 2828.010 25.120 ;
        RECT 2221.410 24.920 2828.010 25.060 ;
        RECT 2221.410 24.860 2221.730 24.920 ;
        RECT 2827.690 24.860 2828.010 24.920 ;
      LAYER via ;
        RECT 2215.920 1686.780 2216.180 1687.040 ;
        RECT 2221.440 1686.780 2221.700 1687.040 ;
        RECT 2221.440 24.860 2221.700 25.120 ;
        RECT 2827.720 24.860 2827.980 25.120 ;
      LAYER met2 ;
        RECT 2215.845 1700.000 2216.125 1704.000 ;
        RECT 2215.980 1687.070 2216.120 1700.000 ;
        RECT 2215.920 1686.750 2216.180 1687.070 ;
        RECT 2221.440 1686.750 2221.700 1687.070 ;
        RECT 2221.500 25.150 2221.640 1686.750 ;
        RECT 2221.440 24.830 2221.700 25.150 ;
        RECT 2827.720 24.830 2827.980 25.150 ;
        RECT 2827.780 2.400 2827.920 24.830 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2222.790 1686.980 2223.110 1687.040 ;
        RECT 2227.850 1686.980 2228.170 1687.040 ;
        RECT 2222.790 1686.840 2228.170 1686.980 ;
        RECT 2222.790 1686.780 2223.110 1686.840 ;
        RECT 2227.850 1686.780 2228.170 1686.840 ;
        RECT 2227.850 24.720 2228.170 24.780 ;
        RECT 2845.170 24.720 2845.490 24.780 ;
        RECT 2227.850 24.580 2845.490 24.720 ;
        RECT 2227.850 24.520 2228.170 24.580 ;
        RECT 2845.170 24.520 2845.490 24.580 ;
      LAYER via ;
        RECT 2222.820 1686.780 2223.080 1687.040 ;
        RECT 2227.880 1686.780 2228.140 1687.040 ;
        RECT 2227.880 24.520 2228.140 24.780 ;
        RECT 2845.200 24.520 2845.460 24.780 ;
      LAYER met2 ;
        RECT 2222.745 1700.000 2223.025 1704.000 ;
        RECT 2222.880 1687.070 2223.020 1700.000 ;
        RECT 2222.820 1686.750 2223.080 1687.070 ;
        RECT 2227.880 1686.750 2228.140 1687.070 ;
        RECT 2227.940 24.810 2228.080 1686.750 ;
        RECT 2227.880 24.490 2228.140 24.810 ;
        RECT 2845.200 24.490 2845.460 24.810 ;
        RECT 2845.260 2.400 2845.400 24.490 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2229.690 1688.340 2230.010 1688.400 ;
        RECT 2235.210 1688.340 2235.530 1688.400 ;
        RECT 2229.690 1688.200 2235.530 1688.340 ;
        RECT 2229.690 1688.140 2230.010 1688.200 ;
        RECT 2235.210 1688.140 2235.530 1688.200 ;
        RECT 2235.210 24.380 2235.530 24.440 ;
        RECT 2863.110 24.380 2863.430 24.440 ;
        RECT 2235.210 24.240 2863.430 24.380 ;
        RECT 2235.210 24.180 2235.530 24.240 ;
        RECT 2863.110 24.180 2863.430 24.240 ;
      LAYER via ;
        RECT 2229.720 1688.140 2229.980 1688.400 ;
        RECT 2235.240 1688.140 2235.500 1688.400 ;
        RECT 2235.240 24.180 2235.500 24.440 ;
        RECT 2863.140 24.180 2863.400 24.440 ;
      LAYER met2 ;
        RECT 2229.645 1700.000 2229.925 1704.000 ;
        RECT 2229.780 1688.430 2229.920 1700.000 ;
        RECT 2229.720 1688.110 2229.980 1688.430 ;
        RECT 2235.240 1688.110 2235.500 1688.430 ;
        RECT 2235.300 24.470 2235.440 1688.110 ;
        RECT 2235.240 24.150 2235.500 24.470 ;
        RECT 2863.140 24.150 2863.400 24.470 ;
        RECT 2863.200 2.400 2863.340 24.150 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2236.130 1688.340 2236.450 1688.400 ;
        RECT 2242.110 1688.340 2242.430 1688.400 ;
        RECT 2236.130 1688.200 2242.430 1688.340 ;
        RECT 2236.130 1688.140 2236.450 1688.200 ;
        RECT 2242.110 1688.140 2242.430 1688.200 ;
        RECT 2242.110 24.040 2242.430 24.100 ;
        RECT 2881.050 24.040 2881.370 24.100 ;
        RECT 2242.110 23.900 2881.370 24.040 ;
        RECT 2242.110 23.840 2242.430 23.900 ;
        RECT 2881.050 23.840 2881.370 23.900 ;
      LAYER via ;
        RECT 2236.160 1688.140 2236.420 1688.400 ;
        RECT 2242.140 1688.140 2242.400 1688.400 ;
        RECT 2242.140 23.840 2242.400 24.100 ;
        RECT 2881.080 23.840 2881.340 24.100 ;
      LAYER met2 ;
        RECT 2236.085 1700.000 2236.365 1704.000 ;
        RECT 2236.220 1688.430 2236.360 1700.000 ;
        RECT 2236.160 1688.110 2236.420 1688.430 ;
        RECT 2242.140 1688.110 2242.400 1688.430 ;
        RECT 2242.200 24.130 2242.340 1688.110 ;
        RECT 2242.140 23.810 2242.400 24.130 ;
        RECT 2881.080 23.810 2881.340 24.130 ;
        RECT 2881.140 2.400 2881.280 23.810 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2243.030 1688.340 2243.350 1688.400 ;
        RECT 2249.010 1688.340 2249.330 1688.400 ;
        RECT 2243.030 1688.200 2249.330 1688.340 ;
        RECT 2243.030 1688.140 2243.350 1688.200 ;
        RECT 2249.010 1688.140 2249.330 1688.200 ;
      LAYER via ;
        RECT 2243.060 1688.140 2243.320 1688.400 ;
        RECT 2249.040 1688.140 2249.300 1688.400 ;
      LAYER met2 ;
        RECT 2242.985 1700.000 2243.265 1704.000 ;
        RECT 2243.120 1688.430 2243.260 1700.000 ;
        RECT 2243.060 1688.110 2243.320 1688.430 ;
        RECT 2249.040 1688.110 2249.300 1688.430 ;
        RECT 2249.100 24.325 2249.240 1688.110 ;
        RECT 2249.030 23.955 2249.310 24.325 ;
        RECT 2899.010 23.955 2899.290 24.325 ;
        RECT 2899.080 2.400 2899.220 23.955 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 2249.030 24.000 2249.310 24.280 ;
        RECT 2899.010 24.000 2899.290 24.280 ;
      LAYER met3 ;
        RECT 2249.005 24.290 2249.335 24.305 ;
        RECT 2898.985 24.290 2899.315 24.305 ;
        RECT 2249.005 23.990 2899.315 24.290 ;
        RECT 2249.005 23.975 2249.335 23.990 ;
        RECT 2898.985 23.975 2899.315 23.990 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1464.325 1545.725 1464.495 1593.835 ;
        RECT 1463.865 131.325 1464.035 153.595 ;
      LAYER mcon ;
        RECT 1464.325 1593.665 1464.495 1593.835 ;
        RECT 1463.865 153.425 1464.035 153.595 ;
      LAYER met1 ;
        RECT 1463.790 1642.440 1464.110 1642.500 ;
        RECT 1467.930 1642.440 1468.250 1642.500 ;
        RECT 1463.790 1642.300 1468.250 1642.440 ;
        RECT 1463.790 1642.240 1464.110 1642.300 ;
        RECT 1467.930 1642.240 1468.250 1642.300 ;
        RECT 1463.790 1607.900 1464.110 1608.160 ;
        RECT 1463.880 1607.420 1464.020 1607.900 ;
        RECT 1464.250 1607.420 1464.570 1607.480 ;
        RECT 1463.880 1607.280 1464.570 1607.420 ;
        RECT 1464.250 1607.220 1464.570 1607.280 ;
        RECT 1464.250 1593.820 1464.570 1593.880 ;
        RECT 1464.055 1593.680 1464.570 1593.820 ;
        RECT 1464.250 1593.620 1464.570 1593.680 ;
        RECT 1464.250 1545.880 1464.570 1545.940 ;
        RECT 1464.055 1545.740 1464.570 1545.880 ;
        RECT 1464.250 1545.680 1464.570 1545.740 ;
        RECT 1464.250 593.680 1464.570 593.940 ;
        RECT 1464.340 593.260 1464.480 593.680 ;
        RECT 1464.250 593.000 1464.570 593.260 ;
        RECT 1463.790 324.260 1464.110 324.320 ;
        RECT 1464.250 324.260 1464.570 324.320 ;
        RECT 1463.790 324.120 1464.570 324.260 ;
        RECT 1463.790 324.060 1464.110 324.120 ;
        RECT 1464.250 324.060 1464.570 324.120 ;
        RECT 1463.805 153.580 1464.095 153.625 ;
        RECT 1464.250 153.580 1464.570 153.640 ;
        RECT 1463.805 153.440 1464.570 153.580 ;
        RECT 1463.805 153.395 1464.095 153.440 ;
        RECT 1464.250 153.380 1464.570 153.440 ;
        RECT 1463.790 131.480 1464.110 131.540 ;
        RECT 1463.595 131.340 1464.110 131.480 ;
        RECT 1463.790 131.280 1464.110 131.340 ;
        RECT 1463.790 96.800 1464.110 96.860 ;
        RECT 1464.250 96.800 1464.570 96.860 ;
        RECT 1463.790 96.660 1464.570 96.800 ;
        RECT 1463.790 96.600 1464.110 96.660 ;
        RECT 1464.250 96.600 1464.570 96.660 ;
        RECT 846.930 61.780 847.250 61.840 ;
        RECT 1464.710 61.780 1465.030 61.840 ;
        RECT 846.930 61.640 1465.030 61.780 ;
        RECT 846.930 61.580 847.250 61.640 ;
        RECT 1464.710 61.580 1465.030 61.640 ;
      LAYER via ;
        RECT 1463.820 1642.240 1464.080 1642.500 ;
        RECT 1467.960 1642.240 1468.220 1642.500 ;
        RECT 1463.820 1607.900 1464.080 1608.160 ;
        RECT 1464.280 1607.220 1464.540 1607.480 ;
        RECT 1464.280 1593.620 1464.540 1593.880 ;
        RECT 1464.280 1545.680 1464.540 1545.940 ;
        RECT 1464.280 593.680 1464.540 593.940 ;
        RECT 1464.280 593.000 1464.540 593.260 ;
        RECT 1463.820 324.060 1464.080 324.320 ;
        RECT 1464.280 324.060 1464.540 324.320 ;
        RECT 1464.280 153.380 1464.540 153.640 ;
        RECT 1463.820 131.280 1464.080 131.540 ;
        RECT 1463.820 96.600 1464.080 96.860 ;
        RECT 1464.280 96.600 1464.540 96.860 ;
        RECT 846.960 61.580 847.220 61.840 ;
        RECT 1464.740 61.580 1465.000 61.840 ;
      LAYER met2 ;
        RECT 1468.345 1700.410 1468.625 1704.000 ;
        RECT 1468.020 1700.270 1468.625 1700.410 ;
        RECT 1468.020 1642.530 1468.160 1700.270 ;
        RECT 1468.345 1700.000 1468.625 1700.270 ;
        RECT 1463.820 1642.210 1464.080 1642.530 ;
        RECT 1467.960 1642.210 1468.220 1642.530 ;
        RECT 1463.880 1608.190 1464.020 1642.210 ;
        RECT 1463.820 1607.870 1464.080 1608.190 ;
        RECT 1464.280 1607.190 1464.540 1607.510 ;
        RECT 1464.340 1593.910 1464.480 1607.190 ;
        RECT 1464.280 1593.590 1464.540 1593.910 ;
        RECT 1464.280 1545.650 1464.540 1545.970 ;
        RECT 1464.340 883.050 1464.480 1545.650 ;
        RECT 1463.880 882.910 1464.480 883.050 ;
        RECT 1463.880 881.690 1464.020 882.910 ;
        RECT 1463.880 881.550 1464.480 881.690 ;
        RECT 1464.340 593.970 1464.480 881.550 ;
        RECT 1464.280 593.650 1464.540 593.970 ;
        RECT 1464.280 592.970 1464.540 593.290 ;
        RECT 1464.340 497.490 1464.480 592.970 ;
        RECT 1463.880 497.350 1464.480 497.490 ;
        RECT 1463.880 496.810 1464.020 497.350 ;
        RECT 1463.880 496.670 1464.480 496.810 ;
        RECT 1464.340 400.930 1464.480 496.670 ;
        RECT 1464.340 400.790 1464.940 400.930 ;
        RECT 1464.800 400.080 1464.940 400.790 ;
        RECT 1464.340 399.940 1464.940 400.080 ;
        RECT 1464.340 355.370 1464.480 399.940 ;
        RECT 1463.880 355.230 1464.480 355.370 ;
        RECT 1463.880 324.350 1464.020 355.230 ;
        RECT 1463.820 324.030 1464.080 324.350 ;
        RECT 1464.280 324.030 1464.540 324.350 ;
        RECT 1464.340 235.010 1464.480 324.030 ;
        RECT 1463.880 234.870 1464.480 235.010 ;
        RECT 1463.880 203.730 1464.020 234.870 ;
        RECT 1463.880 203.590 1464.480 203.730 ;
        RECT 1464.340 153.670 1464.480 203.590 ;
        RECT 1464.280 153.350 1464.540 153.670 ;
        RECT 1463.820 131.250 1464.080 131.570 ;
        RECT 1463.880 96.890 1464.020 131.250 ;
        RECT 1463.820 96.570 1464.080 96.890 ;
        RECT 1464.280 96.570 1464.540 96.890 ;
        RECT 1464.340 62.290 1464.480 96.570 ;
        RECT 1464.340 62.150 1464.940 62.290 ;
        RECT 1464.800 61.870 1464.940 62.150 ;
        RECT 846.960 61.550 847.220 61.870 ;
        RECT 1464.740 61.550 1465.000 61.870 ;
        RECT 847.020 2.400 847.160 61.550 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1470.230 1678.140 1470.550 1678.200 ;
        RECT 1473.910 1678.140 1474.230 1678.200 ;
        RECT 1470.230 1678.000 1474.230 1678.140 ;
        RECT 1470.230 1677.940 1470.550 1678.000 ;
        RECT 1473.910 1677.940 1474.230 1678.000 ;
        RECT 869.010 62.120 869.330 62.180 ;
        RECT 1470.230 62.120 1470.550 62.180 ;
        RECT 869.010 61.980 1470.550 62.120 ;
        RECT 869.010 61.920 869.330 61.980 ;
        RECT 1470.230 61.920 1470.550 61.980 ;
        RECT 864.870 2.960 865.190 3.020 ;
        RECT 869.010 2.960 869.330 3.020 ;
        RECT 864.870 2.820 869.330 2.960 ;
        RECT 864.870 2.760 865.190 2.820 ;
        RECT 869.010 2.760 869.330 2.820 ;
      LAYER via ;
        RECT 1470.260 1677.940 1470.520 1678.200 ;
        RECT 1473.940 1677.940 1474.200 1678.200 ;
        RECT 869.040 61.920 869.300 62.180 ;
        RECT 1470.260 61.920 1470.520 62.180 ;
        RECT 864.900 2.760 865.160 3.020 ;
        RECT 869.040 2.760 869.300 3.020 ;
      LAYER met2 ;
        RECT 1475.245 1700.410 1475.525 1704.000 ;
        RECT 1474.000 1700.270 1475.525 1700.410 ;
        RECT 1474.000 1678.230 1474.140 1700.270 ;
        RECT 1475.245 1700.000 1475.525 1700.270 ;
        RECT 1470.260 1677.910 1470.520 1678.230 ;
        RECT 1473.940 1677.910 1474.200 1678.230 ;
        RECT 1470.320 62.210 1470.460 1677.910 ;
        RECT 869.040 61.890 869.300 62.210 ;
        RECT 1470.260 61.890 1470.520 62.210 ;
        RECT 869.100 3.050 869.240 61.890 ;
        RECT 864.900 2.730 865.160 3.050 ;
        RECT 869.040 2.730 869.300 3.050 ;
        RECT 864.960 2.400 865.100 2.730 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1477.130 1658.080 1477.450 1658.140 ;
        RECT 1480.350 1658.080 1480.670 1658.140 ;
        RECT 1477.130 1657.940 1480.670 1658.080 ;
        RECT 1477.130 1657.880 1477.450 1657.940 ;
        RECT 1480.350 1657.880 1480.670 1657.940 ;
        RECT 881.890 58.380 882.210 58.440 ;
        RECT 1477.130 58.380 1477.450 58.440 ;
        RECT 881.890 58.240 1477.450 58.380 ;
        RECT 881.890 58.180 882.210 58.240 ;
        RECT 1477.130 58.180 1477.450 58.240 ;
      LAYER via ;
        RECT 1477.160 1657.880 1477.420 1658.140 ;
        RECT 1480.380 1657.880 1480.640 1658.140 ;
        RECT 881.920 58.180 882.180 58.440 ;
        RECT 1477.160 58.180 1477.420 58.440 ;
      LAYER met2 ;
        RECT 1482.145 1700.410 1482.425 1704.000 ;
        RECT 1480.440 1700.270 1482.425 1700.410 ;
        RECT 1480.440 1658.170 1480.580 1700.270 ;
        RECT 1482.145 1700.000 1482.425 1700.270 ;
        RECT 1477.160 1657.850 1477.420 1658.170 ;
        RECT 1480.380 1657.850 1480.640 1658.170 ;
        RECT 1477.220 58.470 1477.360 1657.850 ;
        RECT 881.920 58.150 882.180 58.470 ;
        RECT 1477.160 58.150 1477.420 58.470 ;
        RECT 881.980 14.010 882.120 58.150 ;
        RECT 881.980 13.870 883.040 14.010 ;
        RECT 882.900 2.400 883.040 13.870 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1484.030 1678.140 1484.350 1678.200 ;
        RECT 1486.790 1678.140 1487.110 1678.200 ;
        RECT 1484.030 1678.000 1487.110 1678.140 ;
        RECT 1484.030 1677.940 1484.350 1678.000 ;
        RECT 1486.790 1677.940 1487.110 1678.000 ;
        RECT 903.510 58.040 903.830 58.100 ;
        RECT 1484.030 58.040 1484.350 58.100 ;
        RECT 903.510 57.900 1484.350 58.040 ;
        RECT 903.510 57.840 903.830 57.900 ;
        RECT 1484.030 57.840 1484.350 57.900 ;
        RECT 900.750 2.960 901.070 3.020 ;
        RECT 903.510 2.960 903.830 3.020 ;
        RECT 900.750 2.820 903.830 2.960 ;
        RECT 900.750 2.760 901.070 2.820 ;
        RECT 903.510 2.760 903.830 2.820 ;
      LAYER via ;
        RECT 1484.060 1677.940 1484.320 1678.200 ;
        RECT 1486.820 1677.940 1487.080 1678.200 ;
        RECT 903.540 57.840 903.800 58.100 ;
        RECT 1484.060 57.840 1484.320 58.100 ;
        RECT 900.780 2.760 901.040 3.020 ;
        RECT 903.540 2.760 903.800 3.020 ;
      LAYER met2 ;
        RECT 1488.585 1700.410 1488.865 1704.000 ;
        RECT 1486.880 1700.270 1488.865 1700.410 ;
        RECT 1486.880 1678.230 1487.020 1700.270 ;
        RECT 1488.585 1700.000 1488.865 1700.270 ;
        RECT 1484.060 1677.910 1484.320 1678.230 ;
        RECT 1486.820 1677.910 1487.080 1678.230 ;
        RECT 1484.120 58.130 1484.260 1677.910 ;
        RECT 903.540 57.810 903.800 58.130 ;
        RECT 1484.060 57.810 1484.320 58.130 ;
        RECT 903.600 3.050 903.740 57.810 ;
        RECT 900.780 2.730 901.040 3.050 ;
        RECT 903.540 2.730 903.800 3.050 ;
        RECT 900.840 2.400 900.980 2.730 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1492.385 1538.925 1492.555 1587.035 ;
        RECT 1492.385 1449.165 1492.555 1497.275 ;
        RECT 1492.385 1352.945 1492.555 1400.715 ;
        RECT 1492.385 1256.385 1492.555 1304.155 ;
        RECT 1492.385 1207.425 1492.555 1255.875 ;
        RECT 1492.385 966.025 1492.555 980.475 ;
        RECT 1492.385 544.085 1492.555 579.615 ;
      LAYER mcon ;
        RECT 1492.385 1586.865 1492.555 1587.035 ;
        RECT 1492.385 1497.105 1492.555 1497.275 ;
        RECT 1492.385 1400.545 1492.555 1400.715 ;
        RECT 1492.385 1303.985 1492.555 1304.155 ;
        RECT 1492.385 1255.705 1492.555 1255.875 ;
        RECT 1492.385 980.305 1492.555 980.475 ;
        RECT 1492.385 579.445 1492.555 579.615 ;
      LAYER met1 ;
        RECT 1492.310 1657.400 1492.630 1657.460 ;
        RECT 1494.610 1657.400 1494.930 1657.460 ;
        RECT 1492.310 1657.260 1494.930 1657.400 ;
        RECT 1492.310 1657.200 1492.630 1657.260 ;
        RECT 1494.610 1657.200 1494.930 1657.260 ;
        RECT 1492.310 1593.820 1492.630 1593.880 ;
        RECT 1492.770 1593.820 1493.090 1593.880 ;
        RECT 1492.310 1593.680 1493.090 1593.820 ;
        RECT 1492.310 1593.620 1492.630 1593.680 ;
        RECT 1492.770 1593.620 1493.090 1593.680 ;
        RECT 1492.310 1587.020 1492.630 1587.080 ;
        RECT 1492.115 1586.880 1492.630 1587.020 ;
        RECT 1492.310 1586.820 1492.630 1586.880 ;
        RECT 1492.310 1539.080 1492.630 1539.140 ;
        RECT 1492.115 1538.940 1492.630 1539.080 ;
        RECT 1492.310 1538.880 1492.630 1538.940 ;
        RECT 1492.325 1497.260 1492.615 1497.305 ;
        RECT 1492.770 1497.260 1493.090 1497.320 ;
        RECT 1492.325 1497.120 1493.090 1497.260 ;
        RECT 1492.325 1497.075 1492.615 1497.120 ;
        RECT 1492.770 1497.060 1493.090 1497.120 ;
        RECT 1492.310 1449.320 1492.630 1449.380 ;
        RECT 1492.115 1449.180 1492.630 1449.320 ;
        RECT 1492.310 1449.120 1492.630 1449.180 ;
        RECT 1492.310 1414.440 1492.630 1414.700 ;
        RECT 1492.400 1413.960 1492.540 1414.440 ;
        RECT 1492.770 1413.960 1493.090 1414.020 ;
        RECT 1492.400 1413.820 1493.090 1413.960 ;
        RECT 1492.770 1413.760 1493.090 1413.820 ;
        RECT 1492.325 1400.700 1492.615 1400.745 ;
        RECT 1492.770 1400.700 1493.090 1400.760 ;
        RECT 1492.325 1400.560 1493.090 1400.700 ;
        RECT 1492.325 1400.515 1492.615 1400.560 ;
        RECT 1492.770 1400.500 1493.090 1400.560 ;
        RECT 1492.310 1353.100 1492.630 1353.160 ;
        RECT 1492.115 1352.960 1492.630 1353.100 ;
        RECT 1492.310 1352.900 1492.630 1352.960 ;
        RECT 1492.310 1317.880 1492.630 1318.140 ;
        RECT 1492.400 1317.400 1492.540 1317.880 ;
        RECT 1492.770 1317.400 1493.090 1317.460 ;
        RECT 1492.400 1317.260 1493.090 1317.400 ;
        RECT 1492.770 1317.200 1493.090 1317.260 ;
        RECT 1492.325 1304.140 1492.615 1304.185 ;
        RECT 1492.770 1304.140 1493.090 1304.200 ;
        RECT 1492.325 1304.000 1493.090 1304.140 ;
        RECT 1492.325 1303.955 1492.615 1304.000 ;
        RECT 1492.770 1303.940 1493.090 1304.000 ;
        RECT 1492.310 1256.540 1492.630 1256.600 ;
        RECT 1492.115 1256.400 1492.630 1256.540 ;
        RECT 1492.310 1256.340 1492.630 1256.400 ;
        RECT 1492.310 1255.860 1492.630 1255.920 ;
        RECT 1492.115 1255.720 1492.630 1255.860 ;
        RECT 1492.310 1255.660 1492.630 1255.720 ;
        RECT 1492.325 1207.580 1492.615 1207.625 ;
        RECT 1492.770 1207.580 1493.090 1207.640 ;
        RECT 1492.325 1207.440 1493.090 1207.580 ;
        RECT 1492.325 1207.395 1492.615 1207.440 ;
        RECT 1492.770 1207.380 1493.090 1207.440 ;
        RECT 1492.770 1159.100 1493.090 1159.360 ;
        RECT 1492.860 1158.680 1493.000 1159.100 ;
        RECT 1492.770 1158.420 1493.090 1158.680 ;
        RECT 1492.770 1145.360 1493.090 1145.420 ;
        RECT 1493.230 1145.360 1493.550 1145.420 ;
        RECT 1492.770 1145.220 1493.550 1145.360 ;
        RECT 1492.770 1145.160 1493.090 1145.220 ;
        RECT 1493.230 1145.160 1493.550 1145.220 ;
        RECT 1492.770 1007.660 1493.090 1007.720 ;
        RECT 1493.230 1007.660 1493.550 1007.720 ;
        RECT 1492.770 1007.520 1493.550 1007.660 ;
        RECT 1492.770 1007.460 1493.090 1007.520 ;
        RECT 1493.230 1007.460 1493.550 1007.520 ;
        RECT 1492.325 980.460 1492.615 980.505 ;
        RECT 1492.770 980.460 1493.090 980.520 ;
        RECT 1492.325 980.320 1493.090 980.460 ;
        RECT 1492.325 980.275 1492.615 980.320 ;
        RECT 1492.770 980.260 1493.090 980.320 ;
        RECT 1492.310 966.180 1492.630 966.240 ;
        RECT 1492.115 966.040 1492.630 966.180 ;
        RECT 1492.310 965.980 1492.630 966.040 ;
        RECT 1492.310 579.600 1492.630 579.660 ;
        RECT 1492.115 579.460 1492.630 579.600 ;
        RECT 1492.310 579.400 1492.630 579.460 ;
        RECT 1492.325 544.240 1492.615 544.285 ;
        RECT 1492.770 544.240 1493.090 544.300 ;
        RECT 1492.325 544.100 1493.090 544.240 ;
        RECT 1492.325 544.055 1492.615 544.100 ;
        RECT 1492.770 544.040 1493.090 544.100 ;
        RECT 1492.770 497.320 1493.090 497.380 ;
        RECT 1492.400 497.180 1493.090 497.320 ;
        RECT 1492.400 496.700 1492.540 497.180 ;
        RECT 1492.770 497.120 1493.090 497.180 ;
        RECT 1492.310 496.440 1492.630 496.700 ;
        RECT 1492.310 434.760 1492.630 434.820 ;
        RECT 1492.770 434.760 1493.090 434.820 ;
        RECT 1492.310 434.620 1493.090 434.760 ;
        RECT 1492.310 434.560 1492.630 434.620 ;
        RECT 1492.770 434.560 1493.090 434.620 ;
        RECT 1492.770 144.740 1493.090 144.800 ;
        RECT 1493.230 144.740 1493.550 144.800 ;
        RECT 1492.770 144.600 1493.550 144.740 ;
        RECT 1492.770 144.540 1493.090 144.600 ;
        RECT 1493.230 144.540 1493.550 144.600 ;
        RECT 923.750 57.700 924.070 57.760 ;
        RECT 1493.230 57.700 1493.550 57.760 ;
        RECT 923.750 57.560 1493.550 57.700 ;
        RECT 923.750 57.500 924.070 57.560 ;
        RECT 1493.230 57.500 1493.550 57.560 ;
        RECT 918.690 2.960 919.010 3.020 ;
        RECT 923.750 2.960 924.070 3.020 ;
        RECT 918.690 2.820 924.070 2.960 ;
        RECT 918.690 2.760 919.010 2.820 ;
        RECT 923.750 2.760 924.070 2.820 ;
      LAYER via ;
        RECT 1492.340 1657.200 1492.600 1657.460 ;
        RECT 1494.640 1657.200 1494.900 1657.460 ;
        RECT 1492.340 1593.620 1492.600 1593.880 ;
        RECT 1492.800 1593.620 1493.060 1593.880 ;
        RECT 1492.340 1586.820 1492.600 1587.080 ;
        RECT 1492.340 1538.880 1492.600 1539.140 ;
        RECT 1492.800 1497.060 1493.060 1497.320 ;
        RECT 1492.340 1449.120 1492.600 1449.380 ;
        RECT 1492.340 1414.440 1492.600 1414.700 ;
        RECT 1492.800 1413.760 1493.060 1414.020 ;
        RECT 1492.800 1400.500 1493.060 1400.760 ;
        RECT 1492.340 1352.900 1492.600 1353.160 ;
        RECT 1492.340 1317.880 1492.600 1318.140 ;
        RECT 1492.800 1317.200 1493.060 1317.460 ;
        RECT 1492.800 1303.940 1493.060 1304.200 ;
        RECT 1492.340 1256.340 1492.600 1256.600 ;
        RECT 1492.340 1255.660 1492.600 1255.920 ;
        RECT 1492.800 1207.380 1493.060 1207.640 ;
        RECT 1492.800 1159.100 1493.060 1159.360 ;
        RECT 1492.800 1158.420 1493.060 1158.680 ;
        RECT 1492.800 1145.160 1493.060 1145.420 ;
        RECT 1493.260 1145.160 1493.520 1145.420 ;
        RECT 1492.800 1007.460 1493.060 1007.720 ;
        RECT 1493.260 1007.460 1493.520 1007.720 ;
        RECT 1492.800 980.260 1493.060 980.520 ;
        RECT 1492.340 965.980 1492.600 966.240 ;
        RECT 1492.340 579.400 1492.600 579.660 ;
        RECT 1492.800 544.040 1493.060 544.300 ;
        RECT 1492.800 497.120 1493.060 497.380 ;
        RECT 1492.340 496.440 1492.600 496.700 ;
        RECT 1492.340 434.560 1492.600 434.820 ;
        RECT 1492.800 434.560 1493.060 434.820 ;
        RECT 1492.800 144.540 1493.060 144.800 ;
        RECT 1493.260 144.540 1493.520 144.800 ;
        RECT 923.780 57.500 924.040 57.760 ;
        RECT 1493.260 57.500 1493.520 57.760 ;
        RECT 918.720 2.760 918.980 3.020 ;
        RECT 923.780 2.760 924.040 3.020 ;
      LAYER met2 ;
        RECT 1495.485 1700.410 1495.765 1704.000 ;
        RECT 1494.700 1700.270 1495.765 1700.410 ;
        RECT 1494.700 1657.490 1494.840 1700.270 ;
        RECT 1495.485 1700.000 1495.765 1700.270 ;
        RECT 1492.340 1657.170 1492.600 1657.490 ;
        RECT 1494.640 1657.170 1494.900 1657.490 ;
        RECT 1492.400 1606.570 1492.540 1657.170 ;
        RECT 1492.400 1606.430 1493.000 1606.570 ;
        RECT 1492.860 1593.910 1493.000 1606.430 ;
        RECT 1492.340 1593.590 1492.600 1593.910 ;
        RECT 1492.800 1593.590 1493.060 1593.910 ;
        RECT 1492.400 1587.110 1492.540 1593.590 ;
        RECT 1492.340 1586.790 1492.600 1587.110 ;
        RECT 1492.340 1538.850 1492.600 1539.170 ;
        RECT 1492.400 1521.570 1492.540 1538.850 ;
        RECT 1491.940 1521.430 1492.540 1521.570 ;
        RECT 1491.940 1510.010 1492.080 1521.430 ;
        RECT 1491.940 1509.870 1493.000 1510.010 ;
        RECT 1492.860 1497.350 1493.000 1509.870 ;
        RECT 1492.800 1497.030 1493.060 1497.350 ;
        RECT 1492.340 1449.090 1492.600 1449.410 ;
        RECT 1492.400 1414.730 1492.540 1449.090 ;
        RECT 1492.340 1414.410 1492.600 1414.730 ;
        RECT 1492.800 1413.730 1493.060 1414.050 ;
        RECT 1492.860 1400.790 1493.000 1413.730 ;
        RECT 1492.800 1400.470 1493.060 1400.790 ;
        RECT 1492.340 1352.870 1492.600 1353.190 ;
        RECT 1492.400 1318.170 1492.540 1352.870 ;
        RECT 1492.340 1317.850 1492.600 1318.170 ;
        RECT 1492.800 1317.170 1493.060 1317.490 ;
        RECT 1492.860 1304.230 1493.000 1317.170 ;
        RECT 1492.800 1303.910 1493.060 1304.230 ;
        RECT 1492.340 1256.310 1492.600 1256.630 ;
        RECT 1492.400 1255.950 1492.540 1256.310 ;
        RECT 1492.340 1255.630 1492.600 1255.950 ;
        RECT 1492.800 1207.350 1493.060 1207.670 ;
        RECT 1492.860 1159.390 1493.000 1207.350 ;
        RECT 1492.800 1159.070 1493.060 1159.390 ;
        RECT 1492.800 1158.390 1493.060 1158.710 ;
        RECT 1492.860 1145.450 1493.000 1158.390 ;
        RECT 1492.800 1145.130 1493.060 1145.450 ;
        RECT 1493.260 1145.130 1493.520 1145.450 ;
        RECT 1493.320 1007.750 1493.460 1145.130 ;
        RECT 1492.800 1007.430 1493.060 1007.750 ;
        RECT 1493.260 1007.430 1493.520 1007.750 ;
        RECT 1492.860 980.550 1493.000 1007.430 ;
        RECT 1492.800 980.230 1493.060 980.550 ;
        RECT 1492.340 965.950 1492.600 966.270 ;
        RECT 1492.400 931.330 1492.540 965.950 ;
        RECT 1492.400 931.190 1493.000 931.330 ;
        RECT 1492.860 786.660 1493.000 931.190 ;
        RECT 1492.400 786.520 1493.000 786.660 ;
        RECT 1492.400 738.210 1492.540 786.520 ;
        RECT 1492.400 738.070 1493.000 738.210 ;
        RECT 1492.860 579.770 1493.000 738.070 ;
        RECT 1492.400 579.690 1493.000 579.770 ;
        RECT 1492.340 579.630 1493.000 579.690 ;
        RECT 1492.340 579.370 1492.600 579.630 ;
        RECT 1492.400 579.215 1492.540 579.370 ;
        RECT 1492.800 544.010 1493.060 544.330 ;
        RECT 1492.860 497.410 1493.000 544.010 ;
        RECT 1492.800 497.090 1493.060 497.410 ;
        RECT 1492.340 496.410 1492.600 496.730 ;
        RECT 1492.400 434.850 1492.540 496.410 ;
        RECT 1492.340 434.530 1492.600 434.850 ;
        RECT 1492.800 434.530 1493.060 434.850 ;
        RECT 1492.860 410.450 1493.000 434.530 ;
        RECT 1492.400 410.310 1493.000 410.450 ;
        RECT 1492.400 303.010 1492.540 410.310 ;
        RECT 1492.400 302.870 1493.000 303.010 ;
        RECT 1492.860 241.810 1493.000 302.870 ;
        RECT 1492.400 241.670 1493.000 241.810 ;
        RECT 1492.400 205.770 1492.540 241.670 ;
        RECT 1492.400 205.630 1493.000 205.770 ;
        RECT 1492.860 144.830 1493.000 205.630 ;
        RECT 1492.800 144.510 1493.060 144.830 ;
        RECT 1493.260 144.510 1493.520 144.830 ;
        RECT 1493.320 57.790 1493.460 144.510 ;
        RECT 923.780 57.470 924.040 57.790 ;
        RECT 1493.260 57.470 1493.520 57.790 ;
        RECT 923.840 3.050 923.980 57.470 ;
        RECT 918.720 2.730 918.980 3.050 ;
        RECT 923.780 2.730 924.040 3.050 ;
        RECT 918.780 2.400 918.920 2.730 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1499.285 241.485 1499.455 255.935 ;
        RECT 1499.285 75.905 1499.455 83.555 ;
      LAYER mcon ;
        RECT 1499.285 255.765 1499.455 255.935 ;
        RECT 1499.285 83.385 1499.455 83.555 ;
      LAYER met1 ;
        RECT 1499.210 1365.820 1499.530 1366.080 ;
        RECT 1499.300 1365.400 1499.440 1365.820 ;
        RECT 1499.210 1365.140 1499.530 1365.400 ;
        RECT 1499.210 1269.260 1499.530 1269.520 ;
        RECT 1499.300 1268.840 1499.440 1269.260 ;
        RECT 1499.210 1268.580 1499.530 1268.840 ;
        RECT 1499.210 1172.700 1499.530 1172.960 ;
        RECT 1499.300 1172.280 1499.440 1172.700 ;
        RECT 1499.210 1172.020 1499.530 1172.280 ;
        RECT 1499.210 1076.140 1499.530 1076.400 ;
        RECT 1499.300 1075.720 1499.440 1076.140 ;
        RECT 1499.210 1075.460 1499.530 1075.720 ;
        RECT 1499.210 979.580 1499.530 979.840 ;
        RECT 1499.300 979.160 1499.440 979.580 ;
        RECT 1499.210 978.900 1499.530 979.160 ;
        RECT 1499.210 869.960 1499.530 870.020 ;
        RECT 1498.840 869.820 1499.530 869.960 ;
        RECT 1498.840 869.680 1498.980 869.820 ;
        RECT 1499.210 869.760 1499.530 869.820 ;
        RECT 1498.750 869.420 1499.070 869.680 ;
        RECT 1498.750 862.480 1499.070 862.540 ;
        RECT 1500.130 862.480 1500.450 862.540 ;
        RECT 1498.750 862.340 1500.450 862.480 ;
        RECT 1498.750 862.280 1499.070 862.340 ;
        RECT 1500.130 862.280 1500.450 862.340 ;
        RECT 1499.210 400.220 1499.530 400.480 ;
        RECT 1499.300 399.800 1499.440 400.220 ;
        RECT 1499.210 399.540 1499.530 399.800 ;
        RECT 1499.210 255.920 1499.530 255.980 ;
        RECT 1499.015 255.780 1499.530 255.920 ;
        RECT 1499.210 255.720 1499.530 255.780 ;
        RECT 1499.210 241.640 1499.530 241.700 ;
        RECT 1499.015 241.500 1499.530 241.640 ;
        RECT 1499.210 241.440 1499.530 241.500 ;
        RECT 1499.210 227.700 1499.530 227.760 ;
        RECT 1499.670 227.700 1499.990 227.760 ;
        RECT 1499.210 227.560 1499.990 227.700 ;
        RECT 1499.210 227.500 1499.530 227.560 ;
        RECT 1499.670 227.500 1499.990 227.560 ;
        RECT 1498.750 179.420 1499.070 179.480 ;
        RECT 1500.130 179.420 1500.450 179.480 ;
        RECT 1498.750 179.280 1500.450 179.420 ;
        RECT 1498.750 179.220 1499.070 179.280 ;
        RECT 1500.130 179.220 1500.450 179.280 ;
        RECT 1499.225 83.540 1499.515 83.585 ;
        RECT 1500.130 83.540 1500.450 83.600 ;
        RECT 1499.225 83.400 1500.450 83.540 ;
        RECT 1499.225 83.355 1499.515 83.400 ;
        RECT 1500.130 83.340 1500.450 83.400 ;
        RECT 1499.210 76.060 1499.530 76.120 ;
        RECT 1499.015 75.920 1499.530 76.060 ;
        RECT 1499.210 75.860 1499.530 75.920 ;
        RECT 938.010 57.360 938.330 57.420 ;
        RECT 1499.210 57.360 1499.530 57.420 ;
        RECT 938.010 57.220 1499.530 57.360 ;
        RECT 938.010 57.160 938.330 57.220 ;
        RECT 1499.210 57.160 1499.530 57.220 ;
      LAYER via ;
        RECT 1499.240 1365.820 1499.500 1366.080 ;
        RECT 1499.240 1365.140 1499.500 1365.400 ;
        RECT 1499.240 1269.260 1499.500 1269.520 ;
        RECT 1499.240 1268.580 1499.500 1268.840 ;
        RECT 1499.240 1172.700 1499.500 1172.960 ;
        RECT 1499.240 1172.020 1499.500 1172.280 ;
        RECT 1499.240 1076.140 1499.500 1076.400 ;
        RECT 1499.240 1075.460 1499.500 1075.720 ;
        RECT 1499.240 979.580 1499.500 979.840 ;
        RECT 1499.240 978.900 1499.500 979.160 ;
        RECT 1499.240 869.760 1499.500 870.020 ;
        RECT 1498.780 869.420 1499.040 869.680 ;
        RECT 1498.780 862.280 1499.040 862.540 ;
        RECT 1500.160 862.280 1500.420 862.540 ;
        RECT 1499.240 400.220 1499.500 400.480 ;
        RECT 1499.240 399.540 1499.500 399.800 ;
        RECT 1499.240 255.720 1499.500 255.980 ;
        RECT 1499.240 241.440 1499.500 241.700 ;
        RECT 1499.240 227.500 1499.500 227.760 ;
        RECT 1499.700 227.500 1499.960 227.760 ;
        RECT 1498.780 179.220 1499.040 179.480 ;
        RECT 1500.160 179.220 1500.420 179.480 ;
        RECT 1500.160 83.340 1500.420 83.600 ;
        RECT 1499.240 75.860 1499.500 76.120 ;
        RECT 938.040 57.160 938.300 57.420 ;
        RECT 1499.240 57.160 1499.500 57.420 ;
      LAYER met2 ;
        RECT 1502.385 1700.410 1502.665 1704.000 ;
        RECT 1501.140 1700.270 1502.665 1700.410 ;
        RECT 1501.140 1656.210 1501.280 1700.270 ;
        RECT 1502.385 1700.000 1502.665 1700.270 ;
        RECT 1499.300 1656.070 1501.280 1656.210 ;
        RECT 1499.300 1559.650 1499.440 1656.070 ;
        RECT 1498.840 1559.510 1499.440 1559.650 ;
        RECT 1498.840 1558.970 1498.980 1559.510 ;
        RECT 1498.840 1558.830 1499.440 1558.970 ;
        RECT 1499.300 1463.090 1499.440 1558.830 ;
        RECT 1498.840 1462.950 1499.440 1463.090 ;
        RECT 1498.840 1462.410 1498.980 1462.950 ;
        RECT 1498.840 1462.270 1499.440 1462.410 ;
        RECT 1499.300 1366.110 1499.440 1462.270 ;
        RECT 1499.240 1365.790 1499.500 1366.110 ;
        RECT 1499.240 1365.110 1499.500 1365.430 ;
        RECT 1499.300 1269.550 1499.440 1365.110 ;
        RECT 1499.240 1269.230 1499.500 1269.550 ;
        RECT 1499.240 1268.550 1499.500 1268.870 ;
        RECT 1499.300 1172.990 1499.440 1268.550 ;
        RECT 1499.240 1172.670 1499.500 1172.990 ;
        RECT 1499.240 1171.990 1499.500 1172.310 ;
        RECT 1499.300 1076.430 1499.440 1171.990 ;
        RECT 1499.240 1076.110 1499.500 1076.430 ;
        RECT 1499.240 1075.430 1499.500 1075.750 ;
        RECT 1499.300 979.870 1499.440 1075.430 ;
        RECT 1499.240 979.550 1499.500 979.870 ;
        RECT 1499.240 978.870 1499.500 979.190 ;
        RECT 1499.300 870.050 1499.440 978.870 ;
        RECT 1499.240 869.730 1499.500 870.050 ;
        RECT 1498.780 869.390 1499.040 869.710 ;
        RECT 1498.840 862.570 1498.980 869.390 ;
        RECT 1498.780 862.250 1499.040 862.570 ;
        RECT 1500.160 862.250 1500.420 862.570 ;
        RECT 1500.220 785.130 1500.360 862.250 ;
        RECT 1499.300 784.990 1500.360 785.130 ;
        RECT 1499.300 594.050 1499.440 784.990 ;
        RECT 1498.840 593.910 1499.440 594.050 ;
        RECT 1498.840 593.370 1498.980 593.910 ;
        RECT 1498.840 593.230 1499.440 593.370 ;
        RECT 1499.300 400.510 1499.440 593.230 ;
        RECT 1499.240 400.190 1499.500 400.510 ;
        RECT 1499.240 399.510 1499.500 399.830 ;
        RECT 1499.300 256.010 1499.440 399.510 ;
        RECT 1499.240 255.690 1499.500 256.010 ;
        RECT 1499.240 241.410 1499.500 241.730 ;
        RECT 1499.300 227.790 1499.440 241.410 ;
        RECT 1499.240 227.470 1499.500 227.790 ;
        RECT 1499.700 227.470 1499.960 227.790 ;
        RECT 1499.760 180.045 1499.900 227.470 ;
        RECT 1498.770 179.675 1499.050 180.045 ;
        RECT 1499.690 179.675 1499.970 180.045 ;
        RECT 1498.840 179.510 1498.980 179.675 ;
        RECT 1498.780 179.190 1499.040 179.510 ;
        RECT 1500.160 179.190 1500.420 179.510 ;
        RECT 1500.220 83.630 1500.360 179.190 ;
        RECT 1500.160 83.310 1500.420 83.630 ;
        RECT 1499.240 75.830 1499.500 76.150 ;
        RECT 1499.300 57.450 1499.440 75.830 ;
        RECT 938.040 57.130 938.300 57.450 ;
        RECT 1499.240 57.130 1499.500 57.450 ;
        RECT 938.100 3.130 938.240 57.130 ;
        RECT 936.720 2.990 938.240 3.130 ;
        RECT 936.720 2.960 936.860 2.990 ;
        RECT 936.260 2.820 936.860 2.960 ;
        RECT 936.260 2.400 936.400 2.820 ;
        RECT 936.050 -4.800 936.610 2.400 ;
      LAYER via2 ;
        RECT 1498.770 179.720 1499.050 180.000 ;
        RECT 1499.690 179.720 1499.970 180.000 ;
      LAYER met3 ;
        RECT 1498.745 180.010 1499.075 180.025 ;
        RECT 1499.665 180.010 1499.995 180.025 ;
        RECT 1498.745 179.710 1499.995 180.010 ;
        RECT 1498.745 179.695 1499.075 179.710 ;
        RECT 1499.665 179.695 1499.995 179.710 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1504.730 1664.200 1505.050 1664.260 ;
        RECT 1507.030 1664.200 1507.350 1664.260 ;
        RECT 1504.730 1664.060 1507.350 1664.200 ;
        RECT 1504.730 1664.000 1505.050 1664.060 ;
        RECT 1507.030 1664.000 1507.350 1664.060 ;
        RECT 958.710 57.020 959.030 57.080 ;
        RECT 1504.730 57.020 1505.050 57.080 ;
        RECT 958.710 56.880 1505.050 57.020 ;
        RECT 958.710 56.820 959.030 56.880 ;
        RECT 1504.730 56.820 1505.050 56.880 ;
        RECT 954.110 2.960 954.430 3.020 ;
        RECT 958.710 2.960 959.030 3.020 ;
        RECT 954.110 2.820 959.030 2.960 ;
        RECT 954.110 2.760 954.430 2.820 ;
        RECT 958.710 2.760 959.030 2.820 ;
      LAYER via ;
        RECT 1504.760 1664.000 1505.020 1664.260 ;
        RECT 1507.060 1664.000 1507.320 1664.260 ;
        RECT 958.740 56.820 959.000 57.080 ;
        RECT 1504.760 56.820 1505.020 57.080 ;
        RECT 954.140 2.760 954.400 3.020 ;
        RECT 958.740 2.760 959.000 3.020 ;
      LAYER met2 ;
        RECT 1508.825 1700.410 1509.105 1704.000 ;
        RECT 1507.120 1700.270 1509.105 1700.410 ;
        RECT 1507.120 1664.290 1507.260 1700.270 ;
        RECT 1508.825 1700.000 1509.105 1700.270 ;
        RECT 1504.760 1663.970 1505.020 1664.290 ;
        RECT 1507.060 1663.970 1507.320 1664.290 ;
        RECT 1504.820 57.110 1504.960 1663.970 ;
        RECT 958.740 56.790 959.000 57.110 ;
        RECT 1504.760 56.790 1505.020 57.110 ;
        RECT 958.800 3.050 958.940 56.790 ;
        RECT 954.140 2.730 954.400 3.050 ;
        RECT 958.740 2.730 959.000 3.050 ;
        RECT 954.200 2.400 954.340 2.730 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1511.630 1678.140 1511.950 1678.200 ;
        RECT 1514.390 1678.140 1514.710 1678.200 ;
        RECT 1511.630 1678.000 1514.710 1678.140 ;
        RECT 1511.630 1677.940 1511.950 1678.000 ;
        RECT 1514.390 1677.940 1514.710 1678.000 ;
        RECT 972.050 56.680 972.370 56.740 ;
        RECT 1511.630 56.680 1511.950 56.740 ;
        RECT 972.050 56.540 1511.950 56.680 ;
        RECT 972.050 56.480 972.370 56.540 ;
        RECT 1511.630 56.480 1511.950 56.540 ;
      LAYER via ;
        RECT 1511.660 1677.940 1511.920 1678.200 ;
        RECT 1514.420 1677.940 1514.680 1678.200 ;
        RECT 972.080 56.480 972.340 56.740 ;
        RECT 1511.660 56.480 1511.920 56.740 ;
      LAYER met2 ;
        RECT 1515.725 1700.410 1516.005 1704.000 ;
        RECT 1514.480 1700.270 1516.005 1700.410 ;
        RECT 1514.480 1678.230 1514.620 1700.270 ;
        RECT 1515.725 1700.000 1516.005 1700.270 ;
        RECT 1511.660 1677.910 1511.920 1678.230 ;
        RECT 1514.420 1677.910 1514.680 1678.230 ;
        RECT 1511.720 56.770 1511.860 1677.910 ;
        RECT 972.080 56.450 972.340 56.770 ;
        RECT 1511.660 56.450 1511.920 56.770 ;
        RECT 972.140 2.400 972.280 56.450 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 26.760 651.290 26.820 ;
        RECT 1393.870 26.760 1394.190 26.820 ;
        RECT 650.970 26.620 1394.190 26.760 ;
        RECT 650.970 26.560 651.290 26.620 ;
        RECT 1393.870 26.560 1394.190 26.620 ;
      LAYER via ;
        RECT 651.000 26.560 651.260 26.820 ;
        RECT 1393.900 26.560 1394.160 26.820 ;
      LAYER met2 ;
        RECT 1394.285 1700.410 1394.565 1704.000 ;
        RECT 1393.960 1700.270 1394.565 1700.410 ;
        RECT 1393.960 26.850 1394.100 1700.270 ;
        RECT 1394.285 1700.000 1394.565 1700.270 ;
        RECT 651.000 26.530 651.260 26.850 ;
        RECT 1393.900 26.530 1394.160 26.850 ;
        RECT 651.060 2.400 651.200 26.530 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1518.990 1678.140 1519.310 1678.200 ;
        RECT 1520.830 1678.140 1521.150 1678.200 ;
        RECT 1518.990 1678.000 1521.150 1678.140 ;
        RECT 1518.990 1677.940 1519.310 1678.000 ;
        RECT 1520.830 1677.940 1521.150 1678.000 ;
        RECT 993.210 56.340 993.530 56.400 ;
        RECT 1518.990 56.340 1519.310 56.400 ;
        RECT 993.210 56.200 1519.310 56.340 ;
        RECT 993.210 56.140 993.530 56.200 ;
        RECT 1518.990 56.140 1519.310 56.200 ;
        RECT 989.990 2.960 990.310 3.020 ;
        RECT 993.210 2.960 993.530 3.020 ;
        RECT 989.990 2.820 993.530 2.960 ;
        RECT 989.990 2.760 990.310 2.820 ;
        RECT 993.210 2.760 993.530 2.820 ;
      LAYER via ;
        RECT 1519.020 1677.940 1519.280 1678.200 ;
        RECT 1520.860 1677.940 1521.120 1678.200 ;
        RECT 993.240 56.140 993.500 56.400 ;
        RECT 1519.020 56.140 1519.280 56.400 ;
        RECT 990.020 2.760 990.280 3.020 ;
        RECT 993.240 2.760 993.500 3.020 ;
      LAYER met2 ;
        RECT 1522.625 1700.410 1522.905 1704.000 ;
        RECT 1520.920 1700.270 1522.905 1700.410 ;
        RECT 1520.920 1678.230 1521.060 1700.270 ;
        RECT 1522.625 1700.000 1522.905 1700.270 ;
        RECT 1519.020 1677.910 1519.280 1678.230 ;
        RECT 1520.860 1677.910 1521.120 1678.230 ;
        RECT 1519.080 56.430 1519.220 1677.910 ;
        RECT 993.240 56.110 993.500 56.430 ;
        RECT 1519.020 56.110 1519.280 56.430 ;
        RECT 993.300 3.050 993.440 56.110 ;
        RECT 990.020 2.730 990.280 3.050 ;
        RECT 993.240 2.730 993.500 3.050 ;
        RECT 990.080 2.400 990.220 2.730 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1335.065 1642.285 1335.235 1686.315 ;
        RECT 1496.985 1685.125 1497.155 1686.315 ;
        RECT 1497.445 1685.125 1497.615 1686.315 ;
        RECT 1335.065 1497.445 1335.235 1545.215 ;
        RECT 1335.065 1062.585 1335.235 1076.695 ;
        RECT 1335.065 1013.965 1335.235 1055.615 ;
        RECT 1335.065 952.425 1335.235 1000.535 ;
        RECT 1335.525 641.325 1335.695 676.175 ;
        RECT 1335.065 414.205 1335.235 510.595 ;
        RECT 1335.525 338.045 1335.695 389.895 ;
        RECT 1335.065 282.965 1335.235 305.575 ;
        RECT 1335.525 193.205 1335.695 241.315 ;
        RECT 1335.065 138.125 1335.235 186.235 ;
      LAYER mcon ;
        RECT 1335.065 1686.145 1335.235 1686.315 ;
        RECT 1496.985 1686.145 1497.155 1686.315 ;
        RECT 1497.445 1686.145 1497.615 1686.315 ;
        RECT 1335.065 1545.045 1335.235 1545.215 ;
        RECT 1335.065 1076.525 1335.235 1076.695 ;
        RECT 1335.065 1055.445 1335.235 1055.615 ;
        RECT 1335.065 1000.365 1335.235 1000.535 ;
        RECT 1335.525 676.005 1335.695 676.175 ;
        RECT 1335.065 510.425 1335.235 510.595 ;
        RECT 1335.525 389.725 1335.695 389.895 ;
        RECT 1335.065 305.405 1335.235 305.575 ;
        RECT 1335.525 241.145 1335.695 241.315 ;
        RECT 1335.065 186.065 1335.235 186.235 ;
      LAYER met1 ;
        RECT 1335.005 1686.300 1335.295 1686.345 ;
        RECT 1496.925 1686.300 1497.215 1686.345 ;
        RECT 1335.005 1686.160 1497.215 1686.300 ;
        RECT 1335.005 1686.115 1335.295 1686.160 ;
        RECT 1496.925 1686.115 1497.215 1686.160 ;
        RECT 1497.385 1686.300 1497.675 1686.345 ;
        RECT 1529.110 1686.300 1529.430 1686.360 ;
        RECT 1497.385 1686.160 1529.430 1686.300 ;
        RECT 1497.385 1686.115 1497.675 1686.160 ;
        RECT 1529.110 1686.100 1529.430 1686.160 ;
        RECT 1496.925 1685.280 1497.215 1685.325 ;
        RECT 1497.385 1685.280 1497.675 1685.325 ;
        RECT 1496.925 1685.140 1497.675 1685.280 ;
        RECT 1496.925 1685.095 1497.215 1685.140 ;
        RECT 1497.385 1685.095 1497.675 1685.140 ;
        RECT 1334.990 1642.440 1335.310 1642.500 ;
        RECT 1334.795 1642.300 1335.310 1642.440 ;
        RECT 1334.990 1642.240 1335.310 1642.300 ;
        RECT 1335.450 1608.100 1335.770 1608.160 ;
        RECT 1335.080 1607.960 1335.770 1608.100 ;
        RECT 1335.080 1607.140 1335.220 1607.960 ;
        RECT 1335.450 1607.900 1335.770 1607.960 ;
        RECT 1334.990 1606.880 1335.310 1607.140 ;
        RECT 1334.530 1545.880 1334.850 1545.940 ;
        RECT 1334.990 1545.880 1335.310 1545.940 ;
        RECT 1334.530 1545.740 1335.310 1545.880 ;
        RECT 1334.530 1545.680 1334.850 1545.740 ;
        RECT 1334.990 1545.680 1335.310 1545.740 ;
        RECT 1334.990 1545.200 1335.310 1545.260 ;
        RECT 1334.795 1545.060 1335.310 1545.200 ;
        RECT 1334.990 1545.000 1335.310 1545.060 ;
        RECT 1335.005 1497.600 1335.295 1497.645 ;
        RECT 1336.370 1497.600 1336.690 1497.660 ;
        RECT 1335.005 1497.460 1336.690 1497.600 ;
        RECT 1335.005 1497.415 1335.295 1497.460 ;
        RECT 1336.370 1497.400 1336.690 1497.460 ;
        RECT 1334.990 1462.920 1335.310 1462.980 ;
        RECT 1336.370 1462.920 1336.690 1462.980 ;
        RECT 1334.990 1462.780 1336.690 1462.920 ;
        RECT 1334.990 1462.720 1335.310 1462.780 ;
        RECT 1336.370 1462.720 1336.690 1462.780 ;
        RECT 1334.990 1448.980 1335.310 1449.040 ;
        RECT 1336.370 1448.980 1336.690 1449.040 ;
        RECT 1334.990 1448.840 1336.690 1448.980 ;
        RECT 1334.990 1448.780 1335.310 1448.840 ;
        RECT 1336.370 1448.780 1336.690 1448.840 ;
        RECT 1335.910 1297.340 1336.230 1297.400 ;
        RECT 1336.370 1297.340 1336.690 1297.400 ;
        RECT 1335.910 1297.200 1336.690 1297.340 ;
        RECT 1335.910 1297.140 1336.230 1297.200 ;
        RECT 1336.370 1297.140 1336.690 1297.200 ;
        RECT 1334.990 1249.060 1335.310 1249.120 ;
        RECT 1336.370 1249.060 1336.690 1249.120 ;
        RECT 1334.990 1248.920 1336.690 1249.060 ;
        RECT 1334.990 1248.860 1335.310 1248.920 ;
        RECT 1336.370 1248.860 1336.690 1248.920 ;
        RECT 1334.990 1207.380 1335.310 1207.640 ;
        RECT 1335.080 1206.960 1335.220 1207.380 ;
        RECT 1334.990 1206.700 1335.310 1206.960 ;
        RECT 1334.070 1152.500 1334.390 1152.560 ;
        RECT 1334.990 1152.500 1335.310 1152.560 ;
        RECT 1334.070 1152.360 1335.310 1152.500 ;
        RECT 1334.070 1152.300 1334.390 1152.360 ;
        RECT 1334.990 1152.300 1335.310 1152.360 ;
        RECT 1334.530 1104.220 1334.850 1104.280 ;
        RECT 1334.990 1104.220 1335.310 1104.280 ;
        RECT 1334.530 1104.080 1335.310 1104.220 ;
        RECT 1334.530 1104.020 1334.850 1104.080 ;
        RECT 1334.990 1104.020 1335.310 1104.080 ;
        RECT 1334.990 1076.680 1335.310 1076.740 ;
        RECT 1334.795 1076.540 1335.310 1076.680 ;
        RECT 1334.990 1076.480 1335.310 1076.540 ;
        RECT 1334.990 1062.740 1335.310 1062.800 ;
        RECT 1334.795 1062.600 1335.310 1062.740 ;
        RECT 1334.990 1062.540 1335.310 1062.600 ;
        RECT 1334.990 1055.600 1335.310 1055.660 ;
        RECT 1334.795 1055.460 1335.310 1055.600 ;
        RECT 1334.990 1055.400 1335.310 1055.460 ;
        RECT 1335.005 1014.120 1335.295 1014.165 ;
        RECT 1335.450 1014.120 1335.770 1014.180 ;
        RECT 1335.005 1013.980 1335.770 1014.120 ;
        RECT 1335.005 1013.935 1335.295 1013.980 ;
        RECT 1335.450 1013.920 1335.770 1013.980 ;
        RECT 1335.005 1000.520 1335.295 1000.565 ;
        RECT 1335.450 1000.520 1335.770 1000.580 ;
        RECT 1335.005 1000.380 1335.770 1000.520 ;
        RECT 1335.005 1000.335 1335.295 1000.380 ;
        RECT 1335.450 1000.320 1335.770 1000.380 ;
        RECT 1334.990 952.580 1335.310 952.640 ;
        RECT 1334.795 952.440 1335.310 952.580 ;
        RECT 1334.990 952.380 1335.310 952.440 ;
        RECT 1335.450 869.960 1335.770 870.020 ;
        RECT 1335.080 869.820 1335.770 869.960 ;
        RECT 1335.080 869.680 1335.220 869.820 ;
        RECT 1335.450 869.760 1335.770 869.820 ;
        RECT 1334.990 869.420 1335.310 869.680 ;
        RECT 1335.910 690.440 1336.230 690.500 ;
        RECT 1335.540 690.300 1336.230 690.440 ;
        RECT 1335.540 689.820 1335.680 690.300 ;
        RECT 1335.910 690.240 1336.230 690.300 ;
        RECT 1335.450 689.560 1335.770 689.820 ;
        RECT 1335.450 676.160 1335.770 676.220 ;
        RECT 1335.255 676.020 1335.770 676.160 ;
        RECT 1335.450 675.960 1335.770 676.020 ;
        RECT 1335.450 641.480 1335.770 641.540 ;
        RECT 1335.255 641.340 1335.770 641.480 ;
        RECT 1335.450 641.280 1335.770 641.340 ;
        RECT 1334.990 593.540 1335.310 593.600 ;
        RECT 1335.910 593.540 1336.230 593.600 ;
        RECT 1334.990 593.400 1336.230 593.540 ;
        RECT 1334.990 593.340 1335.310 593.400 ;
        RECT 1335.910 593.340 1336.230 593.400 ;
        RECT 1334.990 579.600 1335.310 579.660 ;
        RECT 1335.910 579.600 1336.230 579.660 ;
        RECT 1334.990 579.460 1336.230 579.600 ;
        RECT 1334.990 579.400 1335.310 579.460 ;
        RECT 1335.910 579.400 1336.230 579.460 ;
        RECT 1335.005 510.580 1335.295 510.625 ;
        RECT 1335.450 510.580 1335.770 510.640 ;
        RECT 1335.005 510.440 1335.770 510.580 ;
        RECT 1335.005 510.395 1335.295 510.440 ;
        RECT 1335.450 510.380 1335.770 510.440 ;
        RECT 1335.005 414.360 1335.295 414.405 ;
        RECT 1335.450 414.360 1335.770 414.420 ;
        RECT 1335.005 414.220 1335.770 414.360 ;
        RECT 1335.005 414.175 1335.295 414.220 ;
        RECT 1335.450 414.160 1335.770 414.220 ;
        RECT 1335.450 389.880 1335.770 389.940 ;
        RECT 1335.255 389.740 1335.770 389.880 ;
        RECT 1335.450 389.680 1335.770 389.740 ;
        RECT 1335.450 338.200 1335.770 338.260 ;
        RECT 1335.255 338.060 1335.770 338.200 ;
        RECT 1335.450 338.000 1335.770 338.060 ;
        RECT 1335.005 305.560 1335.295 305.605 ;
        RECT 1335.450 305.560 1335.770 305.620 ;
        RECT 1335.005 305.420 1335.770 305.560 ;
        RECT 1335.005 305.375 1335.295 305.420 ;
        RECT 1335.450 305.360 1335.770 305.420 ;
        RECT 1334.990 283.120 1335.310 283.180 ;
        RECT 1334.795 282.980 1335.310 283.120 ;
        RECT 1334.990 282.920 1335.310 282.980 ;
        RECT 1335.465 241.300 1335.755 241.345 ;
        RECT 1335.910 241.300 1336.230 241.360 ;
        RECT 1335.465 241.160 1336.230 241.300 ;
        RECT 1335.465 241.115 1335.755 241.160 ;
        RECT 1335.910 241.100 1336.230 241.160 ;
        RECT 1335.450 193.360 1335.770 193.420 ;
        RECT 1335.255 193.220 1335.770 193.360 ;
        RECT 1335.450 193.160 1335.770 193.220 ;
        RECT 1335.005 186.220 1335.295 186.265 ;
        RECT 1335.450 186.220 1335.770 186.280 ;
        RECT 1335.005 186.080 1335.770 186.220 ;
        RECT 1335.005 186.035 1335.295 186.080 ;
        RECT 1335.450 186.020 1335.770 186.080 ;
        RECT 1334.990 138.280 1335.310 138.340 ;
        RECT 1334.795 138.140 1335.310 138.280 ;
        RECT 1334.990 138.080 1335.310 138.140 ;
        RECT 1007.470 21.660 1007.790 21.720 ;
        RECT 1336.370 21.660 1336.690 21.720 ;
        RECT 1007.470 21.520 1336.690 21.660 ;
        RECT 1007.470 21.460 1007.790 21.520 ;
        RECT 1336.370 21.460 1336.690 21.520 ;
      LAYER via ;
        RECT 1529.140 1686.100 1529.400 1686.360 ;
        RECT 1335.020 1642.240 1335.280 1642.500 ;
        RECT 1335.480 1607.900 1335.740 1608.160 ;
        RECT 1335.020 1606.880 1335.280 1607.140 ;
        RECT 1334.560 1545.680 1334.820 1545.940 ;
        RECT 1335.020 1545.680 1335.280 1545.940 ;
        RECT 1335.020 1545.000 1335.280 1545.260 ;
        RECT 1336.400 1497.400 1336.660 1497.660 ;
        RECT 1335.020 1462.720 1335.280 1462.980 ;
        RECT 1336.400 1462.720 1336.660 1462.980 ;
        RECT 1335.020 1448.780 1335.280 1449.040 ;
        RECT 1336.400 1448.780 1336.660 1449.040 ;
        RECT 1335.940 1297.140 1336.200 1297.400 ;
        RECT 1336.400 1297.140 1336.660 1297.400 ;
        RECT 1335.020 1248.860 1335.280 1249.120 ;
        RECT 1336.400 1248.860 1336.660 1249.120 ;
        RECT 1335.020 1207.380 1335.280 1207.640 ;
        RECT 1335.020 1206.700 1335.280 1206.960 ;
        RECT 1334.100 1152.300 1334.360 1152.560 ;
        RECT 1335.020 1152.300 1335.280 1152.560 ;
        RECT 1334.560 1104.020 1334.820 1104.280 ;
        RECT 1335.020 1104.020 1335.280 1104.280 ;
        RECT 1335.020 1076.480 1335.280 1076.740 ;
        RECT 1335.020 1062.540 1335.280 1062.800 ;
        RECT 1335.020 1055.400 1335.280 1055.660 ;
        RECT 1335.480 1013.920 1335.740 1014.180 ;
        RECT 1335.480 1000.320 1335.740 1000.580 ;
        RECT 1335.020 952.380 1335.280 952.640 ;
        RECT 1335.480 869.760 1335.740 870.020 ;
        RECT 1335.020 869.420 1335.280 869.680 ;
        RECT 1335.940 690.240 1336.200 690.500 ;
        RECT 1335.480 689.560 1335.740 689.820 ;
        RECT 1335.480 675.960 1335.740 676.220 ;
        RECT 1335.480 641.280 1335.740 641.540 ;
        RECT 1335.020 593.340 1335.280 593.600 ;
        RECT 1335.940 593.340 1336.200 593.600 ;
        RECT 1335.020 579.400 1335.280 579.660 ;
        RECT 1335.940 579.400 1336.200 579.660 ;
        RECT 1335.480 510.380 1335.740 510.640 ;
        RECT 1335.480 414.160 1335.740 414.420 ;
        RECT 1335.480 389.680 1335.740 389.940 ;
        RECT 1335.480 338.000 1335.740 338.260 ;
        RECT 1335.480 305.360 1335.740 305.620 ;
        RECT 1335.020 282.920 1335.280 283.180 ;
        RECT 1335.940 241.100 1336.200 241.360 ;
        RECT 1335.480 193.160 1335.740 193.420 ;
        RECT 1335.480 186.020 1335.740 186.280 ;
        RECT 1335.020 138.080 1335.280 138.340 ;
        RECT 1007.500 21.460 1007.760 21.720 ;
        RECT 1336.400 21.460 1336.660 21.720 ;
      LAYER met2 ;
        RECT 1529.065 1700.000 1529.345 1704.000 ;
        RECT 1529.200 1686.390 1529.340 1700.000 ;
        RECT 1529.140 1686.070 1529.400 1686.390 ;
        RECT 1335.020 1642.210 1335.280 1642.530 ;
        RECT 1335.080 1641.930 1335.220 1642.210 ;
        RECT 1335.080 1641.790 1335.680 1641.930 ;
        RECT 1335.540 1608.190 1335.680 1641.790 ;
        RECT 1335.480 1607.870 1335.740 1608.190 ;
        RECT 1335.020 1606.850 1335.280 1607.170 ;
        RECT 1335.080 1559.650 1335.220 1606.850 ;
        RECT 1334.620 1559.510 1335.220 1559.650 ;
        RECT 1334.620 1545.970 1334.760 1559.510 ;
        RECT 1334.560 1545.650 1334.820 1545.970 ;
        RECT 1335.020 1545.650 1335.280 1545.970 ;
        RECT 1335.080 1545.290 1335.220 1545.650 ;
        RECT 1335.020 1544.970 1335.280 1545.290 ;
        RECT 1336.400 1497.370 1336.660 1497.690 ;
        RECT 1336.460 1463.010 1336.600 1497.370 ;
        RECT 1335.020 1462.690 1335.280 1463.010 ;
        RECT 1336.400 1462.690 1336.660 1463.010 ;
        RECT 1335.080 1449.070 1335.220 1462.690 ;
        RECT 1335.020 1448.750 1335.280 1449.070 ;
        RECT 1336.400 1448.750 1336.660 1449.070 ;
        RECT 1336.460 1353.725 1336.600 1448.750 ;
        RECT 1336.390 1353.355 1336.670 1353.725 ;
        RECT 1335.010 1352.675 1335.290 1353.045 ;
        RECT 1335.080 1345.565 1335.220 1352.675 ;
        RECT 1335.010 1345.195 1335.290 1345.565 ;
        RECT 1335.930 1345.195 1336.210 1345.565 ;
        RECT 1336.000 1297.430 1336.140 1345.195 ;
        RECT 1335.940 1297.110 1336.200 1297.430 ;
        RECT 1336.400 1297.110 1336.660 1297.430 ;
        RECT 1336.460 1249.150 1336.600 1297.110 ;
        RECT 1335.020 1248.830 1335.280 1249.150 ;
        RECT 1336.400 1248.830 1336.660 1249.150 ;
        RECT 1335.080 1207.670 1335.220 1248.830 ;
        RECT 1335.020 1207.350 1335.280 1207.670 ;
        RECT 1335.020 1206.670 1335.280 1206.990 ;
        RECT 1335.080 1152.590 1335.220 1206.670 ;
        RECT 1334.100 1152.330 1334.360 1152.590 ;
        RECT 1334.100 1152.270 1334.760 1152.330 ;
        RECT 1335.020 1152.270 1335.280 1152.590 ;
        RECT 1334.160 1152.190 1334.760 1152.270 ;
        RECT 1334.620 1104.310 1334.760 1152.190 ;
        RECT 1334.560 1103.990 1334.820 1104.310 ;
        RECT 1335.020 1103.990 1335.280 1104.310 ;
        RECT 1335.080 1076.770 1335.220 1103.990 ;
        RECT 1335.020 1076.450 1335.280 1076.770 ;
        RECT 1335.020 1062.510 1335.280 1062.830 ;
        RECT 1335.080 1055.690 1335.220 1062.510 ;
        RECT 1335.020 1055.370 1335.280 1055.690 ;
        RECT 1335.480 1013.890 1335.740 1014.210 ;
        RECT 1335.540 1000.610 1335.680 1013.890 ;
        RECT 1335.480 1000.290 1335.740 1000.610 ;
        RECT 1335.020 952.350 1335.280 952.670 ;
        RECT 1335.080 934.730 1335.220 952.350 ;
        RECT 1335.080 934.590 1335.680 934.730 ;
        RECT 1335.540 870.050 1335.680 934.590 ;
        RECT 1335.480 869.730 1335.740 870.050 ;
        RECT 1335.020 869.390 1335.280 869.710 ;
        RECT 1335.080 821.285 1335.220 869.390 ;
        RECT 1335.010 820.915 1335.290 821.285 ;
        RECT 1336.390 820.235 1336.670 820.605 ;
        RECT 1336.460 773.005 1336.600 820.235 ;
        RECT 1335.010 772.635 1335.290 773.005 ;
        RECT 1336.390 772.635 1336.670 773.005 ;
        RECT 1335.080 738.210 1335.220 772.635 ;
        RECT 1335.080 738.070 1336.140 738.210 ;
        RECT 1336.000 690.530 1336.140 738.070 ;
        RECT 1335.940 690.210 1336.200 690.530 ;
        RECT 1335.480 689.530 1335.740 689.850 ;
        RECT 1335.540 676.250 1335.680 689.530 ;
        RECT 1335.480 675.930 1335.740 676.250 ;
        RECT 1335.480 641.250 1335.740 641.570 ;
        RECT 1335.540 628.050 1335.680 641.250 ;
        RECT 1335.540 627.910 1336.140 628.050 ;
        RECT 1336.000 593.630 1336.140 627.910 ;
        RECT 1335.020 593.310 1335.280 593.630 ;
        RECT 1335.940 593.310 1336.200 593.630 ;
        RECT 1335.080 579.690 1335.220 593.310 ;
        RECT 1335.020 579.370 1335.280 579.690 ;
        RECT 1335.940 579.370 1336.200 579.690 ;
        RECT 1336.000 543.730 1336.140 579.370 ;
        RECT 1335.540 543.590 1336.140 543.730 ;
        RECT 1335.540 510.670 1335.680 543.590 ;
        RECT 1335.480 510.350 1335.740 510.670 ;
        RECT 1335.480 414.130 1335.740 414.450 ;
        RECT 1335.540 389.970 1335.680 414.130 ;
        RECT 1335.480 389.650 1335.740 389.970 ;
        RECT 1335.480 337.970 1335.740 338.290 ;
        RECT 1335.540 305.650 1335.680 337.970 ;
        RECT 1335.480 305.330 1335.740 305.650 ;
        RECT 1335.020 282.890 1335.280 283.210 ;
        RECT 1335.080 280.570 1335.220 282.890 ;
        RECT 1335.080 280.430 1336.140 280.570 ;
        RECT 1336.000 241.390 1336.140 280.430 ;
        RECT 1335.940 241.070 1336.200 241.390 ;
        RECT 1335.480 193.130 1335.740 193.450 ;
        RECT 1335.540 186.310 1335.680 193.130 ;
        RECT 1335.480 185.990 1335.740 186.310 ;
        RECT 1335.020 138.050 1335.280 138.370 ;
        RECT 1335.080 96.405 1335.220 138.050 ;
        RECT 1335.010 96.035 1335.290 96.405 ;
        RECT 1336.390 95.355 1336.670 95.725 ;
        RECT 1336.460 21.750 1336.600 95.355 ;
        RECT 1007.500 21.430 1007.760 21.750 ;
        RECT 1336.400 21.430 1336.660 21.750 ;
        RECT 1007.560 2.400 1007.700 21.430 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER via2 ;
        RECT 1336.390 1353.400 1336.670 1353.680 ;
        RECT 1335.010 1352.720 1335.290 1353.000 ;
        RECT 1335.010 1345.240 1335.290 1345.520 ;
        RECT 1335.930 1345.240 1336.210 1345.520 ;
        RECT 1335.010 820.960 1335.290 821.240 ;
        RECT 1336.390 820.280 1336.670 820.560 ;
        RECT 1335.010 772.680 1335.290 772.960 ;
        RECT 1336.390 772.680 1336.670 772.960 ;
        RECT 1335.010 96.080 1335.290 96.360 ;
        RECT 1336.390 95.400 1336.670 95.680 ;
      LAYER met3 ;
        RECT 1336.365 1353.690 1336.695 1353.705 ;
        RECT 1334.310 1353.390 1336.695 1353.690 ;
        RECT 1334.310 1353.010 1334.610 1353.390 ;
        RECT 1336.365 1353.375 1336.695 1353.390 ;
        RECT 1334.985 1353.010 1335.315 1353.025 ;
        RECT 1334.310 1352.710 1335.315 1353.010 ;
        RECT 1334.985 1352.695 1335.315 1352.710 ;
        RECT 1334.985 1345.530 1335.315 1345.545 ;
        RECT 1335.905 1345.530 1336.235 1345.545 ;
        RECT 1334.985 1345.230 1336.235 1345.530 ;
        RECT 1334.985 1345.215 1335.315 1345.230 ;
        RECT 1335.905 1345.215 1336.235 1345.230 ;
        RECT 1334.985 821.250 1335.315 821.265 ;
        RECT 1334.985 820.950 1336.450 821.250 ;
        RECT 1334.985 820.935 1335.315 820.950 ;
        RECT 1336.150 820.585 1336.450 820.950 ;
        RECT 1336.150 820.270 1336.695 820.585 ;
        RECT 1336.365 820.255 1336.695 820.270 ;
        RECT 1334.985 772.970 1335.315 772.985 ;
        RECT 1336.365 772.970 1336.695 772.985 ;
        RECT 1334.985 772.670 1336.695 772.970 ;
        RECT 1334.985 772.655 1335.315 772.670 ;
        RECT 1336.365 772.655 1336.695 772.670 ;
        RECT 1334.985 96.370 1335.315 96.385 ;
        RECT 1334.310 96.070 1335.315 96.370 ;
        RECT 1334.310 95.690 1334.610 96.070 ;
        RECT 1334.985 96.055 1335.315 96.070 ;
        RECT 1336.365 95.690 1336.695 95.705 ;
        RECT 1334.310 95.390 1336.695 95.690 ;
        RECT 1336.365 95.375 1336.695 95.390 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.870 1678.140 1532.190 1678.200 ;
        RECT 1534.630 1678.140 1534.950 1678.200 ;
        RECT 1531.870 1678.000 1534.950 1678.140 ;
        RECT 1531.870 1677.940 1532.190 1678.000 ;
        RECT 1534.630 1677.940 1534.950 1678.000 ;
      LAYER via ;
        RECT 1531.900 1677.940 1532.160 1678.200 ;
        RECT 1534.660 1677.940 1534.920 1678.200 ;
      LAYER met2 ;
        RECT 1535.965 1700.410 1536.245 1704.000 ;
        RECT 1534.720 1700.270 1536.245 1700.410 ;
        RECT 1534.720 1678.230 1534.860 1700.270 ;
        RECT 1535.965 1700.000 1536.245 1700.270 ;
        RECT 1531.900 1677.910 1532.160 1678.230 ;
        RECT 1534.660 1677.910 1534.920 1678.230 ;
        RECT 1531.960 24.325 1532.100 1677.910 ;
        RECT 1025.430 23.955 1025.710 24.325 ;
        RECT 1531.890 23.955 1532.170 24.325 ;
        RECT 1025.500 2.400 1025.640 23.955 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
      LAYER via2 ;
        RECT 1025.430 24.000 1025.710 24.280 ;
        RECT 1531.890 24.000 1532.170 24.280 ;
      LAYER met3 ;
        RECT 1025.405 24.290 1025.735 24.305 ;
        RECT 1531.865 24.290 1532.195 24.305 ;
        RECT 1025.405 23.990 1532.195 24.290 ;
        RECT 1025.405 23.975 1025.735 23.990 ;
        RECT 1531.865 23.975 1532.195 23.990 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.770 1678.140 1539.090 1678.200 ;
        RECT 1541.070 1678.140 1541.390 1678.200 ;
        RECT 1538.770 1678.000 1541.390 1678.140 ;
        RECT 1538.770 1677.940 1539.090 1678.000 ;
        RECT 1541.070 1677.940 1541.390 1678.000 ;
        RECT 1043.350 23.700 1043.670 23.760 ;
        RECT 1043.350 23.560 1525.200 23.700 ;
        RECT 1043.350 23.500 1043.670 23.560 ;
        RECT 1525.060 23.360 1525.200 23.560 ;
        RECT 1538.770 23.360 1539.090 23.420 ;
        RECT 1525.060 23.220 1539.090 23.360 ;
        RECT 1538.770 23.160 1539.090 23.220 ;
      LAYER via ;
        RECT 1538.800 1677.940 1539.060 1678.200 ;
        RECT 1541.100 1677.940 1541.360 1678.200 ;
        RECT 1043.380 23.500 1043.640 23.760 ;
        RECT 1538.800 23.160 1539.060 23.420 ;
      LAYER met2 ;
        RECT 1542.405 1700.410 1542.685 1704.000 ;
        RECT 1541.160 1700.270 1542.685 1700.410 ;
        RECT 1541.160 1678.230 1541.300 1700.270 ;
        RECT 1542.405 1700.000 1542.685 1700.270 ;
        RECT 1538.800 1677.910 1539.060 1678.230 ;
        RECT 1541.100 1677.910 1541.360 1678.230 ;
        RECT 1043.380 23.470 1043.640 23.790 ;
        RECT 1043.440 2.400 1043.580 23.470 ;
        RECT 1538.860 23.450 1539.000 1677.910 ;
        RECT 1538.800 23.130 1539.060 23.450 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.670 1678.140 1545.990 1678.200 ;
        RECT 1547.510 1678.140 1547.830 1678.200 ;
        RECT 1545.670 1678.000 1547.830 1678.140 ;
        RECT 1545.670 1677.940 1545.990 1678.000 ;
        RECT 1547.510 1677.940 1547.830 1678.000 ;
        RECT 1061.290 23.360 1061.610 23.420 ;
        RECT 1061.290 23.220 1524.740 23.360 ;
        RECT 1061.290 23.160 1061.610 23.220 ;
        RECT 1524.600 23.020 1524.740 23.220 ;
        RECT 1545.210 23.020 1545.530 23.080 ;
        RECT 1524.600 22.880 1545.530 23.020 ;
        RECT 1545.210 22.820 1545.530 22.880 ;
      LAYER via ;
        RECT 1545.700 1677.940 1545.960 1678.200 ;
        RECT 1547.540 1677.940 1547.800 1678.200 ;
        RECT 1061.320 23.160 1061.580 23.420 ;
        RECT 1545.240 22.820 1545.500 23.080 ;
      LAYER met2 ;
        RECT 1549.305 1700.410 1549.585 1704.000 ;
        RECT 1547.600 1700.270 1549.585 1700.410 ;
        RECT 1547.600 1678.230 1547.740 1700.270 ;
        RECT 1549.305 1700.000 1549.585 1700.270 ;
        RECT 1545.700 1677.910 1545.960 1678.230 ;
        RECT 1547.540 1677.910 1547.800 1678.230 ;
        RECT 1545.760 23.530 1545.900 1677.910 ;
        RECT 1061.320 23.130 1061.580 23.450 ;
        RECT 1545.300 23.390 1545.900 23.530 ;
        RECT 1061.380 2.400 1061.520 23.130 ;
        RECT 1545.300 23.110 1545.440 23.390 ;
        RECT 1545.240 22.790 1545.500 23.110 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1534.245 23.885 1535.335 24.055 ;
        RECT 1524.125 23.545 1525.675 23.715 ;
        RECT 1534.245 23.545 1534.415 23.885 ;
        RECT 1524.125 22.865 1524.295 23.545 ;
        RECT 1535.165 22.355 1535.335 23.885 ;
        RECT 1535.165 22.185 1535.795 22.355 ;
      LAYER mcon ;
        RECT 1525.505 23.545 1525.675 23.715 ;
        RECT 1535.625 22.185 1535.795 22.355 ;
      LAYER met1 ;
        RECT 1552.570 1678.140 1552.890 1678.200 ;
        RECT 1554.870 1678.140 1555.190 1678.200 ;
        RECT 1552.570 1678.000 1555.190 1678.140 ;
        RECT 1552.570 1677.940 1552.890 1678.000 ;
        RECT 1554.870 1677.940 1555.190 1678.000 ;
        RECT 1525.445 23.700 1525.735 23.745 ;
        RECT 1534.185 23.700 1534.475 23.745 ;
        RECT 1525.445 23.560 1534.475 23.700 ;
        RECT 1525.445 23.515 1525.735 23.560 ;
        RECT 1534.185 23.515 1534.475 23.560 ;
        RECT 1079.230 23.020 1079.550 23.080 ;
        RECT 1524.065 23.020 1524.355 23.065 ;
        RECT 1079.230 22.880 1524.355 23.020 ;
        RECT 1079.230 22.820 1079.550 22.880 ;
        RECT 1524.065 22.835 1524.355 22.880 ;
        RECT 1535.565 22.340 1535.855 22.385 ;
        RECT 1553.030 22.340 1553.350 22.400 ;
        RECT 1535.565 22.200 1553.350 22.340 ;
        RECT 1535.565 22.155 1535.855 22.200 ;
        RECT 1553.030 22.140 1553.350 22.200 ;
      LAYER via ;
        RECT 1552.600 1677.940 1552.860 1678.200 ;
        RECT 1554.900 1677.940 1555.160 1678.200 ;
        RECT 1079.260 22.820 1079.520 23.080 ;
        RECT 1553.060 22.140 1553.320 22.400 ;
      LAYER met2 ;
        RECT 1556.205 1700.410 1556.485 1704.000 ;
        RECT 1554.960 1700.270 1556.485 1700.410 ;
        RECT 1554.960 1678.230 1555.100 1700.270 ;
        RECT 1556.205 1700.000 1556.485 1700.270 ;
        RECT 1552.600 1677.910 1552.860 1678.230 ;
        RECT 1554.900 1677.910 1555.160 1678.230 ;
        RECT 1552.660 24.210 1552.800 1677.910 ;
        RECT 1552.660 24.070 1553.260 24.210 ;
        RECT 1079.260 22.790 1079.520 23.110 ;
        RECT 1079.320 2.400 1079.460 22.790 ;
        RECT 1553.120 22.430 1553.260 24.070 ;
        RECT 1553.060 22.110 1553.320 22.430 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.470 1678.820 1559.790 1678.880 ;
        RECT 1561.310 1678.820 1561.630 1678.880 ;
        RECT 1559.470 1678.680 1561.630 1678.820 ;
        RECT 1559.470 1678.620 1559.790 1678.680 ;
        RECT 1561.310 1678.620 1561.630 1678.680 ;
        RECT 1096.710 22.680 1097.030 22.740 ;
        RECT 1559.010 22.680 1559.330 22.740 ;
        RECT 1096.710 22.540 1559.330 22.680 ;
        RECT 1096.710 22.480 1097.030 22.540 ;
        RECT 1559.010 22.480 1559.330 22.540 ;
      LAYER via ;
        RECT 1559.500 1678.620 1559.760 1678.880 ;
        RECT 1561.340 1678.620 1561.600 1678.880 ;
        RECT 1096.740 22.480 1097.000 22.740 ;
        RECT 1559.040 22.480 1559.300 22.740 ;
      LAYER met2 ;
        RECT 1562.645 1700.410 1562.925 1704.000 ;
        RECT 1561.400 1700.270 1562.925 1700.410 ;
        RECT 1561.400 1678.910 1561.540 1700.270 ;
        RECT 1562.645 1700.000 1562.925 1700.270 ;
        RECT 1559.500 1678.590 1559.760 1678.910 ;
        RECT 1561.340 1678.590 1561.600 1678.910 ;
        RECT 1559.560 22.850 1559.700 1678.590 ;
        RECT 1559.100 22.770 1559.700 22.850 ;
        RECT 1096.740 22.450 1097.000 22.770 ;
        RECT 1559.040 22.710 1559.700 22.770 ;
        RECT 1559.040 22.450 1559.300 22.710 ;
        RECT 1096.800 2.400 1096.940 22.450 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1566.370 1678.140 1566.690 1678.200 ;
        RECT 1567.750 1678.140 1568.070 1678.200 ;
        RECT 1566.370 1678.000 1568.070 1678.140 ;
        RECT 1566.370 1677.940 1566.690 1678.000 ;
        RECT 1567.750 1677.940 1568.070 1678.000 ;
        RECT 1114.650 22.340 1114.970 22.400 ;
        RECT 1114.650 22.200 1535.320 22.340 ;
        RECT 1114.650 22.140 1114.970 22.200 ;
        RECT 1535.180 22.000 1535.320 22.200 ;
        RECT 1566.370 22.000 1566.690 22.060 ;
        RECT 1535.180 21.860 1566.690 22.000 ;
        RECT 1566.370 21.800 1566.690 21.860 ;
      LAYER via ;
        RECT 1566.400 1677.940 1566.660 1678.200 ;
        RECT 1567.780 1677.940 1568.040 1678.200 ;
        RECT 1114.680 22.140 1114.940 22.400 ;
        RECT 1566.400 21.800 1566.660 22.060 ;
      LAYER met2 ;
        RECT 1569.545 1700.410 1569.825 1704.000 ;
        RECT 1567.840 1700.270 1569.825 1700.410 ;
        RECT 1567.840 1678.230 1567.980 1700.270 ;
        RECT 1569.545 1700.000 1569.825 1700.270 ;
        RECT 1566.400 1677.910 1566.660 1678.230 ;
        RECT 1567.780 1677.910 1568.040 1678.230 ;
        RECT 1114.680 22.110 1114.940 22.430 ;
        RECT 1114.740 2.400 1114.880 22.110 ;
        RECT 1566.460 22.090 1566.600 1677.910 ;
        RECT 1566.400 21.770 1566.660 22.090 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1534.705 21.845 1534.875 23.715 ;
      LAYER mcon ;
        RECT 1534.705 23.545 1534.875 23.715 ;
      LAYER met1 ;
        RECT 1573.270 1676.440 1573.590 1676.500 ;
        RECT 1575.110 1676.440 1575.430 1676.500 ;
        RECT 1573.270 1676.300 1575.430 1676.440 ;
        RECT 1573.270 1676.240 1573.590 1676.300 ;
        RECT 1575.110 1676.240 1575.430 1676.300 ;
        RECT 1534.645 23.700 1534.935 23.745 ;
        RECT 1573.270 23.700 1573.590 23.760 ;
        RECT 1534.645 23.560 1573.590 23.700 ;
        RECT 1534.645 23.515 1534.935 23.560 ;
        RECT 1573.270 23.500 1573.590 23.560 ;
        RECT 1132.590 22.000 1132.910 22.060 ;
        RECT 1534.645 22.000 1534.935 22.045 ;
        RECT 1132.590 21.860 1534.935 22.000 ;
        RECT 1132.590 21.800 1132.910 21.860 ;
        RECT 1534.645 21.815 1534.935 21.860 ;
      LAYER via ;
        RECT 1573.300 1676.240 1573.560 1676.500 ;
        RECT 1575.140 1676.240 1575.400 1676.500 ;
        RECT 1573.300 23.500 1573.560 23.760 ;
        RECT 1132.620 21.800 1132.880 22.060 ;
      LAYER met2 ;
        RECT 1576.445 1700.410 1576.725 1704.000 ;
        RECT 1575.200 1700.270 1576.725 1700.410 ;
        RECT 1575.200 1676.530 1575.340 1700.270 ;
        RECT 1576.445 1700.000 1576.725 1700.270 ;
        RECT 1573.300 1676.210 1573.560 1676.530 ;
        RECT 1575.140 1676.210 1575.400 1676.530 ;
        RECT 1573.360 23.790 1573.500 1676.210 ;
        RECT 1573.300 23.470 1573.560 23.790 ;
        RECT 1132.620 21.770 1132.880 22.090 ;
        RECT 1132.680 2.400 1132.820 21.770 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1580.170 1655.020 1580.490 1655.080 ;
        RECT 1581.550 1655.020 1581.870 1655.080 ;
        RECT 1580.170 1654.880 1581.870 1655.020 ;
        RECT 1580.170 1654.820 1580.490 1654.880 ;
        RECT 1581.550 1654.820 1581.870 1654.880 ;
        RECT 1150.530 24.040 1150.850 24.100 ;
        RECT 1580.170 24.040 1580.490 24.100 ;
        RECT 1150.530 23.900 1580.490 24.040 ;
        RECT 1150.530 23.840 1150.850 23.900 ;
        RECT 1580.170 23.840 1580.490 23.900 ;
      LAYER via ;
        RECT 1580.200 1654.820 1580.460 1655.080 ;
        RECT 1581.580 1654.820 1581.840 1655.080 ;
        RECT 1150.560 23.840 1150.820 24.100 ;
        RECT 1580.200 23.840 1580.460 24.100 ;
      LAYER met2 ;
        RECT 1582.885 1700.410 1583.165 1704.000 ;
        RECT 1581.640 1700.270 1583.165 1700.410 ;
        RECT 1581.640 1655.110 1581.780 1700.270 ;
        RECT 1582.885 1700.000 1583.165 1700.270 ;
        RECT 1580.200 1654.790 1580.460 1655.110 ;
        RECT 1581.580 1654.790 1581.840 1655.110 ;
        RECT 1580.260 24.130 1580.400 1654.790 ;
        RECT 1150.560 23.810 1150.820 24.130 ;
        RECT 1580.200 23.810 1580.460 24.130 ;
        RECT 1150.620 2.400 1150.760 23.810 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 27.100 669.230 27.160 ;
        RECT 1400.770 27.100 1401.090 27.160 ;
        RECT 668.910 26.960 1401.090 27.100 ;
        RECT 668.910 26.900 669.230 26.960 ;
        RECT 1400.770 26.900 1401.090 26.960 ;
      LAYER via ;
        RECT 668.940 26.900 669.200 27.160 ;
        RECT 1400.800 26.900 1401.060 27.160 ;
      LAYER met2 ;
        RECT 1401.185 1700.410 1401.465 1704.000 ;
        RECT 1400.860 1700.270 1401.465 1700.410 ;
        RECT 1400.860 27.190 1401.000 1700.270 ;
        RECT 1401.185 1700.000 1401.465 1700.270 ;
        RECT 668.940 26.870 669.200 27.190 ;
        RECT 1400.800 26.870 1401.060 27.190 ;
        RECT 669.000 2.400 669.140 26.870 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.070 1678.480 1587.390 1678.540 ;
        RECT 1587.990 1678.480 1588.310 1678.540 ;
        RECT 1587.070 1678.340 1588.310 1678.480 ;
        RECT 1587.070 1678.280 1587.390 1678.340 ;
        RECT 1587.990 1678.280 1588.310 1678.340 ;
        RECT 1168.470 24.380 1168.790 24.440 ;
        RECT 1587.070 24.380 1587.390 24.440 ;
        RECT 1168.470 24.240 1587.390 24.380 ;
        RECT 1168.470 24.180 1168.790 24.240 ;
        RECT 1587.070 24.180 1587.390 24.240 ;
      LAYER via ;
        RECT 1587.100 1678.280 1587.360 1678.540 ;
        RECT 1588.020 1678.280 1588.280 1678.540 ;
        RECT 1168.500 24.180 1168.760 24.440 ;
        RECT 1587.100 24.180 1587.360 24.440 ;
      LAYER met2 ;
        RECT 1589.785 1700.410 1590.065 1704.000 ;
        RECT 1588.080 1700.270 1590.065 1700.410 ;
        RECT 1588.080 1678.570 1588.220 1700.270 ;
        RECT 1589.785 1700.000 1590.065 1700.270 ;
        RECT 1587.100 1678.250 1587.360 1678.570 ;
        RECT 1588.020 1678.250 1588.280 1678.570 ;
        RECT 1587.160 24.470 1587.300 1678.250 ;
        RECT 1168.500 24.150 1168.760 24.470 ;
        RECT 1587.100 24.150 1587.360 24.470 ;
        RECT 1168.560 2.400 1168.700 24.150 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.970 1665.900 1594.290 1665.960 ;
        RECT 1595.350 1665.900 1595.670 1665.960 ;
        RECT 1593.970 1665.760 1595.670 1665.900 ;
        RECT 1593.970 1665.700 1594.290 1665.760 ;
        RECT 1595.350 1665.700 1595.670 1665.760 ;
        RECT 1185.950 24.720 1186.270 24.780 ;
        RECT 1593.510 24.720 1593.830 24.780 ;
        RECT 1185.950 24.580 1593.830 24.720 ;
        RECT 1185.950 24.520 1186.270 24.580 ;
        RECT 1593.510 24.520 1593.830 24.580 ;
      LAYER via ;
        RECT 1594.000 1665.700 1594.260 1665.960 ;
        RECT 1595.380 1665.700 1595.640 1665.960 ;
        RECT 1185.980 24.520 1186.240 24.780 ;
        RECT 1593.540 24.520 1593.800 24.780 ;
      LAYER met2 ;
        RECT 1596.685 1700.410 1596.965 1704.000 ;
        RECT 1595.440 1700.270 1596.965 1700.410 ;
        RECT 1595.440 1665.990 1595.580 1700.270 ;
        RECT 1596.685 1700.000 1596.965 1700.270 ;
        RECT 1594.000 1665.670 1594.260 1665.990 ;
        RECT 1595.380 1665.670 1595.640 1665.990 ;
        RECT 1594.060 25.400 1594.200 1665.670 ;
        RECT 1593.600 25.260 1594.200 25.400 ;
        RECT 1593.600 24.810 1593.740 25.260 ;
        RECT 1185.980 24.490 1186.240 24.810 ;
        RECT 1593.540 24.490 1593.800 24.810 ;
        RECT 1186.040 2.400 1186.180 24.490 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 25.060 1204.210 25.120 ;
        RECT 1602.250 25.060 1602.570 25.120 ;
        RECT 1203.890 24.920 1602.570 25.060 ;
        RECT 1203.890 24.860 1204.210 24.920 ;
        RECT 1602.250 24.860 1602.570 24.920 ;
      LAYER via ;
        RECT 1203.920 24.860 1204.180 25.120 ;
        RECT 1602.280 24.860 1602.540 25.120 ;
      LAYER met2 ;
        RECT 1603.125 1700.410 1603.405 1704.000 ;
        RECT 1602.340 1700.270 1603.405 1700.410 ;
        RECT 1602.340 25.150 1602.480 1700.270 ;
        RECT 1603.125 1700.000 1603.405 1700.270 ;
        RECT 1203.920 24.830 1204.180 25.150 ;
        RECT 1602.280 24.830 1602.540 25.150 ;
        RECT 1203.980 2.400 1204.120 24.830 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.830 25.400 1222.150 25.460 ;
        RECT 1609.150 25.400 1609.470 25.460 ;
        RECT 1221.830 25.260 1609.470 25.400 ;
        RECT 1221.830 25.200 1222.150 25.260 ;
        RECT 1609.150 25.200 1609.470 25.260 ;
      LAYER via ;
        RECT 1221.860 25.200 1222.120 25.460 ;
        RECT 1609.180 25.200 1609.440 25.460 ;
      LAYER met2 ;
        RECT 1610.025 1700.410 1610.305 1704.000 ;
        RECT 1609.240 1700.270 1610.305 1700.410 ;
        RECT 1609.240 25.490 1609.380 1700.270 ;
        RECT 1610.025 1700.000 1610.305 1700.270 ;
        RECT 1221.860 25.170 1222.120 25.490 ;
        RECT 1609.180 25.170 1609.440 25.490 ;
        RECT 1221.920 2.400 1222.060 25.170 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1239.770 25.740 1240.090 25.800 ;
        RECT 1616.510 25.740 1616.830 25.800 ;
        RECT 1239.770 25.600 1616.830 25.740 ;
        RECT 1239.770 25.540 1240.090 25.600 ;
        RECT 1616.510 25.540 1616.830 25.600 ;
      LAYER via ;
        RECT 1239.800 25.540 1240.060 25.800 ;
        RECT 1616.540 25.540 1616.800 25.800 ;
      LAYER met2 ;
        RECT 1616.465 1700.000 1616.745 1704.000 ;
        RECT 1616.600 25.830 1616.740 1700.000 ;
        RECT 1239.800 25.510 1240.060 25.830 ;
        RECT 1616.540 25.510 1616.800 25.830 ;
        RECT 1239.860 2.400 1240.000 25.510 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1257.250 26.080 1257.570 26.140 ;
        RECT 1621.570 26.080 1621.890 26.140 ;
        RECT 1257.250 25.940 1621.890 26.080 ;
        RECT 1257.250 25.880 1257.570 25.940 ;
        RECT 1621.570 25.880 1621.890 25.940 ;
      LAYER via ;
        RECT 1257.280 25.880 1257.540 26.140 ;
        RECT 1621.600 25.880 1621.860 26.140 ;
      LAYER met2 ;
        RECT 1623.365 1700.410 1623.645 1704.000 ;
        RECT 1621.660 1700.270 1623.645 1700.410 ;
        RECT 1621.660 26.170 1621.800 1700.270 ;
        RECT 1623.365 1700.000 1623.645 1700.270 ;
        RECT 1257.280 25.850 1257.540 26.170 ;
        RECT 1621.600 25.850 1621.860 26.170 ;
        RECT 1257.340 2.400 1257.480 25.850 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1318.045 17.255 1318.215 17.595 ;
        RECT 1317.585 17.085 1318.215 17.255 ;
        RECT 1352.545 17.085 1353.175 17.255 ;
        RECT 1400.385 16.065 1400.555 17.255 ;
        RECT 1400.845 15.385 1401.015 16.575 ;
        RECT 1448.685 15.385 1448.855 17.255 ;
        RECT 1462.025 17.085 1463.115 17.255 ;
        RECT 1511.245 14.705 1511.415 17.255 ;
      LAYER mcon ;
        RECT 1318.045 17.425 1318.215 17.595 ;
        RECT 1353.005 17.085 1353.175 17.255 ;
        RECT 1400.385 17.085 1400.555 17.255 ;
        RECT 1448.685 17.085 1448.855 17.255 ;
        RECT 1462.945 17.085 1463.115 17.255 ;
        RECT 1511.245 17.085 1511.415 17.255 ;
        RECT 1400.845 16.405 1401.015 16.575 ;
      LAYER met1 ;
        RECT 1545.670 23.020 1545.990 23.080 ;
        RECT 1628.470 23.020 1628.790 23.080 ;
        RECT 1545.670 22.880 1628.790 23.020 ;
        RECT 1545.670 22.820 1545.990 22.880 ;
        RECT 1628.470 22.820 1628.790 22.880 ;
        RECT 1317.985 17.580 1318.275 17.625 ;
        RECT 1317.985 17.440 1352.700 17.580 ;
        RECT 1317.985 17.395 1318.275 17.440 ;
        RECT 1275.190 17.240 1275.510 17.300 ;
        RECT 1352.560 17.285 1352.700 17.440 ;
        RECT 1317.525 17.240 1317.815 17.285 ;
        RECT 1275.190 17.100 1317.815 17.240 ;
        RECT 1275.190 17.040 1275.510 17.100 ;
        RECT 1317.525 17.055 1317.815 17.100 ;
        RECT 1352.485 17.055 1352.775 17.285 ;
        RECT 1352.945 17.240 1353.235 17.285 ;
        RECT 1400.325 17.240 1400.615 17.285 ;
        RECT 1352.945 17.100 1400.615 17.240 ;
        RECT 1352.945 17.055 1353.235 17.100 ;
        RECT 1400.325 17.055 1400.615 17.100 ;
        RECT 1448.625 17.240 1448.915 17.285 ;
        RECT 1461.965 17.240 1462.255 17.285 ;
        RECT 1448.625 17.100 1462.255 17.240 ;
        RECT 1448.625 17.055 1448.915 17.100 ;
        RECT 1461.965 17.055 1462.255 17.100 ;
        RECT 1462.885 17.240 1463.175 17.285 ;
        RECT 1511.185 17.240 1511.475 17.285 ;
        RECT 1462.885 17.100 1511.475 17.240 ;
        RECT 1462.885 17.055 1463.175 17.100 ;
        RECT 1511.185 17.055 1511.475 17.100 ;
        RECT 1400.785 16.560 1401.075 16.605 ;
        RECT 1400.400 16.420 1401.075 16.560 ;
        RECT 1400.400 16.265 1400.540 16.420 ;
        RECT 1400.785 16.375 1401.075 16.420 ;
        RECT 1400.325 16.035 1400.615 16.265 ;
        RECT 1400.785 15.540 1401.075 15.585 ;
        RECT 1448.625 15.540 1448.915 15.585 ;
        RECT 1400.785 15.400 1448.915 15.540 ;
        RECT 1400.785 15.355 1401.075 15.400 ;
        RECT 1448.625 15.355 1448.915 15.400 ;
        RECT 1511.185 14.860 1511.475 14.905 ;
        RECT 1511.185 14.720 1518.300 14.860 ;
        RECT 1511.185 14.675 1511.475 14.720 ;
        RECT 1518.160 14.520 1518.300 14.720 ;
        RECT 1545.670 14.520 1545.990 14.580 ;
        RECT 1518.160 14.380 1545.990 14.520 ;
        RECT 1545.670 14.320 1545.990 14.380 ;
      LAYER via ;
        RECT 1545.700 22.820 1545.960 23.080 ;
        RECT 1628.500 22.820 1628.760 23.080 ;
        RECT 1275.220 17.040 1275.480 17.300 ;
        RECT 1545.700 14.320 1545.960 14.580 ;
      LAYER met2 ;
        RECT 1630.265 1700.410 1630.545 1704.000 ;
        RECT 1628.560 1700.270 1630.545 1700.410 ;
        RECT 1628.560 23.110 1628.700 1700.270 ;
        RECT 1630.265 1700.000 1630.545 1700.270 ;
        RECT 1545.700 22.790 1545.960 23.110 ;
        RECT 1628.500 22.790 1628.760 23.110 ;
        RECT 1275.220 17.010 1275.480 17.330 ;
        RECT 1275.280 2.400 1275.420 17.010 ;
        RECT 1545.760 14.610 1545.900 22.790 ;
        RECT 1545.700 14.290 1545.960 14.610 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1552.570 23.360 1552.890 23.420 ;
        RECT 1635.370 23.360 1635.690 23.420 ;
        RECT 1552.570 23.220 1635.690 23.360 ;
        RECT 1552.570 23.160 1552.890 23.220 ;
        RECT 1635.370 23.160 1635.690 23.220 ;
        RECT 1293.130 17.920 1293.450 17.980 ;
        RECT 1552.570 17.920 1552.890 17.980 ;
        RECT 1293.130 17.780 1552.890 17.920 ;
        RECT 1293.130 17.720 1293.450 17.780 ;
        RECT 1552.570 17.720 1552.890 17.780 ;
      LAYER via ;
        RECT 1552.600 23.160 1552.860 23.420 ;
        RECT 1635.400 23.160 1635.660 23.420 ;
        RECT 1293.160 17.720 1293.420 17.980 ;
        RECT 1552.600 17.720 1552.860 17.980 ;
      LAYER met2 ;
        RECT 1636.705 1700.410 1636.985 1704.000 ;
        RECT 1635.460 1700.270 1636.985 1700.410 ;
        RECT 1635.460 23.450 1635.600 1700.270 ;
        RECT 1636.705 1700.000 1636.985 1700.270 ;
        RECT 1552.600 23.130 1552.860 23.450 ;
        RECT 1635.400 23.130 1635.660 23.450 ;
        RECT 1552.660 18.010 1552.800 23.130 ;
        RECT 1293.160 17.690 1293.420 18.010 ;
        RECT 1552.600 17.690 1552.860 18.010 ;
        RECT 1293.220 2.400 1293.360 17.690 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1643.190 1559.280 1643.510 1559.540 ;
        RECT 1643.280 1558.520 1643.420 1559.280 ;
        RECT 1643.190 1558.260 1643.510 1558.520 ;
        RECT 1565.910 22.340 1566.230 22.400 ;
        RECT 1643.190 22.340 1643.510 22.400 ;
        RECT 1565.910 22.200 1643.510 22.340 ;
        RECT 1565.910 22.140 1566.230 22.200 ;
        RECT 1643.190 22.140 1643.510 22.200 ;
        RECT 1311.070 18.940 1311.390 19.000 ;
        RECT 1565.910 18.940 1566.230 19.000 ;
        RECT 1311.070 18.800 1566.230 18.940 ;
        RECT 1311.070 18.740 1311.390 18.800 ;
        RECT 1565.910 18.740 1566.230 18.800 ;
      LAYER via ;
        RECT 1643.220 1559.280 1643.480 1559.540 ;
        RECT 1643.220 1558.260 1643.480 1558.520 ;
        RECT 1565.940 22.140 1566.200 22.400 ;
        RECT 1643.220 22.140 1643.480 22.400 ;
        RECT 1311.100 18.740 1311.360 19.000 ;
        RECT 1565.940 18.740 1566.200 19.000 ;
      LAYER met2 ;
        RECT 1643.605 1700.000 1643.885 1704.000 ;
        RECT 1643.740 1656.210 1643.880 1700.000 ;
        RECT 1643.280 1656.070 1643.880 1656.210 ;
        RECT 1643.280 1559.570 1643.420 1656.070 ;
        RECT 1643.220 1559.250 1643.480 1559.570 ;
        RECT 1643.220 1558.230 1643.480 1558.550 ;
        RECT 1643.280 22.430 1643.420 1558.230 ;
        RECT 1565.940 22.110 1566.200 22.430 ;
        RECT 1643.220 22.110 1643.480 22.430 ;
        RECT 1566.000 19.030 1566.140 22.110 ;
        RECT 1311.100 18.710 1311.360 19.030 ;
        RECT 1565.940 18.710 1566.200 19.030 ;
        RECT 1311.160 2.400 1311.300 18.710 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1572.810 22.680 1573.130 22.740 ;
        RECT 1650.090 22.680 1650.410 22.740 ;
        RECT 1572.810 22.540 1650.410 22.680 ;
        RECT 1572.810 22.480 1573.130 22.540 ;
        RECT 1650.090 22.480 1650.410 22.540 ;
        RECT 1329.010 19.960 1329.330 20.020 ;
        RECT 1329.010 19.820 1359.600 19.960 ;
        RECT 1329.010 19.760 1329.330 19.820 ;
        RECT 1359.460 19.280 1359.600 19.820 ;
        RECT 1572.810 19.280 1573.130 19.340 ;
        RECT 1359.460 19.140 1573.130 19.280 ;
        RECT 1572.810 19.080 1573.130 19.140 ;
      LAYER via ;
        RECT 1572.840 22.480 1573.100 22.740 ;
        RECT 1650.120 22.480 1650.380 22.740 ;
        RECT 1329.040 19.760 1329.300 20.020 ;
        RECT 1572.840 19.080 1573.100 19.340 ;
      LAYER met2 ;
        RECT 1650.505 1700.410 1650.785 1704.000 ;
        RECT 1650.180 1700.270 1650.785 1700.410 ;
        RECT 1650.180 22.770 1650.320 1700.270 ;
        RECT 1650.505 1700.000 1650.785 1700.270 ;
        RECT 1572.840 22.450 1573.100 22.770 ;
        RECT 1650.120 22.450 1650.380 22.770 ;
        RECT 1329.040 19.730 1329.300 20.050 ;
        RECT 1329.100 2.400 1329.240 19.730 ;
        RECT 1572.900 19.370 1573.040 22.450 ;
        RECT 1572.840 19.050 1573.100 19.370 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 27.440 686.710 27.500 ;
        RECT 1407.670 27.440 1407.990 27.500 ;
        RECT 686.390 27.300 1407.990 27.440 ;
        RECT 686.390 27.240 686.710 27.300 ;
        RECT 1407.670 27.240 1407.990 27.300 ;
      LAYER via ;
        RECT 686.420 27.240 686.680 27.500 ;
        RECT 1407.700 27.240 1407.960 27.500 ;
      LAYER met2 ;
        RECT 1408.085 1700.410 1408.365 1704.000 ;
        RECT 1407.760 1700.270 1408.365 1700.410 ;
        RECT 1407.760 27.530 1407.900 1700.270 ;
        RECT 1408.085 1700.000 1408.365 1700.270 ;
        RECT 686.420 27.210 686.680 27.530 ;
        RECT 1407.700 27.210 1407.960 27.530 ;
        RECT 686.480 2.400 686.620 27.210 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1579.710 23.700 1580.030 23.760 ;
        RECT 1656.990 23.700 1657.310 23.760 ;
        RECT 1579.710 23.560 1657.310 23.700 ;
        RECT 1579.710 23.500 1580.030 23.560 ;
        RECT 1656.990 23.500 1657.310 23.560 ;
        RECT 1346.490 20.300 1346.810 20.360 ;
        RECT 1579.710 20.300 1580.030 20.360 ;
        RECT 1346.490 20.160 1580.030 20.300 ;
        RECT 1346.490 20.100 1346.810 20.160 ;
        RECT 1579.710 20.100 1580.030 20.160 ;
      LAYER via ;
        RECT 1579.740 23.500 1580.000 23.760 ;
        RECT 1657.020 23.500 1657.280 23.760 ;
        RECT 1346.520 20.100 1346.780 20.360 ;
        RECT 1579.740 20.100 1580.000 20.360 ;
      LAYER met2 ;
        RECT 1656.945 1700.000 1657.225 1704.000 ;
        RECT 1657.080 23.790 1657.220 1700.000 ;
        RECT 1579.740 23.470 1580.000 23.790 ;
        RECT 1657.020 23.470 1657.280 23.790 ;
        RECT 1579.800 20.390 1579.940 23.470 ;
        RECT 1346.520 20.070 1346.780 20.390 ;
        RECT 1579.740 20.070 1580.000 20.390 ;
        RECT 1346.580 2.400 1346.720 20.070 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.070 22.000 1587.390 22.060 ;
        RECT 1663.890 22.000 1664.210 22.060 ;
        RECT 1587.070 21.860 1664.210 22.000 ;
        RECT 1587.070 21.800 1587.390 21.860 ;
        RECT 1663.890 21.800 1664.210 21.860 ;
        RECT 1364.430 19.960 1364.750 20.020 ;
        RECT 1587.070 19.960 1587.390 20.020 ;
        RECT 1364.430 19.820 1587.390 19.960 ;
        RECT 1364.430 19.760 1364.750 19.820 ;
        RECT 1587.070 19.760 1587.390 19.820 ;
      LAYER via ;
        RECT 1587.100 21.800 1587.360 22.060 ;
        RECT 1663.920 21.800 1664.180 22.060 ;
        RECT 1364.460 19.760 1364.720 20.020 ;
        RECT 1587.100 19.760 1587.360 20.020 ;
      LAYER met2 ;
        RECT 1663.845 1700.000 1664.125 1704.000 ;
        RECT 1663.980 22.090 1664.120 1700.000 ;
        RECT 1587.100 21.770 1587.360 22.090 ;
        RECT 1663.920 21.770 1664.180 22.090 ;
        RECT 1587.160 20.050 1587.300 21.770 ;
        RECT 1364.460 19.730 1364.720 20.050 ;
        RECT 1587.100 19.730 1587.360 20.050 ;
        RECT 1364.520 2.400 1364.660 19.730 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 31.860 1421.330 31.920 ;
        RECT 1670.790 31.860 1671.110 31.920 ;
        RECT 1421.010 31.720 1671.110 31.860 ;
        RECT 1421.010 31.660 1421.330 31.720 ;
        RECT 1670.790 31.660 1671.110 31.720 ;
        RECT 1382.370 18.600 1382.690 18.660 ;
        RECT 1421.010 18.600 1421.330 18.660 ;
        RECT 1382.370 18.460 1421.330 18.600 ;
        RECT 1382.370 18.400 1382.690 18.460 ;
        RECT 1421.010 18.400 1421.330 18.460 ;
      LAYER via ;
        RECT 1421.040 31.660 1421.300 31.920 ;
        RECT 1670.820 31.660 1671.080 31.920 ;
        RECT 1382.400 18.400 1382.660 18.660 ;
        RECT 1421.040 18.400 1421.300 18.660 ;
      LAYER met2 ;
        RECT 1670.745 1700.000 1671.025 1704.000 ;
        RECT 1670.880 31.950 1671.020 1700.000 ;
        RECT 1421.040 31.630 1421.300 31.950 ;
        RECT 1670.820 31.630 1671.080 31.950 ;
        RECT 1421.100 18.690 1421.240 31.630 ;
        RECT 1382.400 18.370 1382.660 18.690 ;
        RECT 1421.040 18.370 1421.300 18.690 ;
        RECT 1382.460 2.400 1382.600 18.370 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 26.420 1400.630 26.480 ;
        RECT 1677.690 26.420 1678.010 26.480 ;
        RECT 1400.310 26.280 1678.010 26.420 ;
        RECT 1400.310 26.220 1400.630 26.280 ;
        RECT 1677.690 26.220 1678.010 26.280 ;
      LAYER via ;
        RECT 1400.340 26.220 1400.600 26.480 ;
        RECT 1677.720 26.220 1677.980 26.480 ;
      LAYER met2 ;
        RECT 1677.185 1700.410 1677.465 1704.000 ;
        RECT 1677.185 1700.270 1677.920 1700.410 ;
        RECT 1677.185 1700.000 1677.465 1700.270 ;
        RECT 1677.780 26.510 1677.920 1700.270 ;
        RECT 1400.340 26.190 1400.600 26.510 ;
        RECT 1677.720 26.190 1677.980 26.510 ;
        RECT 1400.400 2.400 1400.540 26.190 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.250 26.760 1418.570 26.820 ;
        RECT 1684.130 26.760 1684.450 26.820 ;
        RECT 1418.250 26.620 1684.450 26.760 ;
        RECT 1418.250 26.560 1418.570 26.620 ;
        RECT 1684.130 26.560 1684.450 26.620 ;
      LAYER via ;
        RECT 1418.280 26.560 1418.540 26.820 ;
        RECT 1684.160 26.560 1684.420 26.820 ;
      LAYER met2 ;
        RECT 1684.085 1700.000 1684.365 1704.000 ;
        RECT 1684.220 26.850 1684.360 1700.000 ;
        RECT 1418.280 26.530 1418.540 26.850 ;
        RECT 1684.160 26.530 1684.420 26.850 ;
        RECT 1418.340 2.400 1418.480 26.530 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1435.730 27.100 1436.050 27.160 ;
        RECT 1691.030 27.100 1691.350 27.160 ;
        RECT 1435.730 26.960 1691.350 27.100 ;
        RECT 1435.730 26.900 1436.050 26.960 ;
        RECT 1691.030 26.900 1691.350 26.960 ;
      LAYER via ;
        RECT 1435.760 26.900 1436.020 27.160 ;
        RECT 1691.060 26.900 1691.320 27.160 ;
      LAYER met2 ;
        RECT 1690.525 1700.410 1690.805 1704.000 ;
        RECT 1690.525 1700.270 1691.260 1700.410 ;
        RECT 1690.525 1700.000 1690.805 1700.270 ;
        RECT 1691.120 27.190 1691.260 1700.270 ;
        RECT 1435.760 26.870 1436.020 27.190 ;
        RECT 1691.060 26.870 1691.320 27.190 ;
        RECT 1435.820 2.400 1435.960 26.870 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1453.670 27.440 1453.990 27.500 ;
        RECT 1697.930 27.440 1698.250 27.500 ;
        RECT 1453.670 27.300 1698.250 27.440 ;
        RECT 1453.670 27.240 1453.990 27.300 ;
        RECT 1697.930 27.240 1698.250 27.300 ;
      LAYER via ;
        RECT 1453.700 27.240 1453.960 27.500 ;
        RECT 1697.960 27.240 1698.220 27.500 ;
      LAYER met2 ;
        RECT 1697.425 1700.410 1697.705 1704.000 ;
        RECT 1697.425 1700.270 1698.160 1700.410 ;
        RECT 1697.425 1700.000 1697.705 1700.270 ;
        RECT 1698.020 27.530 1698.160 1700.270 ;
        RECT 1453.700 27.210 1453.960 27.530 ;
        RECT 1697.960 27.210 1698.220 27.530 ;
        RECT 1453.760 2.400 1453.900 27.210 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.610 21.660 1471.930 21.720 ;
        RECT 1704.830 21.660 1705.150 21.720 ;
        RECT 1471.610 21.520 1705.150 21.660 ;
        RECT 1471.610 21.460 1471.930 21.520 ;
        RECT 1704.830 21.460 1705.150 21.520 ;
      LAYER via ;
        RECT 1471.640 21.460 1471.900 21.720 ;
        RECT 1704.860 21.460 1705.120 21.720 ;
      LAYER met2 ;
        RECT 1704.325 1700.410 1704.605 1704.000 ;
        RECT 1704.325 1700.270 1705.060 1700.410 ;
        RECT 1704.325 1700.000 1704.605 1700.270 ;
        RECT 1704.920 21.750 1705.060 1700.270 ;
        RECT 1471.640 21.430 1471.900 21.750 ;
        RECT 1704.860 21.430 1705.120 21.750 ;
        RECT 1471.700 2.400 1471.840 21.430 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 21.320 1490.330 21.380 ;
        RECT 1705.290 21.320 1705.610 21.380 ;
        RECT 1490.010 21.180 1705.610 21.320 ;
        RECT 1490.010 21.120 1490.330 21.180 ;
        RECT 1705.290 21.120 1705.610 21.180 ;
      LAYER via ;
        RECT 1490.040 21.120 1490.300 21.380 ;
        RECT 1705.320 21.120 1705.580 21.380 ;
      LAYER met2 ;
        RECT 1710.765 1700.410 1711.045 1704.000 ;
        RECT 1709.520 1700.270 1711.045 1700.410 ;
        RECT 1709.520 1677.970 1709.660 1700.270 ;
        RECT 1710.765 1700.000 1711.045 1700.270 ;
        RECT 1705.380 1677.830 1709.660 1677.970 ;
        RECT 1705.380 21.410 1705.520 1677.830 ;
        RECT 1490.040 21.090 1490.300 21.410 ;
        RECT 1705.320 21.090 1705.580 21.410 ;
        RECT 1490.100 10.610 1490.240 21.090 ;
        RECT 1489.640 10.470 1490.240 10.610 ;
        RECT 1489.640 2.400 1489.780 10.470 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1712.725 1545.725 1712.895 1593.835 ;
        RECT 1712.265 1490.645 1712.435 1538.755 ;
        RECT 1712.725 1352.605 1712.895 1400.715 ;
        RECT 1712.725 1256.045 1712.895 1304.155 ;
        RECT 1712.725 524.705 1712.895 572.475 ;
        RECT 1712.725 476.085 1712.895 524.195 ;
        RECT 1712.725 234.685 1712.895 255.935 ;
        RECT 1712.265 48.365 1712.435 137.955 ;
      LAYER mcon ;
        RECT 1712.725 1593.665 1712.895 1593.835 ;
        RECT 1712.265 1538.585 1712.435 1538.755 ;
        RECT 1712.725 1400.545 1712.895 1400.715 ;
        RECT 1712.725 1303.985 1712.895 1304.155 ;
        RECT 1712.725 572.305 1712.895 572.475 ;
        RECT 1712.725 524.025 1712.895 524.195 ;
        RECT 1712.725 255.765 1712.895 255.935 ;
        RECT 1712.265 137.785 1712.435 137.955 ;
      LAYER met1 ;
        RECT 1712.650 1593.820 1712.970 1593.880 ;
        RECT 1712.455 1593.680 1712.970 1593.820 ;
        RECT 1712.650 1593.620 1712.970 1593.680 ;
        RECT 1712.650 1545.880 1712.970 1545.940 ;
        RECT 1712.455 1545.740 1712.970 1545.880 ;
        RECT 1712.650 1545.680 1712.970 1545.740 ;
        RECT 1712.190 1538.740 1712.510 1538.800 ;
        RECT 1711.995 1538.600 1712.510 1538.740 ;
        RECT 1712.190 1538.540 1712.510 1538.600 ;
        RECT 1712.205 1490.800 1712.495 1490.845 ;
        RECT 1712.650 1490.800 1712.970 1490.860 ;
        RECT 1712.205 1490.660 1712.970 1490.800 ;
        RECT 1712.205 1490.615 1712.495 1490.660 ;
        RECT 1712.650 1490.600 1712.970 1490.660 ;
        RECT 1712.650 1463.060 1712.970 1463.320 ;
        RECT 1712.740 1462.640 1712.880 1463.060 ;
        RECT 1712.650 1462.380 1712.970 1462.640 ;
        RECT 1712.650 1400.700 1712.970 1400.760 ;
        RECT 1712.455 1400.560 1712.970 1400.700 ;
        RECT 1712.650 1400.500 1712.970 1400.560 ;
        RECT 1712.650 1352.760 1712.970 1352.820 ;
        RECT 1712.455 1352.620 1712.970 1352.760 ;
        RECT 1712.650 1352.560 1712.970 1352.620 ;
        RECT 1712.650 1304.140 1712.970 1304.200 ;
        RECT 1712.455 1304.000 1712.970 1304.140 ;
        RECT 1712.650 1303.940 1712.970 1304.000 ;
        RECT 1712.650 1256.200 1712.970 1256.260 ;
        RECT 1712.455 1256.060 1712.970 1256.200 ;
        RECT 1712.650 1256.000 1712.970 1256.060 ;
        RECT 1711.730 1159.300 1712.050 1159.360 ;
        RECT 1712.650 1159.300 1712.970 1159.360 ;
        RECT 1711.730 1159.160 1712.970 1159.300 ;
        RECT 1711.730 1159.100 1712.050 1159.160 ;
        RECT 1712.650 1159.100 1712.970 1159.160 ;
        RECT 1711.730 1062.740 1712.050 1062.800 ;
        RECT 1712.650 1062.740 1712.970 1062.800 ;
        RECT 1711.730 1062.600 1712.970 1062.740 ;
        RECT 1711.730 1062.540 1712.050 1062.600 ;
        RECT 1712.650 1062.540 1712.970 1062.600 ;
        RECT 1711.730 917.900 1712.050 917.960 ;
        RECT 1712.650 917.900 1712.970 917.960 ;
        RECT 1711.730 917.760 1712.970 917.900 ;
        RECT 1711.730 917.700 1712.050 917.760 ;
        RECT 1712.650 917.700 1712.970 917.760 ;
        RECT 1712.650 814.200 1712.970 814.260 ;
        RECT 1713.110 814.200 1713.430 814.260 ;
        RECT 1712.650 814.060 1713.430 814.200 ;
        RECT 1712.650 814.000 1712.970 814.060 ;
        RECT 1713.110 814.000 1713.430 814.060 ;
        RECT 1712.650 572.460 1712.970 572.520 ;
        RECT 1712.455 572.320 1712.970 572.460 ;
        RECT 1712.650 572.260 1712.970 572.320 ;
        RECT 1712.650 524.860 1712.970 524.920 ;
        RECT 1712.455 524.720 1712.970 524.860 ;
        RECT 1712.650 524.660 1712.970 524.720 ;
        RECT 1712.650 524.180 1712.970 524.240 ;
        RECT 1712.455 524.040 1712.970 524.180 ;
        RECT 1712.650 523.980 1712.970 524.040 ;
        RECT 1712.650 476.240 1712.970 476.300 ;
        RECT 1712.455 476.100 1712.970 476.240 ;
        RECT 1712.650 476.040 1712.970 476.100 ;
        RECT 1712.650 400.560 1712.970 400.820 ;
        RECT 1712.740 400.140 1712.880 400.560 ;
        RECT 1712.650 399.880 1712.970 400.140 ;
        RECT 1712.650 255.920 1712.970 255.980 ;
        RECT 1712.455 255.780 1712.970 255.920 ;
        RECT 1712.650 255.720 1712.970 255.780 ;
        RECT 1712.650 234.840 1712.970 234.900 ;
        RECT 1712.455 234.700 1712.970 234.840 ;
        RECT 1712.650 234.640 1712.970 234.700 ;
        RECT 1712.190 145.220 1712.510 145.480 ;
        RECT 1712.280 145.080 1712.420 145.220 ;
        RECT 1712.650 145.080 1712.970 145.140 ;
        RECT 1712.280 144.940 1712.970 145.080 ;
        RECT 1712.650 144.880 1712.970 144.940 ;
        RECT 1712.205 137.940 1712.495 137.985 ;
        RECT 1712.650 137.940 1712.970 138.000 ;
        RECT 1712.205 137.800 1712.970 137.940 ;
        RECT 1712.205 137.755 1712.495 137.800 ;
        RECT 1712.650 137.740 1712.970 137.800 ;
        RECT 1712.190 48.520 1712.510 48.580 ;
        RECT 1711.995 48.380 1712.510 48.520 ;
        RECT 1712.190 48.320 1712.510 48.380 ;
        RECT 1507.030 20.980 1507.350 21.040 ;
        RECT 1712.190 20.980 1712.510 21.040 ;
        RECT 1507.030 20.840 1712.510 20.980 ;
        RECT 1507.030 20.780 1507.350 20.840 ;
        RECT 1712.190 20.780 1712.510 20.840 ;
      LAYER via ;
        RECT 1712.680 1593.620 1712.940 1593.880 ;
        RECT 1712.680 1545.680 1712.940 1545.940 ;
        RECT 1712.220 1538.540 1712.480 1538.800 ;
        RECT 1712.680 1490.600 1712.940 1490.860 ;
        RECT 1712.680 1463.060 1712.940 1463.320 ;
        RECT 1712.680 1462.380 1712.940 1462.640 ;
        RECT 1712.680 1400.500 1712.940 1400.760 ;
        RECT 1712.680 1352.560 1712.940 1352.820 ;
        RECT 1712.680 1303.940 1712.940 1304.200 ;
        RECT 1712.680 1256.000 1712.940 1256.260 ;
        RECT 1711.760 1159.100 1712.020 1159.360 ;
        RECT 1712.680 1159.100 1712.940 1159.360 ;
        RECT 1711.760 1062.540 1712.020 1062.800 ;
        RECT 1712.680 1062.540 1712.940 1062.800 ;
        RECT 1711.760 917.700 1712.020 917.960 ;
        RECT 1712.680 917.700 1712.940 917.960 ;
        RECT 1712.680 814.000 1712.940 814.260 ;
        RECT 1713.140 814.000 1713.400 814.260 ;
        RECT 1712.680 572.260 1712.940 572.520 ;
        RECT 1712.680 524.660 1712.940 524.920 ;
        RECT 1712.680 523.980 1712.940 524.240 ;
        RECT 1712.680 476.040 1712.940 476.300 ;
        RECT 1712.680 400.560 1712.940 400.820 ;
        RECT 1712.680 399.880 1712.940 400.140 ;
        RECT 1712.680 255.720 1712.940 255.980 ;
        RECT 1712.680 234.640 1712.940 234.900 ;
        RECT 1712.220 145.220 1712.480 145.480 ;
        RECT 1712.680 144.880 1712.940 145.140 ;
        RECT 1712.680 137.740 1712.940 138.000 ;
        RECT 1712.220 48.320 1712.480 48.580 ;
        RECT 1507.060 20.780 1507.320 21.040 ;
        RECT 1712.220 20.780 1712.480 21.040 ;
      LAYER met2 ;
        RECT 1717.665 1700.410 1717.945 1704.000 ;
        RECT 1716.420 1700.270 1717.945 1700.410 ;
        RECT 1716.420 1677.970 1716.560 1700.270 ;
        RECT 1717.665 1700.000 1717.945 1700.270 ;
        RECT 1712.740 1677.830 1716.560 1677.970 ;
        RECT 1712.740 1608.610 1712.880 1677.830 ;
        RECT 1712.740 1608.470 1713.340 1608.610 ;
        RECT 1713.200 1594.330 1713.340 1608.470 ;
        RECT 1712.740 1594.190 1713.340 1594.330 ;
        RECT 1712.740 1593.910 1712.880 1594.190 ;
        RECT 1712.680 1593.590 1712.940 1593.910 ;
        RECT 1712.680 1545.880 1712.940 1545.970 ;
        RECT 1712.280 1545.740 1712.940 1545.880 ;
        RECT 1712.280 1538.830 1712.420 1545.740 ;
        RECT 1712.680 1545.650 1712.940 1545.740 ;
        RECT 1712.220 1538.510 1712.480 1538.830 ;
        RECT 1712.680 1490.570 1712.940 1490.890 ;
        RECT 1712.740 1463.350 1712.880 1490.570 ;
        RECT 1712.680 1463.030 1712.940 1463.350 ;
        RECT 1712.680 1462.350 1712.940 1462.670 ;
        RECT 1712.740 1400.790 1712.880 1462.350 ;
        RECT 1712.680 1400.470 1712.940 1400.790 ;
        RECT 1712.680 1352.530 1712.940 1352.850 ;
        RECT 1712.740 1304.230 1712.880 1352.530 ;
        RECT 1712.680 1303.910 1712.940 1304.230 ;
        RECT 1712.680 1255.970 1712.940 1256.290 ;
        RECT 1712.740 1207.525 1712.880 1255.970 ;
        RECT 1711.750 1207.155 1712.030 1207.525 ;
        RECT 1712.670 1207.155 1712.950 1207.525 ;
        RECT 1711.820 1159.390 1711.960 1207.155 ;
        RECT 1711.760 1159.070 1712.020 1159.390 ;
        RECT 1712.680 1159.070 1712.940 1159.390 ;
        RECT 1712.740 1110.965 1712.880 1159.070 ;
        RECT 1711.750 1110.595 1712.030 1110.965 ;
        RECT 1712.670 1110.595 1712.950 1110.965 ;
        RECT 1711.820 1062.830 1711.960 1110.595 ;
        RECT 1711.760 1062.510 1712.020 1062.830 ;
        RECT 1712.680 1062.510 1712.940 1062.830 ;
        RECT 1712.740 980.290 1712.880 1062.510 ;
        RECT 1712.280 980.150 1712.880 980.290 ;
        RECT 1712.280 979.610 1712.420 980.150 ;
        RECT 1712.280 979.470 1712.880 979.610 ;
        RECT 1712.740 966.125 1712.880 979.470 ;
        RECT 1711.750 965.755 1712.030 966.125 ;
        RECT 1712.670 965.755 1712.950 966.125 ;
        RECT 1711.820 917.990 1711.960 965.755 ;
        RECT 1711.760 917.670 1712.020 917.990 ;
        RECT 1712.680 917.670 1712.940 917.990 ;
        RECT 1712.740 821.965 1712.880 917.670 ;
        RECT 1712.670 821.595 1712.950 821.965 ;
        RECT 1712.670 820.915 1712.950 821.285 ;
        RECT 1712.740 814.290 1712.880 820.915 ;
        RECT 1712.680 813.970 1712.940 814.290 ;
        RECT 1713.140 813.970 1713.400 814.290 ;
        RECT 1713.200 676.330 1713.340 813.970 ;
        RECT 1712.740 676.190 1713.340 676.330 ;
        RECT 1712.740 595.410 1712.880 676.190 ;
        RECT 1712.740 595.270 1713.800 595.410 ;
        RECT 1713.660 573.085 1713.800 595.270 ;
        RECT 1712.670 572.715 1712.950 573.085 ;
        RECT 1713.590 572.715 1713.870 573.085 ;
        RECT 1712.740 572.550 1712.880 572.715 ;
        RECT 1712.680 572.230 1712.940 572.550 ;
        RECT 1712.680 524.630 1712.940 524.950 ;
        RECT 1712.740 524.270 1712.880 524.630 ;
        RECT 1712.680 523.950 1712.940 524.270 ;
        RECT 1712.680 476.010 1712.940 476.330 ;
        RECT 1712.740 400.850 1712.880 476.010 ;
        RECT 1712.680 400.530 1712.940 400.850 ;
        RECT 1712.680 399.850 1712.940 400.170 ;
        RECT 1712.740 256.010 1712.880 399.850 ;
        RECT 1712.680 255.690 1712.940 256.010 ;
        RECT 1712.680 234.610 1712.940 234.930 ;
        RECT 1712.740 234.330 1712.880 234.610 ;
        RECT 1712.280 234.190 1712.880 234.330 ;
        RECT 1712.280 145.510 1712.420 234.190 ;
        RECT 1712.220 145.190 1712.480 145.510 ;
        RECT 1712.680 144.850 1712.940 145.170 ;
        RECT 1712.740 138.030 1712.880 144.850 ;
        RECT 1712.680 137.710 1712.940 138.030 ;
        RECT 1712.220 48.290 1712.480 48.610 ;
        RECT 1712.280 21.070 1712.420 48.290 ;
        RECT 1507.060 20.750 1507.320 21.070 ;
        RECT 1712.220 20.750 1712.480 21.070 ;
        RECT 1507.120 2.400 1507.260 20.750 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
      LAYER via2 ;
        RECT 1711.750 1207.200 1712.030 1207.480 ;
        RECT 1712.670 1207.200 1712.950 1207.480 ;
        RECT 1711.750 1110.640 1712.030 1110.920 ;
        RECT 1712.670 1110.640 1712.950 1110.920 ;
        RECT 1711.750 965.800 1712.030 966.080 ;
        RECT 1712.670 965.800 1712.950 966.080 ;
        RECT 1712.670 821.640 1712.950 821.920 ;
        RECT 1712.670 820.960 1712.950 821.240 ;
        RECT 1712.670 572.760 1712.950 573.040 ;
        RECT 1713.590 572.760 1713.870 573.040 ;
      LAYER met3 ;
        RECT 1711.725 1207.490 1712.055 1207.505 ;
        RECT 1712.645 1207.490 1712.975 1207.505 ;
        RECT 1711.725 1207.190 1712.975 1207.490 ;
        RECT 1711.725 1207.175 1712.055 1207.190 ;
        RECT 1712.645 1207.175 1712.975 1207.190 ;
        RECT 1711.725 1110.930 1712.055 1110.945 ;
        RECT 1712.645 1110.930 1712.975 1110.945 ;
        RECT 1711.725 1110.630 1712.975 1110.930 ;
        RECT 1711.725 1110.615 1712.055 1110.630 ;
        RECT 1712.645 1110.615 1712.975 1110.630 ;
        RECT 1711.725 966.090 1712.055 966.105 ;
        RECT 1712.645 966.090 1712.975 966.105 ;
        RECT 1711.725 965.790 1712.975 966.090 ;
        RECT 1711.725 965.775 1712.055 965.790 ;
        RECT 1712.645 965.775 1712.975 965.790 ;
        RECT 1712.645 821.930 1712.975 821.945 ;
        RECT 1712.645 821.630 1713.650 821.930 ;
        RECT 1712.645 821.615 1712.975 821.630 ;
        RECT 1712.645 821.250 1712.975 821.265 ;
        RECT 1713.350 821.250 1713.650 821.630 ;
        RECT 1712.645 820.950 1713.650 821.250 ;
        RECT 1712.645 820.935 1712.975 820.950 ;
        RECT 1712.645 573.050 1712.975 573.065 ;
        RECT 1713.565 573.050 1713.895 573.065 ;
        RECT 1712.645 572.750 1713.895 573.050 ;
        RECT 1712.645 572.735 1712.975 572.750 ;
        RECT 1713.565 572.735 1713.895 572.750 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 704.330 59.740 704.650 59.800 ;
        RECT 1415.490 59.740 1415.810 59.800 ;
        RECT 704.330 59.600 1415.810 59.740 ;
        RECT 704.330 59.540 704.650 59.600 ;
        RECT 1415.490 59.540 1415.810 59.600 ;
      LAYER via ;
        RECT 704.360 59.540 704.620 59.800 ;
        RECT 1415.520 59.540 1415.780 59.800 ;
      LAYER met2 ;
        RECT 1414.525 1700.410 1414.805 1704.000 ;
        RECT 1414.525 1700.270 1415.720 1700.410 ;
        RECT 1414.525 1700.000 1414.805 1700.270 ;
        RECT 1415.580 59.830 1415.720 1700.270 ;
        RECT 704.360 59.510 704.620 59.830 ;
        RECT 1415.520 59.510 1415.780 59.830 ;
        RECT 704.420 2.400 704.560 59.510 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1719.165 1642.285 1719.335 1677.815 ;
        RECT 1718.705 1013.965 1718.875 1055.615 ;
        RECT 1719.625 766.105 1719.795 814.215 ;
        RECT 1719.165 676.345 1719.335 741.795 ;
        RECT 1718.705 379.865 1718.875 427.635 ;
        RECT 1718.705 331.245 1718.875 379.355 ;
      LAYER mcon ;
        RECT 1719.165 1677.645 1719.335 1677.815 ;
        RECT 1718.705 1055.445 1718.875 1055.615 ;
        RECT 1719.625 814.045 1719.795 814.215 ;
        RECT 1719.165 741.625 1719.335 741.795 ;
        RECT 1718.705 427.465 1718.875 427.635 ;
        RECT 1718.705 379.185 1718.875 379.355 ;
      LAYER met1 ;
        RECT 1719.105 1677.800 1719.395 1677.845 ;
        RECT 1722.770 1677.800 1723.090 1677.860 ;
        RECT 1719.105 1677.660 1723.090 1677.800 ;
        RECT 1719.105 1677.615 1719.395 1677.660 ;
        RECT 1722.770 1677.600 1723.090 1677.660 ;
        RECT 1719.090 1642.440 1719.410 1642.500 ;
        RECT 1718.895 1642.300 1719.410 1642.440 ;
        RECT 1719.090 1642.240 1719.410 1642.300 ;
        RECT 1719.090 1062.740 1719.410 1062.800 ;
        RECT 1718.720 1062.600 1719.410 1062.740 ;
        RECT 1718.720 1062.460 1718.860 1062.600 ;
        RECT 1719.090 1062.540 1719.410 1062.600 ;
        RECT 1718.630 1062.200 1718.950 1062.460 ;
        RECT 1718.630 1055.600 1718.950 1055.660 ;
        RECT 1718.435 1055.460 1718.950 1055.600 ;
        RECT 1718.630 1055.400 1718.950 1055.460 ;
        RECT 1718.630 1014.120 1718.950 1014.180 ;
        RECT 1718.435 1013.980 1718.950 1014.120 ;
        RECT 1718.630 1013.920 1718.950 1013.980 ;
        RECT 1719.090 917.560 1719.410 917.620 ;
        RECT 1719.550 917.560 1719.870 917.620 ;
        RECT 1719.090 917.420 1719.870 917.560 ;
        RECT 1719.090 917.360 1719.410 917.420 ;
        RECT 1719.550 917.360 1719.870 917.420 ;
        RECT 1719.550 910.760 1719.870 910.820 ;
        RECT 1720.470 910.760 1720.790 910.820 ;
        RECT 1719.550 910.620 1720.790 910.760 ;
        RECT 1719.550 910.560 1719.870 910.620 ;
        RECT 1720.470 910.560 1720.790 910.620 ;
        RECT 1719.550 814.200 1719.870 814.260 ;
        RECT 1719.355 814.060 1719.870 814.200 ;
        RECT 1719.550 814.000 1719.870 814.060 ;
        RECT 1719.550 766.260 1719.870 766.320 ;
        RECT 1719.355 766.120 1719.870 766.260 ;
        RECT 1719.550 766.060 1719.870 766.120 ;
        RECT 1719.105 741.780 1719.395 741.825 ;
        RECT 1719.550 741.780 1719.870 741.840 ;
        RECT 1719.105 741.640 1719.870 741.780 ;
        RECT 1719.105 741.595 1719.395 741.640 ;
        RECT 1719.550 741.580 1719.870 741.640 ;
        RECT 1719.090 676.500 1719.410 676.560 ;
        RECT 1718.895 676.360 1719.410 676.500 ;
        RECT 1719.090 676.300 1719.410 676.360 ;
        RECT 1718.630 434.760 1718.950 434.820 ;
        RECT 1719.090 434.760 1719.410 434.820 ;
        RECT 1718.630 434.620 1719.410 434.760 ;
        RECT 1718.630 434.560 1718.950 434.620 ;
        RECT 1719.090 434.560 1719.410 434.620 ;
        RECT 1718.630 427.620 1718.950 427.680 ;
        RECT 1718.435 427.480 1718.950 427.620 ;
        RECT 1718.630 427.420 1718.950 427.480 ;
        RECT 1718.630 380.020 1718.950 380.080 ;
        RECT 1718.435 379.880 1718.950 380.020 ;
        RECT 1718.630 379.820 1718.950 379.880 ;
        RECT 1718.630 379.340 1718.950 379.400 ;
        RECT 1718.435 379.200 1718.950 379.340 ;
        RECT 1718.630 379.140 1718.950 379.200 ;
        RECT 1718.645 331.400 1718.935 331.445 ;
        RECT 1719.550 331.400 1719.870 331.460 ;
        RECT 1718.645 331.260 1719.870 331.400 ;
        RECT 1718.645 331.215 1718.935 331.260 ;
        RECT 1719.550 331.200 1719.870 331.260 ;
        RECT 1524.970 32.200 1525.290 32.260 ;
        RECT 1718.630 32.200 1718.950 32.260 ;
        RECT 1524.970 32.060 1718.950 32.200 ;
        RECT 1524.970 32.000 1525.290 32.060 ;
        RECT 1718.630 32.000 1718.950 32.060 ;
      LAYER via ;
        RECT 1722.800 1677.600 1723.060 1677.860 ;
        RECT 1719.120 1642.240 1719.380 1642.500 ;
        RECT 1719.120 1062.540 1719.380 1062.800 ;
        RECT 1718.660 1062.200 1718.920 1062.460 ;
        RECT 1718.660 1055.400 1718.920 1055.660 ;
        RECT 1718.660 1013.920 1718.920 1014.180 ;
        RECT 1719.120 917.360 1719.380 917.620 ;
        RECT 1719.580 917.360 1719.840 917.620 ;
        RECT 1719.580 910.560 1719.840 910.820 ;
        RECT 1720.500 910.560 1720.760 910.820 ;
        RECT 1719.580 814.000 1719.840 814.260 ;
        RECT 1719.580 766.060 1719.840 766.320 ;
        RECT 1719.580 741.580 1719.840 741.840 ;
        RECT 1719.120 676.300 1719.380 676.560 ;
        RECT 1718.660 434.560 1718.920 434.820 ;
        RECT 1719.120 434.560 1719.380 434.820 ;
        RECT 1718.660 427.420 1718.920 427.680 ;
        RECT 1718.660 379.820 1718.920 380.080 ;
        RECT 1718.660 379.140 1718.920 379.400 ;
        RECT 1719.580 331.200 1719.840 331.460 ;
        RECT 1525.000 32.000 1525.260 32.260 ;
        RECT 1718.660 32.000 1718.920 32.260 ;
      LAYER met2 ;
        RECT 1724.565 1700.410 1724.845 1704.000 ;
        RECT 1722.860 1700.270 1724.845 1700.410 ;
        RECT 1722.860 1677.890 1723.000 1700.270 ;
        RECT 1724.565 1700.000 1724.845 1700.270 ;
        RECT 1722.800 1677.570 1723.060 1677.890 ;
        RECT 1719.120 1642.210 1719.380 1642.530 ;
        RECT 1719.180 1414.810 1719.320 1642.210 ;
        RECT 1718.720 1414.670 1719.320 1414.810 ;
        RECT 1718.720 1414.130 1718.860 1414.670 ;
        RECT 1718.720 1413.990 1719.320 1414.130 ;
        RECT 1719.180 1318.250 1719.320 1413.990 ;
        RECT 1718.720 1318.110 1719.320 1318.250 ;
        RECT 1718.720 1317.570 1718.860 1318.110 ;
        RECT 1718.720 1317.430 1719.320 1317.570 ;
        RECT 1719.180 1221.690 1719.320 1317.430 ;
        RECT 1718.720 1221.550 1719.320 1221.690 ;
        RECT 1718.720 1221.010 1718.860 1221.550 ;
        RECT 1718.720 1220.870 1719.320 1221.010 ;
        RECT 1719.180 1125.130 1719.320 1220.870 ;
        RECT 1718.720 1124.990 1719.320 1125.130 ;
        RECT 1718.720 1124.450 1718.860 1124.990 ;
        RECT 1718.720 1124.310 1719.320 1124.450 ;
        RECT 1719.180 1062.830 1719.320 1124.310 ;
        RECT 1719.120 1062.510 1719.380 1062.830 ;
        RECT 1718.660 1062.170 1718.920 1062.490 ;
        RECT 1718.720 1055.690 1718.860 1062.170 ;
        RECT 1718.660 1055.370 1718.920 1055.690 ;
        RECT 1718.660 1013.890 1718.920 1014.210 ;
        RECT 1718.720 980.290 1718.860 1013.890 ;
        RECT 1718.260 980.150 1718.860 980.290 ;
        RECT 1718.260 966.010 1718.400 980.150 ;
        RECT 1718.260 965.870 1719.320 966.010 ;
        RECT 1719.180 917.650 1719.320 965.870 ;
        RECT 1719.120 917.330 1719.380 917.650 ;
        RECT 1719.580 917.330 1719.840 917.650 ;
        RECT 1719.640 910.850 1719.780 917.330 ;
        RECT 1719.580 910.530 1719.840 910.850 ;
        RECT 1720.500 910.530 1720.760 910.850 ;
        RECT 1720.560 862.765 1720.700 910.530 ;
        RECT 1719.570 862.395 1719.850 862.765 ;
        RECT 1720.490 862.395 1720.770 862.765 ;
        RECT 1719.640 821.965 1719.780 862.395 ;
        RECT 1719.570 821.595 1719.850 821.965 ;
        RECT 1719.570 820.915 1719.850 821.285 ;
        RECT 1719.640 814.290 1719.780 820.915 ;
        RECT 1719.580 813.970 1719.840 814.290 ;
        RECT 1719.580 766.030 1719.840 766.350 ;
        RECT 1719.640 741.870 1719.780 766.030 ;
        RECT 1719.580 741.550 1719.840 741.870 ;
        RECT 1719.120 676.270 1719.380 676.590 ;
        RECT 1719.180 545.770 1719.320 676.270 ;
        RECT 1718.720 545.630 1719.320 545.770 ;
        RECT 1718.720 545.090 1718.860 545.630 ;
        RECT 1718.720 544.950 1719.320 545.090 ;
        RECT 1719.180 434.850 1719.320 544.950 ;
        RECT 1718.660 434.530 1718.920 434.850 ;
        RECT 1719.120 434.530 1719.380 434.850 ;
        RECT 1718.720 427.710 1718.860 434.530 ;
        RECT 1718.660 427.390 1718.920 427.710 ;
        RECT 1718.660 379.790 1718.920 380.110 ;
        RECT 1718.720 379.430 1718.860 379.790 ;
        RECT 1718.660 379.110 1718.920 379.430 ;
        RECT 1719.580 331.170 1719.840 331.490 ;
        RECT 1719.640 303.690 1719.780 331.170 ;
        RECT 1719.180 303.550 1719.780 303.690 ;
        RECT 1719.180 207.130 1719.320 303.550 ;
        RECT 1718.720 206.990 1719.320 207.130 ;
        RECT 1718.720 206.450 1718.860 206.990 ;
        RECT 1718.720 206.310 1719.320 206.450 ;
        RECT 1719.180 62.290 1719.320 206.310 ;
        RECT 1718.720 62.150 1719.320 62.290 ;
        RECT 1718.720 32.290 1718.860 62.150 ;
        RECT 1525.000 31.970 1525.260 32.290 ;
        RECT 1718.660 31.970 1718.920 32.290 ;
        RECT 1525.060 2.400 1525.200 31.970 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
      LAYER via2 ;
        RECT 1719.570 862.440 1719.850 862.720 ;
        RECT 1720.490 862.440 1720.770 862.720 ;
        RECT 1719.570 821.640 1719.850 821.920 ;
        RECT 1719.570 820.960 1719.850 821.240 ;
      LAYER met3 ;
        RECT 1719.545 862.730 1719.875 862.745 ;
        RECT 1720.465 862.730 1720.795 862.745 ;
        RECT 1719.545 862.430 1720.795 862.730 ;
        RECT 1719.545 862.415 1719.875 862.430 ;
        RECT 1720.465 862.415 1720.795 862.430 ;
        RECT 1719.545 821.930 1719.875 821.945 ;
        RECT 1718.870 821.630 1719.875 821.930 ;
        RECT 1718.870 821.250 1719.170 821.630 ;
        RECT 1719.545 821.615 1719.875 821.630 ;
        RECT 1719.545 821.250 1719.875 821.265 ;
        RECT 1718.870 820.950 1719.875 821.250 ;
        RECT 1719.545 820.935 1719.875 820.950 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1725.530 1678.140 1725.850 1678.200 ;
        RECT 1729.670 1678.140 1729.990 1678.200 ;
        RECT 1725.530 1678.000 1729.990 1678.140 ;
        RECT 1725.530 1677.940 1725.850 1678.000 ;
        RECT 1729.670 1677.940 1729.990 1678.000 ;
        RECT 1725.530 966.320 1725.850 966.580 ;
        RECT 1725.620 965.900 1725.760 966.320 ;
        RECT 1725.530 965.640 1725.850 965.900 ;
        RECT 1583.390 24.040 1583.710 24.100 ;
        RECT 1725.530 24.040 1725.850 24.100 ;
        RECT 1583.390 23.900 1725.850 24.040 ;
        RECT 1583.390 23.840 1583.710 23.900 ;
        RECT 1725.530 23.840 1725.850 23.900 ;
        RECT 1542.910 14.180 1543.230 14.240 ;
        RECT 1583.390 14.180 1583.710 14.240 ;
        RECT 1542.910 14.040 1583.710 14.180 ;
        RECT 1542.910 13.980 1543.230 14.040 ;
        RECT 1583.390 13.980 1583.710 14.040 ;
      LAYER via ;
        RECT 1725.560 1677.940 1725.820 1678.200 ;
        RECT 1729.700 1677.940 1729.960 1678.200 ;
        RECT 1725.560 966.320 1725.820 966.580 ;
        RECT 1725.560 965.640 1725.820 965.900 ;
        RECT 1583.420 23.840 1583.680 24.100 ;
        RECT 1725.560 23.840 1725.820 24.100 ;
        RECT 1542.940 13.980 1543.200 14.240 ;
        RECT 1583.420 13.980 1583.680 14.240 ;
      LAYER met2 ;
        RECT 1731.005 1700.410 1731.285 1704.000 ;
        RECT 1729.760 1700.270 1731.285 1700.410 ;
        RECT 1729.760 1678.230 1729.900 1700.270 ;
        RECT 1731.005 1700.000 1731.285 1700.270 ;
        RECT 1725.560 1677.910 1725.820 1678.230 ;
        RECT 1729.700 1677.910 1729.960 1678.230 ;
        RECT 1725.620 966.610 1725.760 1677.910 ;
        RECT 1725.560 966.290 1725.820 966.610 ;
        RECT 1725.560 965.610 1725.820 965.930 ;
        RECT 1725.620 24.130 1725.760 965.610 ;
        RECT 1583.420 23.810 1583.680 24.130 ;
        RECT 1725.560 23.810 1725.820 24.130 ;
        RECT 1583.480 14.270 1583.620 23.810 ;
        RECT 1542.940 13.950 1543.200 14.270 ;
        RECT 1583.420 13.950 1583.680 14.270 ;
        RECT 1543.000 2.400 1543.140 13.950 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1732.965 227.885 1733.135 255.935 ;
        RECT 1732.045 83.045 1732.215 131.155 ;
      LAYER mcon ;
        RECT 1732.965 255.765 1733.135 255.935 ;
        RECT 1732.045 130.985 1732.215 131.155 ;
      LAYER met1 ;
        RECT 1732.890 1642.440 1733.210 1642.500 ;
        RECT 1736.570 1642.440 1736.890 1642.500 ;
        RECT 1732.890 1642.300 1736.890 1642.440 ;
        RECT 1732.890 1642.240 1733.210 1642.300 ;
        RECT 1736.570 1642.240 1736.890 1642.300 ;
        RECT 1732.890 931.640 1733.210 931.900 ;
        RECT 1732.980 931.160 1733.120 931.640 ;
        RECT 1733.350 931.160 1733.670 931.220 ;
        RECT 1732.980 931.020 1733.670 931.160 ;
        RECT 1733.350 930.960 1733.670 931.020 ;
        RECT 1732.430 835.280 1732.750 835.340 ;
        RECT 1733.350 835.280 1733.670 835.340 ;
        RECT 1732.430 835.140 1733.670 835.280 ;
        RECT 1732.430 835.080 1732.750 835.140 ;
        RECT 1733.350 835.080 1733.670 835.140 ;
        RECT 1732.890 676.500 1733.210 676.560 ;
        RECT 1733.350 676.500 1733.670 676.560 ;
        RECT 1732.890 676.360 1733.670 676.500 ;
        RECT 1732.890 676.300 1733.210 676.360 ;
        RECT 1733.350 676.300 1733.670 676.360 ;
        RECT 1732.890 352.280 1733.210 352.540 ;
        RECT 1732.980 351.860 1733.120 352.280 ;
        RECT 1732.890 351.600 1733.210 351.860 ;
        RECT 1732.890 255.920 1733.210 255.980 ;
        RECT 1732.695 255.780 1733.210 255.920 ;
        RECT 1732.890 255.720 1733.210 255.780 ;
        RECT 1732.890 228.040 1733.210 228.100 ;
        RECT 1732.695 227.900 1733.210 228.040 ;
        RECT 1732.890 227.840 1733.210 227.900 ;
        RECT 1731.985 131.140 1732.275 131.185 ;
        RECT 1732.890 131.140 1733.210 131.200 ;
        RECT 1731.985 131.000 1733.210 131.140 ;
        RECT 1731.985 130.955 1732.275 131.000 ;
        RECT 1732.890 130.940 1733.210 131.000 ;
        RECT 1731.970 83.200 1732.290 83.260 ;
        RECT 1731.775 83.060 1732.290 83.200 ;
        RECT 1731.970 83.000 1732.290 83.060 ;
        RECT 1593.970 24.720 1594.290 24.780 ;
        RECT 1731.970 24.720 1732.290 24.780 ;
        RECT 1593.970 24.580 1732.290 24.720 ;
        RECT 1593.970 24.520 1594.290 24.580 ;
        RECT 1731.970 24.520 1732.290 24.580 ;
        RECT 1560.850 17.920 1561.170 17.980 ;
        RECT 1593.970 17.920 1594.290 17.980 ;
        RECT 1560.850 17.780 1594.290 17.920 ;
        RECT 1560.850 17.720 1561.170 17.780 ;
        RECT 1593.970 17.720 1594.290 17.780 ;
      LAYER via ;
        RECT 1732.920 1642.240 1733.180 1642.500 ;
        RECT 1736.600 1642.240 1736.860 1642.500 ;
        RECT 1732.920 931.640 1733.180 931.900 ;
        RECT 1733.380 930.960 1733.640 931.220 ;
        RECT 1732.460 835.080 1732.720 835.340 ;
        RECT 1733.380 835.080 1733.640 835.340 ;
        RECT 1732.920 676.300 1733.180 676.560 ;
        RECT 1733.380 676.300 1733.640 676.560 ;
        RECT 1732.920 352.280 1733.180 352.540 ;
        RECT 1732.920 351.600 1733.180 351.860 ;
        RECT 1732.920 255.720 1733.180 255.980 ;
        RECT 1732.920 227.840 1733.180 228.100 ;
        RECT 1732.920 130.940 1733.180 131.200 ;
        RECT 1732.000 83.000 1732.260 83.260 ;
        RECT 1594.000 24.520 1594.260 24.780 ;
        RECT 1732.000 24.520 1732.260 24.780 ;
        RECT 1560.880 17.720 1561.140 17.980 ;
        RECT 1594.000 17.720 1594.260 17.980 ;
      LAYER met2 ;
        RECT 1737.905 1700.410 1738.185 1704.000 ;
        RECT 1736.660 1700.270 1738.185 1700.410 ;
        RECT 1736.660 1642.530 1736.800 1700.270 ;
        RECT 1737.905 1700.000 1738.185 1700.270 ;
        RECT 1732.920 1642.210 1733.180 1642.530 ;
        RECT 1736.600 1642.210 1736.860 1642.530 ;
        RECT 1732.980 1414.810 1733.120 1642.210 ;
        RECT 1732.520 1414.670 1733.120 1414.810 ;
        RECT 1732.520 1414.130 1732.660 1414.670 ;
        RECT 1732.520 1413.990 1733.120 1414.130 ;
        RECT 1732.980 1318.250 1733.120 1413.990 ;
        RECT 1732.520 1318.110 1733.120 1318.250 ;
        RECT 1732.520 1317.570 1732.660 1318.110 ;
        RECT 1732.520 1317.430 1733.120 1317.570 ;
        RECT 1732.980 1221.690 1733.120 1317.430 ;
        RECT 1732.520 1221.550 1733.120 1221.690 ;
        RECT 1732.520 1221.010 1732.660 1221.550 ;
        RECT 1732.520 1220.870 1733.120 1221.010 ;
        RECT 1732.980 1125.130 1733.120 1220.870 ;
        RECT 1732.520 1124.990 1733.120 1125.130 ;
        RECT 1732.520 1124.450 1732.660 1124.990 ;
        RECT 1732.520 1124.310 1733.120 1124.450 ;
        RECT 1732.980 1028.570 1733.120 1124.310 ;
        RECT 1732.520 1028.430 1733.120 1028.570 ;
        RECT 1732.520 1027.890 1732.660 1028.430 ;
        RECT 1732.520 1027.750 1733.120 1027.890 ;
        RECT 1732.980 931.930 1733.120 1027.750 ;
        RECT 1732.920 931.610 1733.180 931.930 ;
        RECT 1733.380 930.930 1733.640 931.250 ;
        RECT 1733.440 835.370 1733.580 930.930 ;
        RECT 1732.460 835.050 1732.720 835.370 ;
        RECT 1733.380 835.050 1733.640 835.370 ;
        RECT 1732.520 834.770 1732.660 835.050 ;
        RECT 1732.520 834.630 1733.580 834.770 ;
        RECT 1733.440 676.590 1733.580 834.630 ;
        RECT 1732.920 676.270 1733.180 676.590 ;
        RECT 1733.380 676.270 1733.640 676.590 ;
        RECT 1732.980 545.770 1733.120 676.270 ;
        RECT 1732.520 545.630 1733.120 545.770 ;
        RECT 1732.520 545.090 1732.660 545.630 ;
        RECT 1732.520 544.950 1733.120 545.090 ;
        RECT 1732.980 352.570 1733.120 544.950 ;
        RECT 1732.920 352.250 1733.180 352.570 ;
        RECT 1732.920 351.570 1733.180 351.890 ;
        RECT 1732.980 256.010 1733.120 351.570 ;
        RECT 1732.920 255.690 1733.180 256.010 ;
        RECT 1732.920 227.810 1733.180 228.130 ;
        RECT 1732.980 203.730 1733.120 227.810 ;
        RECT 1732.520 203.590 1733.120 203.730 ;
        RECT 1732.520 162.250 1732.660 203.590 ;
        RECT 1732.520 162.110 1733.120 162.250 ;
        RECT 1732.980 131.230 1733.120 162.110 ;
        RECT 1732.920 130.910 1733.180 131.230 ;
        RECT 1732.000 82.970 1732.260 83.290 ;
        RECT 1732.060 24.810 1732.200 82.970 ;
        RECT 1594.000 24.490 1594.260 24.810 ;
        RECT 1732.000 24.490 1732.260 24.810 ;
        RECT 1594.060 18.010 1594.200 24.490 ;
        RECT 1560.880 17.690 1561.140 18.010 ;
        RECT 1594.000 17.690 1594.260 18.010 ;
        RECT 1560.940 2.400 1561.080 17.690 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.330 1666.580 1739.650 1666.640 ;
        RECT 1743.470 1666.580 1743.790 1666.640 ;
        RECT 1739.330 1666.440 1743.790 1666.580 ;
        RECT 1739.330 1666.380 1739.650 1666.440 ;
        RECT 1743.470 1666.380 1743.790 1666.440 ;
        RECT 1600.870 24.380 1601.190 24.440 ;
        RECT 1739.330 24.380 1739.650 24.440 ;
        RECT 1600.870 24.240 1739.650 24.380 ;
        RECT 1600.870 24.180 1601.190 24.240 ;
        RECT 1739.330 24.180 1739.650 24.240 ;
        RECT 1578.790 18.940 1579.110 19.000 ;
        RECT 1600.870 18.940 1601.190 19.000 ;
        RECT 1578.790 18.800 1601.190 18.940 ;
        RECT 1578.790 18.740 1579.110 18.800 ;
        RECT 1600.870 18.740 1601.190 18.800 ;
      LAYER via ;
        RECT 1739.360 1666.380 1739.620 1666.640 ;
        RECT 1743.500 1666.380 1743.760 1666.640 ;
        RECT 1600.900 24.180 1601.160 24.440 ;
        RECT 1739.360 24.180 1739.620 24.440 ;
        RECT 1578.820 18.740 1579.080 19.000 ;
        RECT 1600.900 18.740 1601.160 19.000 ;
      LAYER met2 ;
        RECT 1744.805 1700.410 1745.085 1704.000 ;
        RECT 1743.560 1700.270 1745.085 1700.410 ;
        RECT 1743.560 1666.670 1743.700 1700.270 ;
        RECT 1744.805 1700.000 1745.085 1700.270 ;
        RECT 1739.360 1666.350 1739.620 1666.670 ;
        RECT 1743.500 1666.350 1743.760 1666.670 ;
        RECT 1739.420 24.470 1739.560 1666.350 ;
        RECT 1600.900 24.150 1601.160 24.470 ;
        RECT 1739.360 24.150 1739.620 24.470 ;
        RECT 1600.960 19.030 1601.100 24.150 ;
        RECT 1578.820 18.710 1579.080 19.030 ;
        RECT 1600.900 18.710 1601.160 19.030 ;
        RECT 1578.880 2.400 1579.020 18.710 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1723.690 1684.600 1724.010 1684.660 ;
        RECT 1751.290 1684.600 1751.610 1684.660 ;
        RECT 1723.690 1684.460 1751.610 1684.600 ;
        RECT 1723.690 1684.400 1724.010 1684.460 ;
        RECT 1751.290 1684.400 1751.610 1684.460 ;
        RECT 1596.270 20.300 1596.590 20.360 ;
        RECT 1721.850 20.300 1722.170 20.360 ;
        RECT 1596.270 20.160 1722.170 20.300 ;
        RECT 1596.270 20.100 1596.590 20.160 ;
        RECT 1721.850 20.100 1722.170 20.160 ;
      LAYER via ;
        RECT 1723.720 1684.400 1723.980 1684.660 ;
        RECT 1751.320 1684.400 1751.580 1684.660 ;
        RECT 1596.300 20.100 1596.560 20.360 ;
        RECT 1721.880 20.100 1722.140 20.360 ;
      LAYER met2 ;
        RECT 1751.245 1700.000 1751.525 1704.000 ;
        RECT 1751.380 1684.690 1751.520 1700.000 ;
        RECT 1723.720 1684.370 1723.980 1684.690 ;
        RECT 1751.320 1684.370 1751.580 1684.690 ;
        RECT 1723.780 1676.610 1723.920 1684.370 ;
        RECT 1721.940 1676.470 1723.920 1676.610 ;
        RECT 1721.940 20.390 1722.080 1676.470 ;
        RECT 1596.300 20.070 1596.560 20.390 ;
        RECT 1721.880 20.070 1722.140 20.390 ;
        RECT 1596.360 2.400 1596.500 20.070 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1632.685 14.365 1632.855 15.215 ;
      LAYER mcon ;
        RECT 1632.685 15.045 1632.855 15.215 ;
      LAYER met1 ;
        RECT 1728.750 1689.700 1729.070 1689.760 ;
        RECT 1758.190 1689.700 1758.510 1689.760 ;
        RECT 1728.750 1689.560 1758.510 1689.700 ;
        RECT 1728.750 1689.500 1729.070 1689.560 ;
        RECT 1758.190 1689.500 1758.510 1689.560 ;
        RECT 1632.625 15.200 1632.915 15.245 ;
        RECT 1728.750 15.200 1729.070 15.260 ;
        RECT 1632.625 15.060 1729.070 15.200 ;
        RECT 1632.625 15.015 1632.915 15.060 ;
        RECT 1728.750 15.000 1729.070 15.060 ;
        RECT 1614.210 14.520 1614.530 14.580 ;
        RECT 1632.625 14.520 1632.915 14.565 ;
        RECT 1614.210 14.380 1632.915 14.520 ;
        RECT 1614.210 14.320 1614.530 14.380 ;
        RECT 1632.625 14.335 1632.915 14.380 ;
      LAYER via ;
        RECT 1728.780 1689.500 1729.040 1689.760 ;
        RECT 1758.220 1689.500 1758.480 1689.760 ;
        RECT 1728.780 15.000 1729.040 15.260 ;
        RECT 1614.240 14.320 1614.500 14.580 ;
      LAYER met2 ;
        RECT 1758.145 1700.000 1758.425 1704.000 ;
        RECT 1758.280 1689.790 1758.420 1700.000 ;
        RECT 1728.780 1689.470 1729.040 1689.790 ;
        RECT 1758.220 1689.470 1758.480 1689.790 ;
        RECT 1728.840 15.290 1728.980 1689.470 ;
        RECT 1728.780 14.970 1729.040 15.290 ;
        RECT 1614.240 14.290 1614.500 14.610 ;
        RECT 1614.300 2.400 1614.440 14.290 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1676.385 14.025 1676.555 19.975 ;
      LAYER mcon ;
        RECT 1676.385 19.805 1676.555 19.975 ;
      LAYER met1 ;
        RECT 1760.030 1689.360 1760.350 1689.420 ;
        RECT 1763.710 1689.360 1764.030 1689.420 ;
        RECT 1760.030 1689.220 1764.030 1689.360 ;
        RECT 1760.030 1689.160 1760.350 1689.220 ;
        RECT 1763.710 1689.160 1764.030 1689.220 ;
        RECT 1676.325 19.960 1676.615 20.005 ;
        RECT 1760.030 19.960 1760.350 20.020 ;
        RECT 1676.325 19.820 1760.350 19.960 ;
        RECT 1676.325 19.775 1676.615 19.820 ;
        RECT 1760.030 19.760 1760.350 19.820 ;
        RECT 1632.150 14.180 1632.470 14.240 ;
        RECT 1676.325 14.180 1676.615 14.225 ;
        RECT 1632.150 14.040 1676.615 14.180 ;
        RECT 1632.150 13.980 1632.470 14.040 ;
        RECT 1676.325 13.995 1676.615 14.040 ;
      LAYER via ;
        RECT 1760.060 1689.160 1760.320 1689.420 ;
        RECT 1763.740 1689.160 1764.000 1689.420 ;
        RECT 1760.060 19.760 1760.320 20.020 ;
        RECT 1632.180 13.980 1632.440 14.240 ;
      LAYER met2 ;
        RECT 1765.045 1700.410 1765.325 1704.000 ;
        RECT 1763.800 1700.270 1765.325 1700.410 ;
        RECT 1763.800 1689.450 1763.940 1700.270 ;
        RECT 1765.045 1700.000 1765.325 1700.270 ;
        RECT 1760.060 1689.130 1760.320 1689.450 ;
        RECT 1763.740 1689.130 1764.000 1689.450 ;
        RECT 1760.120 20.050 1760.260 1689.130 ;
        RECT 1760.060 19.730 1760.320 20.050 ;
        RECT 1632.180 13.950 1632.440 14.270 ;
        RECT 1632.240 2.400 1632.380 13.950 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1700.305 1686.825 1700.475 1688.695 ;
        RECT 1727.445 1683.765 1727.615 1686.995 ;
      LAYER mcon ;
        RECT 1700.305 1688.525 1700.475 1688.695 ;
        RECT 1727.445 1686.825 1727.615 1686.995 ;
      LAYER met1 ;
        RECT 1655.610 1688.680 1655.930 1688.740 ;
        RECT 1700.245 1688.680 1700.535 1688.725 ;
        RECT 1655.610 1688.540 1700.535 1688.680 ;
        RECT 1655.610 1688.480 1655.930 1688.540 ;
        RECT 1700.245 1688.495 1700.535 1688.540 ;
        RECT 1700.245 1686.980 1700.535 1687.025 ;
        RECT 1727.385 1686.980 1727.675 1687.025 ;
        RECT 1700.245 1686.840 1727.675 1686.980 ;
        RECT 1700.245 1686.795 1700.535 1686.840 ;
        RECT 1727.385 1686.795 1727.675 1686.840 ;
        RECT 1727.385 1683.920 1727.675 1683.965 ;
        RECT 1771.530 1683.920 1771.850 1683.980 ;
        RECT 1727.385 1683.780 1771.850 1683.920 ;
        RECT 1727.385 1683.735 1727.675 1683.780 ;
        RECT 1771.530 1683.720 1771.850 1683.780 ;
        RECT 1650.090 19.960 1650.410 20.020 ;
        RECT 1655.610 19.960 1655.930 20.020 ;
        RECT 1650.090 19.820 1655.930 19.960 ;
        RECT 1650.090 19.760 1650.410 19.820 ;
        RECT 1655.610 19.760 1655.930 19.820 ;
      LAYER via ;
        RECT 1655.640 1688.480 1655.900 1688.740 ;
        RECT 1771.560 1683.720 1771.820 1683.980 ;
        RECT 1650.120 19.760 1650.380 20.020 ;
        RECT 1655.640 19.760 1655.900 20.020 ;
      LAYER met2 ;
        RECT 1771.485 1700.000 1771.765 1704.000 ;
        RECT 1655.640 1688.450 1655.900 1688.770 ;
        RECT 1655.700 20.050 1655.840 1688.450 ;
        RECT 1771.620 1684.010 1771.760 1700.000 ;
        RECT 1771.560 1683.690 1771.820 1684.010 ;
        RECT 1650.120 19.730 1650.380 20.050 ;
        RECT 1655.640 19.730 1655.900 20.050 ;
        RECT 1650.180 2.400 1650.320 19.730 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1669.410 1687.320 1669.730 1687.380 ;
        RECT 1778.430 1687.320 1778.750 1687.380 ;
        RECT 1669.410 1687.180 1778.750 1687.320 ;
        RECT 1669.410 1687.120 1669.730 1687.180 ;
        RECT 1778.430 1687.120 1778.750 1687.180 ;
      LAYER via ;
        RECT 1669.440 1687.120 1669.700 1687.380 ;
        RECT 1778.460 1687.120 1778.720 1687.380 ;
      LAYER met2 ;
        RECT 1778.385 1700.000 1778.665 1704.000 ;
        RECT 1778.520 1687.410 1778.660 1700.000 ;
        RECT 1669.440 1687.090 1669.700 1687.410 ;
        RECT 1778.460 1687.090 1778.720 1687.410 ;
        RECT 1669.500 3.130 1669.640 1687.090 ;
        RECT 1668.120 2.990 1669.640 3.130 ;
        RECT 1668.120 2.400 1668.260 2.990 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1701.225 1686.485 1701.395 1688.015 ;
      LAYER mcon ;
        RECT 1701.225 1687.845 1701.395 1688.015 ;
      LAYER met1 ;
        RECT 1701.165 1688.000 1701.455 1688.045 ;
        RECT 1784.870 1688.000 1785.190 1688.060 ;
        RECT 1701.165 1687.860 1785.190 1688.000 ;
        RECT 1701.165 1687.815 1701.455 1687.860 ;
        RECT 1784.870 1687.800 1785.190 1687.860 ;
        RECT 1690.110 1686.640 1690.430 1686.700 ;
        RECT 1701.165 1686.640 1701.455 1686.685 ;
        RECT 1690.110 1686.500 1701.455 1686.640 ;
        RECT 1690.110 1686.440 1690.430 1686.500 ;
        RECT 1701.165 1686.455 1701.455 1686.500 ;
        RECT 1690.110 904.440 1690.430 904.700 ;
        RECT 1690.200 904.020 1690.340 904.440 ;
        RECT 1690.110 903.760 1690.430 904.020 ;
        RECT 1685.510 18.600 1685.830 18.660 ;
        RECT 1690.110 18.600 1690.430 18.660 ;
        RECT 1685.510 18.460 1690.430 18.600 ;
        RECT 1685.510 18.400 1685.830 18.460 ;
        RECT 1690.110 18.400 1690.430 18.460 ;
      LAYER via ;
        RECT 1784.900 1687.800 1785.160 1688.060 ;
        RECT 1690.140 1686.440 1690.400 1686.700 ;
        RECT 1690.140 904.440 1690.400 904.700 ;
        RECT 1690.140 903.760 1690.400 904.020 ;
        RECT 1685.540 18.400 1685.800 18.660 ;
        RECT 1690.140 18.400 1690.400 18.660 ;
      LAYER met2 ;
        RECT 1784.825 1700.000 1785.105 1704.000 ;
        RECT 1784.960 1688.090 1785.100 1700.000 ;
        RECT 1784.900 1687.770 1785.160 1688.090 ;
        RECT 1690.140 1686.410 1690.400 1686.730 ;
        RECT 1690.200 904.730 1690.340 1686.410 ;
        RECT 1690.140 904.410 1690.400 904.730 ;
        RECT 1690.140 903.730 1690.400 904.050 ;
        RECT 1690.200 18.690 1690.340 903.730 ;
        RECT 1685.540 18.370 1685.800 18.690 ;
        RECT 1690.140 18.370 1690.400 18.690 ;
        RECT 1685.600 2.400 1685.740 18.370 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 60.080 724.430 60.140 ;
        RECT 1422.390 60.080 1422.710 60.140 ;
        RECT 724.110 59.940 1422.710 60.080 ;
        RECT 724.110 59.880 724.430 59.940 ;
        RECT 1422.390 59.880 1422.710 59.940 ;
      LAYER via ;
        RECT 724.140 59.880 724.400 60.140 ;
        RECT 1422.420 59.880 1422.680 60.140 ;
      LAYER met2 ;
        RECT 1421.425 1700.410 1421.705 1704.000 ;
        RECT 1421.425 1700.270 1422.620 1700.410 ;
        RECT 1421.425 1700.000 1421.705 1700.270 ;
        RECT 1422.480 60.170 1422.620 1700.270 ;
        RECT 724.140 59.850 724.400 60.170 ;
        RECT 1422.420 59.850 1422.680 60.170 ;
        RECT 724.200 3.130 724.340 59.850 ;
        RECT 722.360 2.990 724.340 3.130 ;
        RECT 722.360 2.400 722.500 2.990 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 1688.340 1704.230 1688.400 ;
        RECT 1791.770 1688.340 1792.090 1688.400 ;
        RECT 1703.910 1688.200 1792.090 1688.340 ;
        RECT 1703.910 1688.140 1704.230 1688.200 ;
        RECT 1791.770 1688.140 1792.090 1688.200 ;
      LAYER via ;
        RECT 1703.940 1688.140 1704.200 1688.400 ;
        RECT 1791.800 1688.140 1792.060 1688.400 ;
      LAYER met2 ;
        RECT 1791.725 1700.000 1792.005 1704.000 ;
        RECT 1791.860 1688.430 1792.000 1700.000 ;
        RECT 1703.940 1688.110 1704.200 1688.430 ;
        RECT 1791.800 1688.110 1792.060 1688.430 ;
        RECT 1704.000 24.380 1704.140 1688.110 ;
        RECT 1703.540 24.240 1704.140 24.380 ;
        RECT 1703.540 2.400 1703.680 24.240 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1724.610 1689.020 1724.930 1689.080 ;
        RECT 1798.670 1689.020 1798.990 1689.080 ;
        RECT 1724.610 1688.880 1798.990 1689.020 ;
        RECT 1724.610 1688.820 1724.930 1688.880 ;
        RECT 1798.670 1688.820 1798.990 1688.880 ;
        RECT 1721.390 20.640 1721.710 20.700 ;
        RECT 1724.610 20.640 1724.930 20.700 ;
        RECT 1721.390 20.500 1724.930 20.640 ;
        RECT 1721.390 20.440 1721.710 20.500 ;
        RECT 1724.610 20.440 1724.930 20.500 ;
      LAYER via ;
        RECT 1724.640 1688.820 1724.900 1689.080 ;
        RECT 1798.700 1688.820 1798.960 1689.080 ;
        RECT 1721.420 20.440 1721.680 20.700 ;
        RECT 1724.640 20.440 1724.900 20.700 ;
      LAYER met2 ;
        RECT 1798.625 1700.000 1798.905 1704.000 ;
        RECT 1798.760 1689.110 1798.900 1700.000 ;
        RECT 1724.640 1688.790 1724.900 1689.110 ;
        RECT 1798.700 1688.790 1798.960 1689.110 ;
        RECT 1724.700 20.730 1724.840 1688.790 ;
        RECT 1721.420 20.410 1721.680 20.730 ;
        RECT 1724.640 20.410 1724.900 20.730 ;
        RECT 1721.480 2.400 1721.620 20.410 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1764.245 1689.205 1764.415 1690.055 ;
      LAYER mcon ;
        RECT 1764.245 1689.885 1764.415 1690.055 ;
      LAYER met1 ;
        RECT 1745.310 1690.040 1745.630 1690.100 ;
        RECT 1764.185 1690.040 1764.475 1690.085 ;
        RECT 1745.310 1689.900 1764.475 1690.040 ;
        RECT 1745.310 1689.840 1745.630 1689.900 ;
        RECT 1764.185 1689.855 1764.475 1689.900 ;
        RECT 1805.110 1689.700 1805.430 1689.760 ;
        RECT 1776.220 1689.560 1805.430 1689.700 ;
        RECT 1764.185 1689.360 1764.475 1689.405 ;
        RECT 1776.220 1689.360 1776.360 1689.560 ;
        RECT 1805.110 1689.500 1805.430 1689.560 ;
        RECT 1764.185 1689.220 1776.360 1689.360 ;
        RECT 1764.185 1689.175 1764.475 1689.220 ;
        RECT 1739.330 17.920 1739.650 17.980 ;
        RECT 1745.310 17.920 1745.630 17.980 ;
        RECT 1739.330 17.780 1745.630 17.920 ;
        RECT 1739.330 17.720 1739.650 17.780 ;
        RECT 1745.310 17.720 1745.630 17.780 ;
      LAYER via ;
        RECT 1745.340 1689.840 1745.600 1690.100 ;
        RECT 1805.140 1689.500 1805.400 1689.760 ;
        RECT 1739.360 17.720 1739.620 17.980 ;
        RECT 1745.340 17.720 1745.600 17.980 ;
      LAYER met2 ;
        RECT 1805.065 1700.000 1805.345 1704.000 ;
        RECT 1745.340 1689.810 1745.600 1690.130 ;
        RECT 1745.400 18.010 1745.540 1689.810 ;
        RECT 1805.200 1689.790 1805.340 1700.000 ;
        RECT 1805.140 1689.470 1805.400 1689.790 ;
        RECT 1739.360 17.690 1739.620 18.010 ;
        RECT 1745.340 17.690 1745.600 18.010 ;
        RECT 1739.420 2.400 1739.560 17.690 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1775.745 1687.505 1775.915 1689.715 ;
      LAYER mcon ;
        RECT 1775.745 1689.545 1775.915 1689.715 ;
      LAYER met1 ;
        RECT 1759.110 1689.700 1759.430 1689.760 ;
        RECT 1775.685 1689.700 1775.975 1689.745 ;
        RECT 1759.110 1689.560 1775.975 1689.700 ;
        RECT 1759.110 1689.500 1759.430 1689.560 ;
        RECT 1775.685 1689.515 1775.975 1689.560 ;
        RECT 1775.685 1687.660 1775.975 1687.705 ;
        RECT 1812.010 1687.660 1812.330 1687.720 ;
        RECT 1775.685 1687.520 1812.330 1687.660 ;
        RECT 1775.685 1687.475 1775.975 1687.520 ;
        RECT 1812.010 1687.460 1812.330 1687.520 ;
        RECT 1756.810 17.580 1757.130 17.640 ;
        RECT 1759.110 17.580 1759.430 17.640 ;
        RECT 1756.810 17.440 1759.430 17.580 ;
        RECT 1756.810 17.380 1757.130 17.440 ;
        RECT 1759.110 17.380 1759.430 17.440 ;
      LAYER via ;
        RECT 1759.140 1689.500 1759.400 1689.760 ;
        RECT 1812.040 1687.460 1812.300 1687.720 ;
        RECT 1756.840 17.380 1757.100 17.640 ;
        RECT 1759.140 17.380 1759.400 17.640 ;
      LAYER met2 ;
        RECT 1811.965 1700.000 1812.245 1704.000 ;
        RECT 1759.140 1689.470 1759.400 1689.790 ;
        RECT 1759.200 17.670 1759.340 1689.470 ;
        RECT 1812.100 1687.750 1812.240 1700.000 ;
        RECT 1812.040 1687.430 1812.300 1687.750 ;
        RECT 1756.840 17.350 1757.100 17.670 ;
        RECT 1759.140 17.350 1759.400 17.670 ;
        RECT 1756.900 2.400 1757.040 17.350 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1779.810 1686.980 1780.130 1687.040 ;
        RECT 1818.910 1686.980 1819.230 1687.040 ;
        RECT 1779.810 1686.840 1819.230 1686.980 ;
        RECT 1779.810 1686.780 1780.130 1686.840 ;
        RECT 1818.910 1686.780 1819.230 1686.840 ;
        RECT 1774.750 17.580 1775.070 17.640 ;
        RECT 1779.810 17.580 1780.130 17.640 ;
        RECT 1774.750 17.440 1780.130 17.580 ;
        RECT 1774.750 17.380 1775.070 17.440 ;
        RECT 1779.810 17.380 1780.130 17.440 ;
      LAYER via ;
        RECT 1779.840 1686.780 1780.100 1687.040 ;
        RECT 1818.940 1686.780 1819.200 1687.040 ;
        RECT 1774.780 17.380 1775.040 17.640 ;
        RECT 1779.840 17.380 1780.100 17.640 ;
      LAYER met2 ;
        RECT 1818.865 1700.000 1819.145 1704.000 ;
        RECT 1819.000 1687.070 1819.140 1700.000 ;
        RECT 1779.840 1686.750 1780.100 1687.070 ;
        RECT 1818.940 1686.750 1819.200 1687.070 ;
        RECT 1779.900 17.670 1780.040 1686.750 ;
        RECT 1774.780 17.350 1775.040 17.670 ;
        RECT 1779.840 17.350 1780.100 17.670 ;
        RECT 1774.840 2.400 1774.980 17.350 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 1685.620 1793.930 1685.680 ;
        RECT 1825.350 1685.620 1825.670 1685.680 ;
        RECT 1793.610 1685.480 1825.670 1685.620 ;
        RECT 1793.610 1685.420 1793.930 1685.480 ;
        RECT 1825.350 1685.420 1825.670 1685.480 ;
        RECT 1792.690 2.960 1793.010 3.020 ;
        RECT 1793.610 2.960 1793.930 3.020 ;
        RECT 1792.690 2.820 1793.930 2.960 ;
        RECT 1792.690 2.760 1793.010 2.820 ;
        RECT 1793.610 2.760 1793.930 2.820 ;
      LAYER via ;
        RECT 1793.640 1685.420 1793.900 1685.680 ;
        RECT 1825.380 1685.420 1825.640 1685.680 ;
        RECT 1792.720 2.760 1792.980 3.020 ;
        RECT 1793.640 2.760 1793.900 3.020 ;
      LAYER met2 ;
        RECT 1825.305 1700.000 1825.585 1704.000 ;
        RECT 1825.440 1685.710 1825.580 1700.000 ;
        RECT 1793.640 1685.390 1793.900 1685.710 ;
        RECT 1825.380 1685.390 1825.640 1685.710 ;
        RECT 1793.700 3.050 1793.840 1685.390 ;
        RECT 1792.720 2.730 1792.980 3.050 ;
        RECT 1793.640 2.730 1793.900 3.050 ;
        RECT 1792.780 2.400 1792.920 2.730 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.310 1683.920 1814.630 1683.980 ;
        RECT 1832.250 1683.920 1832.570 1683.980 ;
        RECT 1814.310 1683.780 1832.570 1683.920 ;
        RECT 1814.310 1683.720 1814.630 1683.780 ;
        RECT 1832.250 1683.720 1832.570 1683.780 ;
        RECT 1810.630 20.640 1810.950 20.700 ;
        RECT 1814.310 20.640 1814.630 20.700 ;
        RECT 1810.630 20.500 1814.630 20.640 ;
        RECT 1810.630 20.440 1810.950 20.500 ;
        RECT 1814.310 20.440 1814.630 20.500 ;
      LAYER via ;
        RECT 1814.340 1683.720 1814.600 1683.980 ;
        RECT 1832.280 1683.720 1832.540 1683.980 ;
        RECT 1810.660 20.440 1810.920 20.700 ;
        RECT 1814.340 20.440 1814.600 20.700 ;
      LAYER met2 ;
        RECT 1832.205 1700.000 1832.485 1704.000 ;
        RECT 1832.340 1684.010 1832.480 1700.000 ;
        RECT 1814.340 1683.690 1814.600 1684.010 ;
        RECT 1832.280 1683.690 1832.540 1684.010 ;
        RECT 1814.400 20.730 1814.540 1683.690 ;
        RECT 1810.660 20.410 1810.920 20.730 ;
        RECT 1814.340 20.410 1814.600 20.730 ;
        RECT 1810.720 2.400 1810.860 20.410 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1834.550 1684.260 1834.870 1684.320 ;
        RECT 1839.150 1684.260 1839.470 1684.320 ;
        RECT 1834.550 1684.120 1839.470 1684.260 ;
        RECT 1834.550 1684.060 1834.870 1684.120 ;
        RECT 1839.150 1684.060 1839.470 1684.120 ;
        RECT 1828.570 16.560 1828.890 16.620 ;
        RECT 1834.550 16.560 1834.870 16.620 ;
        RECT 1828.570 16.420 1834.870 16.560 ;
        RECT 1828.570 16.360 1828.890 16.420 ;
        RECT 1834.550 16.360 1834.870 16.420 ;
      LAYER via ;
        RECT 1834.580 1684.060 1834.840 1684.320 ;
        RECT 1839.180 1684.060 1839.440 1684.320 ;
        RECT 1828.600 16.360 1828.860 16.620 ;
        RECT 1834.580 16.360 1834.840 16.620 ;
      LAYER met2 ;
        RECT 1839.105 1700.000 1839.385 1704.000 ;
        RECT 1839.240 1684.350 1839.380 1700.000 ;
        RECT 1834.580 1684.030 1834.840 1684.350 ;
        RECT 1839.180 1684.030 1839.440 1684.350 ;
        RECT 1834.640 16.650 1834.780 1684.030 ;
        RECT 1828.600 16.330 1828.860 16.650 ;
        RECT 1834.580 16.330 1834.840 16.650 ;
        RECT 1828.660 2.400 1828.800 16.330 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1842.830 20.640 1843.150 20.700 ;
        RECT 1846.050 20.640 1846.370 20.700 ;
        RECT 1842.830 20.500 1846.370 20.640 ;
        RECT 1842.830 20.440 1843.150 20.500 ;
        RECT 1846.050 20.440 1846.370 20.500 ;
      LAYER via ;
        RECT 1842.860 20.440 1843.120 20.700 ;
        RECT 1846.080 20.440 1846.340 20.700 ;
      LAYER met2 ;
        RECT 1845.545 1700.410 1845.825 1704.000 ;
        RECT 1844.300 1700.270 1845.825 1700.410 ;
        RECT 1844.300 1677.970 1844.440 1700.270 ;
        RECT 1845.545 1700.000 1845.825 1700.270 ;
        RECT 1842.920 1677.830 1844.440 1677.970 ;
        RECT 1842.920 20.730 1843.060 1677.830 ;
        RECT 1842.860 20.410 1843.120 20.730 ;
        RECT 1846.080 20.410 1846.340 20.730 ;
        RECT 1846.140 2.400 1846.280 20.410 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1852.490 1685.960 1852.810 1686.020 ;
        RECT 1863.530 1685.960 1863.850 1686.020 ;
        RECT 1852.490 1685.820 1863.850 1685.960 ;
        RECT 1852.490 1685.760 1852.810 1685.820 ;
        RECT 1863.530 1685.760 1863.850 1685.820 ;
      LAYER via ;
        RECT 1852.520 1685.760 1852.780 1686.020 ;
        RECT 1863.560 1685.760 1863.820 1686.020 ;
      LAYER met2 ;
        RECT 1852.445 1700.000 1852.725 1704.000 ;
        RECT 1852.580 1686.050 1852.720 1700.000 ;
        RECT 1852.520 1685.730 1852.780 1686.050 ;
        RECT 1863.560 1685.730 1863.820 1686.050 ;
        RECT 1863.620 17.410 1863.760 1685.730 ;
        RECT 1863.620 17.270 1864.220 17.410 ;
        RECT 1864.080 2.400 1864.220 17.270 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 744.810 60.420 745.130 60.480 ;
        RECT 1429.750 60.420 1430.070 60.480 ;
        RECT 744.810 60.280 1430.070 60.420 ;
        RECT 744.810 60.220 745.130 60.280 ;
        RECT 1429.750 60.220 1430.070 60.280 ;
        RECT 740.210 2.960 740.530 3.020 ;
        RECT 744.810 2.960 745.130 3.020 ;
        RECT 740.210 2.820 745.130 2.960 ;
        RECT 740.210 2.760 740.530 2.820 ;
        RECT 744.810 2.760 745.130 2.820 ;
      LAYER via ;
        RECT 744.840 60.220 745.100 60.480 ;
        RECT 1429.780 60.220 1430.040 60.480 ;
        RECT 740.240 2.760 740.500 3.020 ;
        RECT 744.840 2.760 745.100 3.020 ;
      LAYER met2 ;
        RECT 1428.325 1700.410 1428.605 1704.000 ;
        RECT 1428.325 1700.270 1429.980 1700.410 ;
        RECT 1428.325 1700.000 1428.605 1700.270 ;
        RECT 1429.840 60.510 1429.980 1700.270 ;
        RECT 744.840 60.190 745.100 60.510 ;
        RECT 1429.780 60.190 1430.040 60.510 ;
        RECT 744.900 3.050 745.040 60.190 ;
        RECT 740.240 2.730 740.500 3.050 ;
        RECT 744.840 2.730 745.100 3.050 ;
        RECT 740.300 2.400 740.440 2.730 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1858.930 1685.280 1859.250 1685.340 ;
        RECT 1878.250 1685.280 1878.570 1685.340 ;
        RECT 1858.930 1685.140 1878.570 1685.280 ;
        RECT 1858.930 1685.080 1859.250 1685.140 ;
        RECT 1878.250 1685.080 1878.570 1685.140 ;
      LAYER via ;
        RECT 1858.960 1685.080 1859.220 1685.340 ;
        RECT 1878.280 1685.080 1878.540 1685.340 ;
      LAYER met2 ;
        RECT 1858.885 1700.000 1859.165 1704.000 ;
        RECT 1859.020 1685.370 1859.160 1700.000 ;
        RECT 1858.960 1685.050 1859.220 1685.370 ;
        RECT 1878.280 1685.050 1878.540 1685.370 ;
        RECT 1878.340 16.730 1878.480 1685.050 ;
        RECT 1878.340 16.590 1882.160 16.730 ;
        RECT 1882.020 2.400 1882.160 16.590 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1865.830 1687.320 1866.150 1687.380 ;
        RECT 1865.830 1687.180 1882.620 1687.320 ;
        RECT 1865.830 1687.120 1866.150 1687.180 ;
        RECT 1882.480 1686.980 1882.620 1687.180 ;
        RECT 1898.030 1686.980 1898.350 1687.040 ;
        RECT 1882.480 1686.840 1898.350 1686.980 ;
        RECT 1898.030 1686.780 1898.350 1686.840 ;
        RECT 1898.030 2.960 1898.350 3.020 ;
        RECT 1899.870 2.960 1900.190 3.020 ;
        RECT 1898.030 2.820 1900.190 2.960 ;
        RECT 1898.030 2.760 1898.350 2.820 ;
        RECT 1899.870 2.760 1900.190 2.820 ;
      LAYER via ;
        RECT 1865.860 1687.120 1866.120 1687.380 ;
        RECT 1898.060 1686.780 1898.320 1687.040 ;
        RECT 1898.060 2.760 1898.320 3.020 ;
        RECT 1899.900 2.760 1900.160 3.020 ;
      LAYER met2 ;
        RECT 1865.785 1700.000 1866.065 1704.000 ;
        RECT 1865.920 1687.410 1866.060 1700.000 ;
        RECT 1865.860 1687.090 1866.120 1687.410 ;
        RECT 1898.060 1686.750 1898.320 1687.070 ;
        RECT 1898.120 3.050 1898.260 1686.750 ;
        RECT 1898.060 2.730 1898.320 3.050 ;
        RECT 1899.900 2.730 1900.160 3.050 ;
        RECT 1899.960 2.400 1900.100 2.730 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1872.730 1689.020 1873.050 1689.080 ;
        RECT 1880.090 1689.020 1880.410 1689.080 ;
        RECT 1872.730 1688.880 1880.410 1689.020 ;
        RECT 1872.730 1688.820 1873.050 1688.880 ;
        RECT 1880.090 1688.820 1880.410 1688.880 ;
        RECT 1880.090 19.280 1880.410 19.340 ;
        RECT 1917.350 19.280 1917.670 19.340 ;
        RECT 1880.090 19.140 1917.670 19.280 ;
        RECT 1880.090 19.080 1880.410 19.140 ;
        RECT 1917.350 19.080 1917.670 19.140 ;
      LAYER via ;
        RECT 1872.760 1688.820 1873.020 1689.080 ;
        RECT 1880.120 1688.820 1880.380 1689.080 ;
        RECT 1880.120 19.080 1880.380 19.340 ;
        RECT 1917.380 19.080 1917.640 19.340 ;
      LAYER met2 ;
        RECT 1872.685 1700.000 1872.965 1704.000 ;
        RECT 1872.820 1689.110 1872.960 1700.000 ;
        RECT 1872.760 1688.790 1873.020 1689.110 ;
        RECT 1880.120 1688.790 1880.380 1689.110 ;
        RECT 1880.180 19.370 1880.320 1688.790 ;
        RECT 1880.120 19.050 1880.380 19.370 ;
        RECT 1917.380 19.050 1917.640 19.370 ;
        RECT 1917.440 16.050 1917.580 19.050 ;
        RECT 1917.440 15.910 1918.040 16.050 ;
        RECT 1917.900 2.400 1918.040 15.910 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1879.170 1688.340 1879.490 1688.400 ;
        RECT 1886.990 1688.340 1887.310 1688.400 ;
        RECT 1879.170 1688.200 1887.310 1688.340 ;
        RECT 1879.170 1688.140 1879.490 1688.200 ;
        RECT 1886.990 1688.140 1887.310 1688.200 ;
        RECT 1886.990 18.260 1887.310 18.320 ;
        RECT 1935.290 18.260 1935.610 18.320 ;
        RECT 1886.990 18.120 1935.610 18.260 ;
        RECT 1886.990 18.060 1887.310 18.120 ;
        RECT 1935.290 18.060 1935.610 18.120 ;
      LAYER via ;
        RECT 1879.200 1688.140 1879.460 1688.400 ;
        RECT 1887.020 1688.140 1887.280 1688.400 ;
        RECT 1887.020 18.060 1887.280 18.320 ;
        RECT 1935.320 18.060 1935.580 18.320 ;
      LAYER met2 ;
        RECT 1879.125 1700.000 1879.405 1704.000 ;
        RECT 1879.260 1688.430 1879.400 1700.000 ;
        RECT 1879.200 1688.110 1879.460 1688.430 ;
        RECT 1887.020 1688.110 1887.280 1688.430 ;
        RECT 1887.080 18.350 1887.220 1688.110 ;
        RECT 1887.020 18.030 1887.280 18.350 ;
        RECT 1935.320 18.030 1935.580 18.350 ;
        RECT 1935.380 2.400 1935.520 18.030 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1935.825 16.745 1935.995 17.595 ;
      LAYER mcon ;
        RECT 1935.825 17.425 1935.995 17.595 ;
      LAYER met1 ;
        RECT 1886.070 1688.680 1886.390 1688.740 ;
        RECT 1889.750 1688.680 1890.070 1688.740 ;
        RECT 1886.070 1688.540 1890.070 1688.680 ;
        RECT 1886.070 1688.480 1886.390 1688.540 ;
        RECT 1889.750 1688.480 1890.070 1688.540 ;
        RECT 1889.750 17.580 1890.070 17.640 ;
        RECT 1935.765 17.580 1936.055 17.625 ;
        RECT 1889.750 17.440 1936.055 17.580 ;
        RECT 1889.750 17.380 1890.070 17.440 ;
        RECT 1935.765 17.395 1936.055 17.440 ;
        RECT 1935.765 16.900 1936.055 16.945 ;
        RECT 1953.230 16.900 1953.550 16.960 ;
        RECT 1935.765 16.760 1953.550 16.900 ;
        RECT 1935.765 16.715 1936.055 16.760 ;
        RECT 1953.230 16.700 1953.550 16.760 ;
      LAYER via ;
        RECT 1886.100 1688.480 1886.360 1688.740 ;
        RECT 1889.780 1688.480 1890.040 1688.740 ;
        RECT 1889.780 17.380 1890.040 17.640 ;
        RECT 1953.260 16.700 1953.520 16.960 ;
      LAYER met2 ;
        RECT 1886.025 1700.000 1886.305 1704.000 ;
        RECT 1886.160 1688.770 1886.300 1700.000 ;
        RECT 1886.100 1688.450 1886.360 1688.770 ;
        RECT 1889.780 1688.450 1890.040 1688.770 ;
        RECT 1889.840 17.670 1889.980 1688.450 ;
        RECT 1889.780 17.350 1890.040 17.670 ;
        RECT 1953.260 16.670 1953.520 16.990 ;
        RECT 1953.320 2.400 1953.460 16.670 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1892.970 1688.340 1893.290 1688.400 ;
        RECT 1900.790 1688.340 1901.110 1688.400 ;
        RECT 1892.970 1688.200 1901.110 1688.340 ;
        RECT 1892.970 1688.140 1893.290 1688.200 ;
        RECT 1900.790 1688.140 1901.110 1688.200 ;
        RECT 1900.790 17.240 1901.110 17.300 ;
        RECT 1971.170 17.240 1971.490 17.300 ;
        RECT 1900.790 17.100 1971.490 17.240 ;
        RECT 1900.790 17.040 1901.110 17.100 ;
        RECT 1971.170 17.040 1971.490 17.100 ;
      LAYER via ;
        RECT 1893.000 1688.140 1893.260 1688.400 ;
        RECT 1900.820 1688.140 1901.080 1688.400 ;
        RECT 1900.820 17.040 1901.080 17.300 ;
        RECT 1971.200 17.040 1971.460 17.300 ;
      LAYER met2 ;
        RECT 1892.925 1700.000 1893.205 1704.000 ;
        RECT 1893.060 1688.430 1893.200 1700.000 ;
        RECT 1893.000 1688.110 1893.260 1688.430 ;
        RECT 1900.820 1688.110 1901.080 1688.430 ;
        RECT 1900.880 17.330 1901.020 1688.110 ;
        RECT 1900.820 17.010 1901.080 17.330 ;
        RECT 1971.200 17.010 1971.460 17.330 ;
        RECT 1971.260 2.400 1971.400 17.010 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1899.410 1688.680 1899.730 1688.740 ;
        RECT 1904.010 1688.680 1904.330 1688.740 ;
        RECT 1899.410 1688.540 1904.330 1688.680 ;
        RECT 1899.410 1688.480 1899.730 1688.540 ;
        RECT 1904.010 1688.480 1904.330 1688.540 ;
        RECT 1904.010 15.200 1904.330 15.260 ;
        RECT 1989.110 15.200 1989.430 15.260 ;
        RECT 1904.010 15.060 1989.430 15.200 ;
        RECT 1904.010 15.000 1904.330 15.060 ;
        RECT 1989.110 15.000 1989.430 15.060 ;
      LAYER via ;
        RECT 1899.440 1688.480 1899.700 1688.740 ;
        RECT 1904.040 1688.480 1904.300 1688.740 ;
        RECT 1904.040 15.000 1904.300 15.260 ;
        RECT 1989.140 15.000 1989.400 15.260 ;
      LAYER met2 ;
        RECT 1899.365 1700.000 1899.645 1704.000 ;
        RECT 1899.500 1688.770 1899.640 1700.000 ;
        RECT 1899.440 1688.450 1899.700 1688.770 ;
        RECT 1904.040 1688.450 1904.300 1688.770 ;
        RECT 1904.100 15.290 1904.240 1688.450 ;
        RECT 1904.040 14.970 1904.300 15.290 ;
        RECT 1989.140 14.970 1989.400 15.290 ;
        RECT 1989.200 2.400 1989.340 14.970 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1906.310 1688.680 1906.630 1688.740 ;
        RECT 1910.910 1688.680 1911.230 1688.740 ;
        RECT 1906.310 1688.540 1911.230 1688.680 ;
        RECT 1906.310 1688.480 1906.630 1688.540 ;
        RECT 1910.910 1688.480 1911.230 1688.540 ;
        RECT 1910.910 15.540 1911.230 15.600 ;
        RECT 2006.590 15.540 2006.910 15.600 ;
        RECT 1910.910 15.400 2006.910 15.540 ;
        RECT 1910.910 15.340 1911.230 15.400 ;
        RECT 2006.590 15.340 2006.910 15.400 ;
      LAYER via ;
        RECT 1906.340 1688.480 1906.600 1688.740 ;
        RECT 1910.940 1688.480 1911.200 1688.740 ;
        RECT 1910.940 15.340 1911.200 15.600 ;
        RECT 2006.620 15.340 2006.880 15.600 ;
      LAYER met2 ;
        RECT 1906.265 1700.000 1906.545 1704.000 ;
        RECT 1906.400 1688.770 1906.540 1700.000 ;
        RECT 1906.340 1688.450 1906.600 1688.770 ;
        RECT 1910.940 1688.450 1911.200 1688.770 ;
        RECT 1911.000 15.630 1911.140 1688.450 ;
        RECT 1910.940 15.310 1911.200 15.630 ;
        RECT 2006.620 15.310 2006.880 15.630 ;
        RECT 2006.680 2.400 2006.820 15.310 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1917.885 1688.865 1918.055 1690.055 ;
      LAYER mcon ;
        RECT 1917.885 1689.885 1918.055 1690.055 ;
      LAYER met1 ;
        RECT 1917.825 1690.040 1918.115 1690.085 ;
        RECT 1917.825 1689.900 1942.420 1690.040 ;
        RECT 1917.825 1689.855 1918.115 1689.900 ;
        RECT 1942.280 1689.700 1942.420 1689.900 ;
        RECT 1969.790 1689.700 1970.110 1689.760 ;
        RECT 1942.280 1689.560 1970.110 1689.700 ;
        RECT 1969.790 1689.500 1970.110 1689.560 ;
        RECT 1913.210 1689.020 1913.530 1689.080 ;
        RECT 1917.825 1689.020 1918.115 1689.065 ;
        RECT 1913.210 1688.880 1918.115 1689.020 ;
        RECT 1913.210 1688.820 1913.530 1688.880 ;
        RECT 1917.825 1688.835 1918.115 1688.880 ;
        RECT 1969.790 14.180 1970.110 14.240 ;
        RECT 2024.530 14.180 2024.850 14.240 ;
        RECT 1969.790 14.040 2024.850 14.180 ;
        RECT 1969.790 13.980 1970.110 14.040 ;
        RECT 2024.530 13.980 2024.850 14.040 ;
      LAYER via ;
        RECT 1969.820 1689.500 1970.080 1689.760 ;
        RECT 1913.240 1688.820 1913.500 1689.080 ;
        RECT 1969.820 13.980 1970.080 14.240 ;
        RECT 2024.560 13.980 2024.820 14.240 ;
      LAYER met2 ;
        RECT 1913.165 1700.000 1913.445 1704.000 ;
        RECT 1913.300 1689.110 1913.440 1700.000 ;
        RECT 1969.820 1689.470 1970.080 1689.790 ;
        RECT 1913.240 1688.790 1913.500 1689.110 ;
        RECT 1969.880 14.270 1970.020 1689.470 ;
        RECT 1969.820 13.950 1970.080 14.270 ;
        RECT 2024.560 13.950 2024.820 14.270 ;
        RECT 2024.620 2.400 2024.760 13.950 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1941.805 16.065 1941.975 19.635 ;
      LAYER mcon ;
        RECT 1941.805 19.465 1941.975 19.635 ;
      LAYER met1 ;
        RECT 1919.650 1688.680 1919.970 1688.740 ;
        RECT 1924.710 1688.680 1925.030 1688.740 ;
        RECT 1919.650 1688.540 1925.030 1688.680 ;
        RECT 1919.650 1688.480 1919.970 1688.540 ;
        RECT 1924.710 1688.480 1925.030 1688.540 ;
        RECT 1924.710 19.620 1925.030 19.680 ;
        RECT 1941.745 19.620 1942.035 19.665 ;
        RECT 1924.710 19.480 1942.035 19.620 ;
        RECT 1924.710 19.420 1925.030 19.480 ;
        RECT 1941.745 19.435 1942.035 19.480 ;
        RECT 1941.745 16.220 1942.035 16.265 ;
        RECT 2042.470 16.220 2042.790 16.280 ;
        RECT 1941.745 16.080 2042.790 16.220 ;
        RECT 1941.745 16.035 1942.035 16.080 ;
        RECT 2042.470 16.020 2042.790 16.080 ;
      LAYER via ;
        RECT 1919.680 1688.480 1919.940 1688.740 ;
        RECT 1924.740 1688.480 1925.000 1688.740 ;
        RECT 1924.740 19.420 1925.000 19.680 ;
        RECT 2042.500 16.020 2042.760 16.280 ;
      LAYER met2 ;
        RECT 1919.605 1700.000 1919.885 1704.000 ;
        RECT 1919.740 1688.770 1919.880 1700.000 ;
        RECT 1919.680 1688.450 1919.940 1688.770 ;
        RECT 1924.740 1688.450 1925.000 1688.770 ;
        RECT 1924.800 19.710 1924.940 1688.450 ;
        RECT 1924.740 19.390 1925.000 19.710 ;
        RECT 2042.500 15.990 2042.760 16.310 ;
        RECT 2042.560 2.400 2042.700 15.990 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1429.290 1678.480 1429.610 1678.540 ;
        RECT 1433.430 1678.480 1433.750 1678.540 ;
        RECT 1429.290 1678.340 1433.750 1678.480 ;
        RECT 1429.290 1678.280 1429.610 1678.340 ;
        RECT 1433.430 1678.280 1433.750 1678.340 ;
        RECT 758.610 60.760 758.930 60.820 ;
        RECT 1429.290 60.760 1429.610 60.820 ;
        RECT 758.610 60.620 1429.610 60.760 ;
        RECT 758.610 60.560 758.930 60.620 ;
        RECT 1429.290 60.560 1429.610 60.620 ;
        RECT 757.690 2.960 758.010 3.020 ;
        RECT 758.610 2.960 758.930 3.020 ;
        RECT 757.690 2.820 758.930 2.960 ;
        RECT 757.690 2.760 758.010 2.820 ;
        RECT 758.610 2.760 758.930 2.820 ;
      LAYER via ;
        RECT 1429.320 1678.280 1429.580 1678.540 ;
        RECT 1433.460 1678.280 1433.720 1678.540 ;
        RECT 758.640 60.560 758.900 60.820 ;
        RECT 1429.320 60.560 1429.580 60.820 ;
        RECT 757.720 2.760 757.980 3.020 ;
        RECT 758.640 2.760 758.900 3.020 ;
      LAYER met2 ;
        RECT 1434.765 1700.410 1435.045 1704.000 ;
        RECT 1433.520 1700.270 1435.045 1700.410 ;
        RECT 1433.520 1678.570 1433.660 1700.270 ;
        RECT 1434.765 1700.000 1435.045 1700.270 ;
        RECT 1429.320 1678.250 1429.580 1678.570 ;
        RECT 1433.460 1678.250 1433.720 1678.570 ;
        RECT 1429.380 60.850 1429.520 1678.250 ;
        RECT 758.640 60.530 758.900 60.850 ;
        RECT 1429.320 60.530 1429.580 60.850 ;
        RECT 758.700 3.050 758.840 60.530 ;
        RECT 757.720 2.730 757.980 3.050 ;
        RECT 758.640 2.730 758.900 3.050 ;
        RECT 757.780 2.400 757.920 2.730 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1966.185 1686.485 1966.355 1687.675 ;
      LAYER mcon ;
        RECT 1966.185 1687.505 1966.355 1687.675 ;
      LAYER met1 ;
        RECT 1966.125 1687.660 1966.415 1687.705 ;
        RECT 2025.450 1687.660 2025.770 1687.720 ;
        RECT 1966.125 1687.520 2025.770 1687.660 ;
        RECT 1966.125 1687.475 1966.415 1687.520 ;
        RECT 2025.450 1687.460 2025.770 1687.520 ;
        RECT 1926.550 1686.640 1926.870 1686.700 ;
        RECT 1966.125 1686.640 1966.415 1686.685 ;
        RECT 1926.550 1686.500 1966.415 1686.640 ;
        RECT 1926.550 1686.440 1926.870 1686.500 ;
        RECT 1966.125 1686.455 1966.415 1686.500 ;
        RECT 2025.450 15.540 2025.770 15.600 ;
        RECT 2060.410 15.540 2060.730 15.600 ;
        RECT 2025.450 15.400 2060.730 15.540 ;
        RECT 2025.450 15.340 2025.770 15.400 ;
        RECT 2060.410 15.340 2060.730 15.400 ;
      LAYER via ;
        RECT 2025.480 1687.460 2025.740 1687.720 ;
        RECT 1926.580 1686.440 1926.840 1686.700 ;
        RECT 2025.480 15.340 2025.740 15.600 ;
        RECT 2060.440 15.340 2060.700 15.600 ;
      LAYER met2 ;
        RECT 1926.505 1700.000 1926.785 1704.000 ;
        RECT 1926.640 1686.730 1926.780 1700.000 ;
        RECT 2025.480 1687.430 2025.740 1687.750 ;
        RECT 1926.580 1686.410 1926.840 1686.730 ;
        RECT 2025.540 15.630 2025.680 1687.430 ;
        RECT 2025.480 15.310 2025.740 15.630 ;
        RECT 2060.440 15.310 2060.700 15.630 ;
        RECT 2060.500 2.400 2060.640 15.310 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1932.990 1688.000 1933.310 1688.060 ;
        RECT 1937.590 1688.000 1937.910 1688.060 ;
        RECT 1932.990 1687.860 1937.910 1688.000 ;
        RECT 1932.990 1687.800 1933.310 1687.860 ;
        RECT 1937.590 1687.800 1937.910 1687.860 ;
        RECT 1937.590 23.360 1937.910 23.420 ;
        RECT 2078.350 23.360 2078.670 23.420 ;
        RECT 1937.590 23.220 2078.670 23.360 ;
        RECT 1937.590 23.160 1937.910 23.220 ;
        RECT 2078.350 23.160 2078.670 23.220 ;
      LAYER via ;
        RECT 1933.020 1687.800 1933.280 1688.060 ;
        RECT 1937.620 1687.800 1937.880 1688.060 ;
        RECT 1937.620 23.160 1937.880 23.420 ;
        RECT 2078.380 23.160 2078.640 23.420 ;
      LAYER met2 ;
        RECT 1932.945 1700.000 1933.225 1704.000 ;
        RECT 1933.080 1688.090 1933.220 1700.000 ;
        RECT 1933.020 1687.770 1933.280 1688.090 ;
        RECT 1937.620 1687.770 1937.880 1688.090 ;
        RECT 1937.680 23.450 1937.820 1687.770 ;
        RECT 1937.620 23.130 1937.880 23.450 ;
        RECT 2078.380 23.130 2078.640 23.450 ;
        RECT 2078.440 2.400 2078.580 23.130 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2038.790 1688.000 2039.110 1688.060 ;
        RECT 1965.740 1687.860 2039.110 1688.000 ;
        RECT 1939.890 1687.660 1940.210 1687.720 ;
        RECT 1965.740 1687.660 1965.880 1687.860 ;
        RECT 2038.790 1687.800 2039.110 1687.860 ;
        RECT 1939.890 1687.520 1965.880 1687.660 ;
        RECT 1939.890 1687.460 1940.210 1687.520 ;
        RECT 2038.790 16.560 2039.110 16.620 ;
        RECT 2095.830 16.560 2096.150 16.620 ;
        RECT 2038.790 16.420 2096.150 16.560 ;
        RECT 2038.790 16.360 2039.110 16.420 ;
        RECT 2095.830 16.360 2096.150 16.420 ;
      LAYER via ;
        RECT 1939.920 1687.460 1940.180 1687.720 ;
        RECT 2038.820 1687.800 2039.080 1688.060 ;
        RECT 2038.820 16.360 2039.080 16.620 ;
        RECT 2095.860 16.360 2096.120 16.620 ;
      LAYER met2 ;
        RECT 1939.845 1700.000 1940.125 1704.000 ;
        RECT 1939.980 1687.750 1940.120 1700.000 ;
        RECT 2038.820 1687.770 2039.080 1688.090 ;
        RECT 1939.920 1687.430 1940.180 1687.750 ;
        RECT 2038.880 16.650 2039.020 1687.770 ;
        RECT 2038.820 16.330 2039.080 16.650 ;
        RECT 2095.860 16.330 2096.120 16.650 ;
        RECT 2095.920 2.400 2096.060 16.330 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1946.790 1688.680 1947.110 1688.740 ;
        RECT 1952.310 1688.680 1952.630 1688.740 ;
        RECT 1946.790 1688.540 1952.630 1688.680 ;
        RECT 1946.790 1688.480 1947.110 1688.540 ;
        RECT 1952.310 1688.480 1952.630 1688.540 ;
        RECT 1952.310 23.700 1952.630 23.760 ;
        RECT 2113.770 23.700 2114.090 23.760 ;
        RECT 1952.310 23.560 2114.090 23.700 ;
        RECT 1952.310 23.500 1952.630 23.560 ;
        RECT 2113.770 23.500 2114.090 23.560 ;
      LAYER via ;
        RECT 1946.820 1688.480 1947.080 1688.740 ;
        RECT 1952.340 1688.480 1952.600 1688.740 ;
        RECT 1952.340 23.500 1952.600 23.760 ;
        RECT 2113.800 23.500 2114.060 23.760 ;
      LAYER met2 ;
        RECT 1946.745 1700.000 1947.025 1704.000 ;
        RECT 1946.880 1688.770 1947.020 1700.000 ;
        RECT 1946.820 1688.450 1947.080 1688.770 ;
        RECT 1952.340 1688.450 1952.600 1688.770 ;
        RECT 1952.400 23.790 1952.540 1688.450 ;
        RECT 1952.340 23.470 1952.600 23.790 ;
        RECT 2113.800 23.470 2114.060 23.790 ;
        RECT 2113.860 2.400 2114.000 23.470 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1953.230 1688.000 1953.550 1688.060 ;
        RECT 1958.290 1688.000 1958.610 1688.060 ;
        RECT 1953.230 1687.860 1958.610 1688.000 ;
        RECT 1953.230 1687.800 1953.550 1687.860 ;
        RECT 1958.290 1687.800 1958.610 1687.860 ;
        RECT 1958.290 27.100 1958.610 27.160 ;
        RECT 2131.710 27.100 2132.030 27.160 ;
        RECT 1958.290 26.960 2132.030 27.100 ;
        RECT 1958.290 26.900 1958.610 26.960 ;
        RECT 2131.710 26.900 2132.030 26.960 ;
      LAYER via ;
        RECT 1953.260 1687.800 1953.520 1688.060 ;
        RECT 1958.320 1687.800 1958.580 1688.060 ;
        RECT 1958.320 26.900 1958.580 27.160 ;
        RECT 2131.740 26.900 2132.000 27.160 ;
      LAYER met2 ;
        RECT 1953.185 1700.000 1953.465 1704.000 ;
        RECT 1953.320 1688.090 1953.460 1700.000 ;
        RECT 1953.260 1687.770 1953.520 1688.090 ;
        RECT 1958.320 1687.770 1958.580 1688.090 ;
        RECT 1958.380 27.190 1958.520 1687.770 ;
        RECT 1958.320 26.870 1958.580 27.190 ;
        RECT 2131.740 26.870 2132.000 27.190 ;
        RECT 2131.800 2.400 2131.940 26.870 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1960.130 1688.000 1960.450 1688.060 ;
        RECT 1965.190 1688.000 1965.510 1688.060 ;
        RECT 1960.130 1687.860 1965.510 1688.000 ;
        RECT 1960.130 1687.800 1960.450 1687.860 ;
        RECT 1965.190 1687.800 1965.510 1687.860 ;
        RECT 1965.190 26.760 1965.510 26.820 ;
        RECT 2149.650 26.760 2149.970 26.820 ;
        RECT 1965.190 26.620 2149.970 26.760 ;
        RECT 1965.190 26.560 1965.510 26.620 ;
        RECT 2149.650 26.560 2149.970 26.620 ;
      LAYER via ;
        RECT 1960.160 1687.800 1960.420 1688.060 ;
        RECT 1965.220 1687.800 1965.480 1688.060 ;
        RECT 1965.220 26.560 1965.480 26.820 ;
        RECT 2149.680 26.560 2149.940 26.820 ;
      LAYER met2 ;
        RECT 1960.085 1700.000 1960.365 1704.000 ;
        RECT 1960.220 1688.090 1960.360 1700.000 ;
        RECT 1960.160 1687.770 1960.420 1688.090 ;
        RECT 1965.220 1687.770 1965.480 1688.090 ;
        RECT 1965.280 26.850 1965.420 1687.770 ;
        RECT 1965.220 26.530 1965.480 26.850 ;
        RECT 2149.680 26.530 2149.940 26.850 ;
        RECT 2149.740 2.400 2149.880 26.530 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1967.030 1685.620 1967.350 1685.680 ;
        RECT 1972.550 1685.620 1972.870 1685.680 ;
        RECT 1967.030 1685.480 1972.870 1685.620 ;
        RECT 1967.030 1685.420 1967.350 1685.480 ;
        RECT 1972.550 1685.420 1972.870 1685.480 ;
        RECT 1972.550 26.420 1972.870 26.480 ;
        RECT 2167.590 26.420 2167.910 26.480 ;
        RECT 1972.550 26.280 2167.910 26.420 ;
        RECT 1972.550 26.220 1972.870 26.280 ;
        RECT 2167.590 26.220 2167.910 26.280 ;
      LAYER via ;
        RECT 1967.060 1685.420 1967.320 1685.680 ;
        RECT 1972.580 1685.420 1972.840 1685.680 ;
        RECT 1972.580 26.220 1972.840 26.480 ;
        RECT 2167.620 26.220 2167.880 26.480 ;
      LAYER met2 ;
        RECT 1966.985 1700.000 1967.265 1704.000 ;
        RECT 1967.120 1685.710 1967.260 1700.000 ;
        RECT 1967.060 1685.390 1967.320 1685.710 ;
        RECT 1972.580 1685.390 1972.840 1685.710 ;
        RECT 1972.640 26.510 1972.780 1685.390 ;
        RECT 1972.580 26.190 1972.840 26.510 ;
        RECT 2167.620 26.190 2167.880 26.510 ;
        RECT 2167.680 2.400 2167.820 26.190 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.470 1687.320 1973.790 1687.380 ;
        RECT 1978.990 1687.320 1979.310 1687.380 ;
        RECT 1973.470 1687.180 1979.310 1687.320 ;
        RECT 1973.470 1687.120 1973.790 1687.180 ;
        RECT 1978.990 1687.120 1979.310 1687.180 ;
        RECT 1978.990 25.740 1979.310 25.800 ;
        RECT 2185.070 25.740 2185.390 25.800 ;
        RECT 1978.990 25.600 2185.390 25.740 ;
        RECT 1978.990 25.540 1979.310 25.600 ;
        RECT 2185.070 25.540 2185.390 25.600 ;
      LAYER via ;
        RECT 1973.500 1687.120 1973.760 1687.380 ;
        RECT 1979.020 1687.120 1979.280 1687.380 ;
        RECT 1979.020 25.540 1979.280 25.800 ;
        RECT 2185.100 25.540 2185.360 25.800 ;
      LAYER met2 ;
        RECT 1973.425 1700.000 1973.705 1704.000 ;
        RECT 1973.560 1687.410 1973.700 1700.000 ;
        RECT 1973.500 1687.090 1973.760 1687.410 ;
        RECT 1979.020 1687.090 1979.280 1687.410 ;
        RECT 1979.080 25.830 1979.220 1687.090 ;
        RECT 1979.020 25.510 1979.280 25.830 ;
        RECT 2185.100 25.510 2185.360 25.830 ;
        RECT 2185.160 2.400 2185.300 25.510 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1980.370 1688.340 1980.690 1688.400 ;
        RECT 1986.810 1688.340 1987.130 1688.400 ;
        RECT 1980.370 1688.200 1987.130 1688.340 ;
        RECT 1980.370 1688.140 1980.690 1688.200 ;
        RECT 1986.810 1688.140 1987.130 1688.200 ;
        RECT 1986.810 25.060 1987.130 25.120 ;
        RECT 2203.010 25.060 2203.330 25.120 ;
        RECT 1986.810 24.920 2203.330 25.060 ;
        RECT 1986.810 24.860 1987.130 24.920 ;
        RECT 2203.010 24.860 2203.330 24.920 ;
      LAYER via ;
        RECT 1980.400 1688.140 1980.660 1688.400 ;
        RECT 1986.840 1688.140 1987.100 1688.400 ;
        RECT 1986.840 24.860 1987.100 25.120 ;
        RECT 2203.040 24.860 2203.300 25.120 ;
      LAYER met2 ;
        RECT 1980.325 1700.000 1980.605 1704.000 ;
        RECT 1980.460 1688.430 1980.600 1700.000 ;
        RECT 1980.400 1688.110 1980.660 1688.430 ;
        RECT 1986.840 1688.110 1987.100 1688.430 ;
        RECT 1986.900 25.150 1987.040 1688.110 ;
        RECT 1986.840 24.830 1987.100 25.150 ;
        RECT 2203.040 24.830 2203.300 25.150 ;
        RECT 2203.100 2.400 2203.240 24.830 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1987.270 1688.340 1987.590 1688.400 ;
        RECT 1993.250 1688.340 1993.570 1688.400 ;
        RECT 1987.270 1688.200 1993.570 1688.340 ;
        RECT 1987.270 1688.140 1987.590 1688.200 ;
        RECT 1993.250 1688.140 1993.570 1688.200 ;
        RECT 1993.250 24.720 1993.570 24.780 ;
        RECT 2220.950 24.720 2221.270 24.780 ;
        RECT 1993.250 24.580 2221.270 24.720 ;
        RECT 1993.250 24.520 1993.570 24.580 ;
        RECT 2220.950 24.520 2221.270 24.580 ;
      LAYER via ;
        RECT 1987.300 1688.140 1987.560 1688.400 ;
        RECT 1993.280 1688.140 1993.540 1688.400 ;
        RECT 1993.280 24.520 1993.540 24.780 ;
        RECT 2220.980 24.520 2221.240 24.780 ;
      LAYER met2 ;
        RECT 1987.225 1700.000 1987.505 1704.000 ;
        RECT 1987.360 1688.430 1987.500 1700.000 ;
        RECT 1987.300 1688.110 1987.560 1688.430 ;
        RECT 1993.280 1688.110 1993.540 1688.430 ;
        RECT 1993.340 24.810 1993.480 1688.110 ;
        RECT 1993.280 24.490 1993.540 24.810 ;
        RECT 2220.980 24.490 2221.240 24.810 ;
        RECT 2221.040 2.400 2221.180 24.490 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1437.185 1635.485 1437.355 1671.695 ;
        RECT 1436.725 1558.985 1436.895 1587.035 ;
        RECT 1436.725 1449.165 1436.895 1497.275 ;
        RECT 1436.725 1352.605 1436.895 1400.715 ;
        RECT 1436.725 1256.045 1436.895 1304.155 ;
        RECT 1436.725 772.905 1436.895 821.015 ;
        RECT 1436.265 688.925 1436.435 717.655 ;
        RECT 1436.725 524.365 1436.895 572.475 ;
      LAYER mcon ;
        RECT 1437.185 1671.525 1437.355 1671.695 ;
        RECT 1436.725 1586.865 1436.895 1587.035 ;
        RECT 1436.725 1497.105 1436.895 1497.275 ;
        RECT 1436.725 1400.545 1436.895 1400.715 ;
        RECT 1436.725 1303.985 1436.895 1304.155 ;
        RECT 1436.725 820.845 1436.895 821.015 ;
        RECT 1436.265 717.485 1436.435 717.655 ;
        RECT 1436.725 572.305 1436.895 572.475 ;
      LAYER met1 ;
        RECT 1437.125 1671.680 1437.415 1671.725 ;
        RECT 1439.870 1671.680 1440.190 1671.740 ;
        RECT 1437.125 1671.540 1440.190 1671.680 ;
        RECT 1437.125 1671.495 1437.415 1671.540 ;
        RECT 1439.870 1671.480 1440.190 1671.540 ;
        RECT 1437.110 1635.640 1437.430 1635.700 ;
        RECT 1436.915 1635.500 1437.430 1635.640 ;
        RECT 1437.110 1635.440 1437.430 1635.500 ;
        RECT 1436.650 1587.020 1436.970 1587.080 ;
        RECT 1436.455 1586.880 1436.970 1587.020 ;
        RECT 1436.650 1586.820 1436.970 1586.880 ;
        RECT 1436.650 1559.140 1436.970 1559.200 ;
        RECT 1436.455 1559.000 1436.970 1559.140 ;
        RECT 1436.650 1558.940 1436.970 1559.000 ;
        RECT 1436.650 1497.260 1436.970 1497.320 ;
        RECT 1436.455 1497.120 1436.970 1497.260 ;
        RECT 1436.650 1497.060 1436.970 1497.120 ;
        RECT 1436.650 1449.320 1436.970 1449.380 ;
        RECT 1436.455 1449.180 1436.970 1449.320 ;
        RECT 1436.650 1449.120 1436.970 1449.180 ;
        RECT 1436.650 1400.700 1436.970 1400.760 ;
        RECT 1436.455 1400.560 1436.970 1400.700 ;
        RECT 1436.650 1400.500 1436.970 1400.560 ;
        RECT 1436.650 1352.760 1436.970 1352.820 ;
        RECT 1436.455 1352.620 1436.970 1352.760 ;
        RECT 1436.650 1352.560 1436.970 1352.620 ;
        RECT 1436.650 1304.140 1436.970 1304.200 ;
        RECT 1436.455 1304.000 1436.970 1304.140 ;
        RECT 1436.650 1303.940 1436.970 1304.000 ;
        RECT 1436.650 1256.200 1436.970 1256.260 ;
        RECT 1436.455 1256.060 1436.970 1256.200 ;
        RECT 1436.650 1256.000 1436.970 1256.060 ;
        RECT 1436.650 1172.700 1436.970 1172.960 ;
        RECT 1436.740 1172.280 1436.880 1172.700 ;
        RECT 1436.650 1172.020 1436.970 1172.280 ;
        RECT 1436.650 1062.740 1436.970 1062.800 ;
        RECT 1437.570 1062.740 1437.890 1062.800 ;
        RECT 1436.650 1062.600 1437.890 1062.740 ;
        RECT 1436.650 1062.540 1436.970 1062.600 ;
        RECT 1437.570 1062.540 1437.890 1062.600 ;
        RECT 1436.650 966.180 1436.970 966.240 ;
        RECT 1437.570 966.180 1437.890 966.240 ;
        RECT 1436.650 966.040 1437.890 966.180 ;
        RECT 1436.650 965.980 1436.970 966.040 ;
        RECT 1437.570 965.980 1437.890 966.040 ;
        RECT 1436.190 883.560 1436.510 883.620 ;
        RECT 1436.190 883.420 1436.880 883.560 ;
        RECT 1436.190 883.360 1436.510 883.420 ;
        RECT 1436.740 883.280 1436.880 883.420 ;
        RECT 1436.650 883.020 1436.970 883.280 ;
        RECT 1436.650 821.000 1436.970 821.060 ;
        RECT 1436.455 820.860 1436.970 821.000 ;
        RECT 1436.650 820.800 1436.970 820.860 ;
        RECT 1436.650 773.060 1436.970 773.120 ;
        RECT 1436.455 772.920 1436.970 773.060 ;
        RECT 1436.650 772.860 1436.970 772.920 ;
        RECT 1436.190 725.120 1436.510 725.180 ;
        RECT 1436.650 725.120 1436.970 725.180 ;
        RECT 1436.190 724.980 1436.970 725.120 ;
        RECT 1436.190 724.920 1436.510 724.980 ;
        RECT 1436.650 724.920 1436.970 724.980 ;
        RECT 1436.190 717.640 1436.510 717.700 ;
        RECT 1435.995 717.500 1436.510 717.640 ;
        RECT 1436.190 717.440 1436.510 717.500 ;
        RECT 1436.205 689.080 1436.495 689.125 ;
        RECT 1437.110 689.080 1437.430 689.140 ;
        RECT 1436.205 688.940 1437.430 689.080 ;
        RECT 1436.205 688.895 1436.495 688.940 ;
        RECT 1437.110 688.880 1437.430 688.940 ;
        RECT 1436.650 669.360 1436.970 669.420 ;
        RECT 1437.570 669.360 1437.890 669.420 ;
        RECT 1436.650 669.220 1437.890 669.360 ;
        RECT 1436.650 669.160 1436.970 669.220 ;
        RECT 1437.570 669.160 1437.890 669.220 ;
        RECT 1436.190 620.540 1436.510 620.800 ;
        RECT 1436.280 620.400 1436.420 620.540 ;
        RECT 1437.110 620.400 1437.430 620.460 ;
        RECT 1436.280 620.260 1437.430 620.400 ;
        RECT 1437.110 620.200 1437.430 620.260 ;
        RECT 1436.650 572.460 1436.970 572.520 ;
        RECT 1436.455 572.320 1436.970 572.460 ;
        RECT 1436.650 572.260 1436.970 572.320 ;
        RECT 1436.650 524.520 1436.970 524.580 ;
        RECT 1436.455 524.380 1436.970 524.520 ;
        RECT 1436.650 524.320 1436.970 524.380 ;
        RECT 1436.650 427.960 1436.970 428.020 ;
        RECT 1437.110 427.960 1437.430 428.020 ;
        RECT 1436.650 427.820 1437.430 427.960 ;
        RECT 1436.650 427.760 1436.970 427.820 ;
        RECT 1437.110 427.760 1437.430 427.820 ;
        RECT 1436.650 400.560 1436.970 400.820 ;
        RECT 1436.740 400.140 1436.880 400.560 ;
        RECT 1436.650 399.880 1436.970 400.140 ;
        RECT 1436.650 352.280 1436.970 352.540 ;
        RECT 1436.740 351.860 1436.880 352.280 ;
        RECT 1436.650 351.600 1436.970 351.860 ;
        RECT 1436.650 289.920 1436.970 289.980 ;
        RECT 1437.110 289.920 1437.430 289.980 ;
        RECT 1436.650 289.780 1437.430 289.920 ;
        RECT 1436.650 289.720 1436.970 289.780 ;
        RECT 1437.110 289.720 1437.430 289.780 ;
        RECT 1436.650 256.260 1436.970 256.320 ;
        RECT 1436.280 256.120 1436.970 256.260 ;
        RECT 1436.280 255.300 1436.420 256.120 ;
        RECT 1436.650 256.060 1436.970 256.120 ;
        RECT 1436.190 255.040 1436.510 255.300 ;
        RECT 1436.190 193.500 1436.510 193.760 ;
        RECT 1436.280 193.080 1436.420 193.500 ;
        RECT 1436.190 192.820 1436.510 193.080 ;
        RECT 779.310 66.540 779.630 66.600 ;
        RECT 1436.650 66.540 1436.970 66.600 ;
        RECT 779.310 66.400 1436.970 66.540 ;
        RECT 779.310 66.340 779.630 66.400 ;
        RECT 1436.650 66.340 1436.970 66.400 ;
        RECT 775.630 2.960 775.950 3.020 ;
        RECT 779.310 2.960 779.630 3.020 ;
        RECT 775.630 2.820 779.630 2.960 ;
        RECT 775.630 2.760 775.950 2.820 ;
        RECT 779.310 2.760 779.630 2.820 ;
      LAYER via ;
        RECT 1439.900 1671.480 1440.160 1671.740 ;
        RECT 1437.140 1635.440 1437.400 1635.700 ;
        RECT 1436.680 1586.820 1436.940 1587.080 ;
        RECT 1436.680 1558.940 1436.940 1559.200 ;
        RECT 1436.680 1497.060 1436.940 1497.320 ;
        RECT 1436.680 1449.120 1436.940 1449.380 ;
        RECT 1436.680 1400.500 1436.940 1400.760 ;
        RECT 1436.680 1352.560 1436.940 1352.820 ;
        RECT 1436.680 1303.940 1436.940 1304.200 ;
        RECT 1436.680 1256.000 1436.940 1256.260 ;
        RECT 1436.680 1172.700 1436.940 1172.960 ;
        RECT 1436.680 1172.020 1436.940 1172.280 ;
        RECT 1436.680 1062.540 1436.940 1062.800 ;
        RECT 1437.600 1062.540 1437.860 1062.800 ;
        RECT 1436.680 965.980 1436.940 966.240 ;
        RECT 1437.600 965.980 1437.860 966.240 ;
        RECT 1436.220 883.360 1436.480 883.620 ;
        RECT 1436.680 883.020 1436.940 883.280 ;
        RECT 1436.680 820.800 1436.940 821.060 ;
        RECT 1436.680 772.860 1436.940 773.120 ;
        RECT 1436.220 724.920 1436.480 725.180 ;
        RECT 1436.680 724.920 1436.940 725.180 ;
        RECT 1436.220 717.440 1436.480 717.700 ;
        RECT 1437.140 688.880 1437.400 689.140 ;
        RECT 1436.680 669.160 1436.940 669.420 ;
        RECT 1437.600 669.160 1437.860 669.420 ;
        RECT 1436.220 620.540 1436.480 620.800 ;
        RECT 1437.140 620.200 1437.400 620.460 ;
        RECT 1436.680 572.260 1436.940 572.520 ;
        RECT 1436.680 524.320 1436.940 524.580 ;
        RECT 1436.680 427.760 1436.940 428.020 ;
        RECT 1437.140 427.760 1437.400 428.020 ;
        RECT 1436.680 400.560 1436.940 400.820 ;
        RECT 1436.680 399.880 1436.940 400.140 ;
        RECT 1436.680 352.280 1436.940 352.540 ;
        RECT 1436.680 351.600 1436.940 351.860 ;
        RECT 1436.680 289.720 1436.940 289.980 ;
        RECT 1437.140 289.720 1437.400 289.980 ;
        RECT 1436.680 256.060 1436.940 256.320 ;
        RECT 1436.220 255.040 1436.480 255.300 ;
        RECT 1436.220 193.500 1436.480 193.760 ;
        RECT 1436.220 192.820 1436.480 193.080 ;
        RECT 779.340 66.340 779.600 66.600 ;
        RECT 1436.680 66.340 1436.940 66.600 ;
        RECT 775.660 2.760 775.920 3.020 ;
        RECT 779.340 2.760 779.600 3.020 ;
      LAYER met2 ;
        RECT 1441.665 1700.410 1441.945 1704.000 ;
        RECT 1439.960 1700.270 1441.945 1700.410 ;
        RECT 1439.960 1671.770 1440.100 1700.270 ;
        RECT 1441.665 1700.000 1441.945 1700.270 ;
        RECT 1439.900 1671.450 1440.160 1671.770 ;
        RECT 1437.140 1635.410 1437.400 1635.730 ;
        RECT 1437.200 1594.330 1437.340 1635.410 ;
        RECT 1436.740 1594.190 1437.340 1594.330 ;
        RECT 1436.740 1587.110 1436.880 1594.190 ;
        RECT 1436.680 1586.790 1436.940 1587.110 ;
        RECT 1436.680 1558.910 1436.940 1559.230 ;
        RECT 1436.740 1497.350 1436.880 1558.910 ;
        RECT 1436.680 1497.030 1436.940 1497.350 ;
        RECT 1436.680 1449.090 1436.940 1449.410 ;
        RECT 1436.740 1400.790 1436.880 1449.090 ;
        RECT 1436.680 1400.470 1436.940 1400.790 ;
        RECT 1436.680 1352.530 1436.940 1352.850 ;
        RECT 1436.740 1304.230 1436.880 1352.530 ;
        RECT 1436.680 1303.910 1436.940 1304.230 ;
        RECT 1436.680 1255.970 1436.940 1256.290 ;
        RECT 1436.740 1172.990 1436.880 1255.970 ;
        RECT 1436.680 1172.670 1436.940 1172.990 ;
        RECT 1436.680 1171.990 1436.940 1172.310 ;
        RECT 1436.740 1110.965 1436.880 1171.990 ;
        RECT 1436.670 1110.595 1436.950 1110.965 ;
        RECT 1437.590 1110.595 1437.870 1110.965 ;
        RECT 1437.660 1062.830 1437.800 1110.595 ;
        RECT 1436.680 1062.510 1436.940 1062.830 ;
        RECT 1437.600 1062.510 1437.860 1062.830 ;
        RECT 1436.740 1014.405 1436.880 1062.510 ;
        RECT 1436.670 1014.035 1436.950 1014.405 ;
        RECT 1437.590 1014.035 1437.870 1014.405 ;
        RECT 1437.660 966.270 1437.800 1014.035 ;
        RECT 1436.680 965.950 1436.940 966.270 ;
        RECT 1437.600 965.950 1437.860 966.270 ;
        RECT 1436.740 917.730 1436.880 965.950 ;
        RECT 1436.280 917.590 1436.880 917.730 ;
        RECT 1436.280 883.650 1436.420 917.590 ;
        RECT 1436.220 883.330 1436.480 883.650 ;
        RECT 1436.680 882.990 1436.940 883.310 ;
        RECT 1436.740 821.090 1436.880 882.990 ;
        RECT 1436.680 820.770 1436.940 821.090 ;
        RECT 1436.680 772.830 1436.940 773.150 ;
        RECT 1436.740 725.210 1436.880 772.830 ;
        RECT 1436.220 724.890 1436.480 725.210 ;
        RECT 1436.680 724.890 1436.940 725.210 ;
        RECT 1436.280 717.730 1436.420 724.890 ;
        RECT 1436.220 717.410 1436.480 717.730 ;
        RECT 1437.140 688.850 1437.400 689.170 ;
        RECT 1437.200 669.530 1437.340 688.850 ;
        RECT 1436.740 669.450 1437.340 669.530 ;
        RECT 1436.680 669.390 1437.340 669.450 ;
        RECT 1436.680 669.130 1436.940 669.390 ;
        RECT 1437.600 669.130 1437.860 669.450 ;
        RECT 1436.740 668.975 1436.880 669.130 ;
        RECT 1437.660 621.365 1437.800 669.130 ;
        RECT 1436.210 620.995 1436.490 621.365 ;
        RECT 1437.590 620.995 1437.870 621.365 ;
        RECT 1436.280 620.830 1436.420 620.995 ;
        RECT 1436.220 620.510 1436.480 620.830 ;
        RECT 1437.140 620.170 1437.400 620.490 ;
        RECT 1437.200 579.090 1437.340 620.170 ;
        RECT 1436.740 578.950 1437.340 579.090 ;
        RECT 1436.740 572.550 1436.880 578.950 ;
        RECT 1436.680 572.230 1436.940 572.550 ;
        RECT 1436.680 524.290 1436.940 524.610 ;
        RECT 1436.740 497.490 1436.880 524.290 ;
        RECT 1436.740 497.350 1437.340 497.490 ;
        RECT 1437.200 428.050 1437.340 497.350 ;
        RECT 1436.680 427.730 1436.940 428.050 ;
        RECT 1437.140 427.730 1437.400 428.050 ;
        RECT 1436.740 400.850 1436.880 427.730 ;
        RECT 1436.680 400.530 1436.940 400.850 ;
        RECT 1436.680 399.850 1436.940 400.170 ;
        RECT 1436.740 352.570 1436.880 399.850 ;
        RECT 1436.680 352.250 1436.940 352.570 ;
        RECT 1436.680 351.570 1436.940 351.890 ;
        RECT 1436.740 338.485 1436.880 351.570 ;
        RECT 1436.670 338.115 1436.950 338.485 ;
        RECT 1437.130 337.435 1437.410 337.805 ;
        RECT 1437.200 290.010 1437.340 337.435 ;
        RECT 1436.680 289.690 1436.940 290.010 ;
        RECT 1437.140 289.690 1437.400 290.010 ;
        RECT 1436.740 256.350 1436.880 289.690 ;
        RECT 1436.680 256.030 1436.940 256.350 ;
        RECT 1436.220 255.010 1436.480 255.330 ;
        RECT 1436.280 193.790 1436.420 255.010 ;
        RECT 1436.220 193.470 1436.480 193.790 ;
        RECT 1436.220 192.790 1436.480 193.110 ;
        RECT 1436.280 144.685 1436.420 192.790 ;
        RECT 1436.210 144.315 1436.490 144.685 ;
        RECT 1436.670 143.635 1436.950 144.005 ;
        RECT 1436.740 66.630 1436.880 143.635 ;
        RECT 779.340 66.310 779.600 66.630 ;
        RECT 1436.680 66.310 1436.940 66.630 ;
        RECT 779.400 3.050 779.540 66.310 ;
        RECT 775.660 2.730 775.920 3.050 ;
        RECT 779.340 2.730 779.600 3.050 ;
        RECT 775.720 2.400 775.860 2.730 ;
        RECT 775.510 -4.800 776.070 2.400 ;
      LAYER via2 ;
        RECT 1436.670 1110.640 1436.950 1110.920 ;
        RECT 1437.590 1110.640 1437.870 1110.920 ;
        RECT 1436.670 1014.080 1436.950 1014.360 ;
        RECT 1437.590 1014.080 1437.870 1014.360 ;
        RECT 1436.210 621.040 1436.490 621.320 ;
        RECT 1437.590 621.040 1437.870 621.320 ;
        RECT 1436.670 338.160 1436.950 338.440 ;
        RECT 1437.130 337.480 1437.410 337.760 ;
        RECT 1436.210 144.360 1436.490 144.640 ;
        RECT 1436.670 143.680 1436.950 143.960 ;
      LAYER met3 ;
        RECT 1436.645 1110.930 1436.975 1110.945 ;
        RECT 1437.565 1110.930 1437.895 1110.945 ;
        RECT 1436.645 1110.630 1437.895 1110.930 ;
        RECT 1436.645 1110.615 1436.975 1110.630 ;
        RECT 1437.565 1110.615 1437.895 1110.630 ;
        RECT 1436.645 1014.370 1436.975 1014.385 ;
        RECT 1437.565 1014.370 1437.895 1014.385 ;
        RECT 1436.645 1014.070 1437.895 1014.370 ;
        RECT 1436.645 1014.055 1436.975 1014.070 ;
        RECT 1437.565 1014.055 1437.895 1014.070 ;
        RECT 1436.185 621.330 1436.515 621.345 ;
        RECT 1437.565 621.330 1437.895 621.345 ;
        RECT 1436.185 621.030 1437.895 621.330 ;
        RECT 1436.185 621.015 1436.515 621.030 ;
        RECT 1437.565 621.015 1437.895 621.030 ;
        RECT 1436.645 338.450 1436.975 338.465 ;
        RECT 1436.430 338.135 1436.975 338.450 ;
        RECT 1436.430 337.770 1436.730 338.135 ;
        RECT 1437.105 337.770 1437.435 337.785 ;
        RECT 1436.430 337.470 1437.435 337.770 ;
        RECT 1437.105 337.455 1437.435 337.470 ;
        RECT 1436.185 144.650 1436.515 144.665 ;
        RECT 1435.510 144.350 1436.515 144.650 ;
        RECT 1435.510 143.970 1435.810 144.350 ;
        RECT 1436.185 144.335 1436.515 144.350 ;
        RECT 1436.645 143.970 1436.975 143.985 ;
        RECT 1435.510 143.670 1436.975 143.970 ;
        RECT 1436.645 143.655 1436.975 143.670 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 24.040 1994.030 24.100 ;
        RECT 2238.890 24.040 2239.210 24.100 ;
        RECT 1993.710 23.900 2239.210 24.040 ;
        RECT 1993.710 23.840 1994.030 23.900 ;
        RECT 2238.890 23.840 2239.210 23.900 ;
      LAYER via ;
        RECT 1993.740 23.840 1994.000 24.100 ;
        RECT 2238.920 23.840 2239.180 24.100 ;
      LAYER met2 ;
        RECT 1993.665 1700.000 1993.945 1704.000 ;
        RECT 1993.800 24.130 1993.940 1700.000 ;
        RECT 1993.740 23.810 1994.000 24.130 ;
        RECT 2238.920 23.810 2239.180 24.130 ;
        RECT 2238.980 2.400 2239.120 23.810 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2000.610 20.980 2000.930 21.040 ;
        RECT 2256.370 20.980 2256.690 21.040 ;
        RECT 2000.610 20.840 2256.690 20.980 ;
        RECT 2000.610 20.780 2000.930 20.840 ;
        RECT 2256.370 20.780 2256.690 20.840 ;
      LAYER via ;
        RECT 2000.640 20.780 2000.900 21.040 ;
        RECT 2256.400 20.780 2256.660 21.040 ;
      LAYER met2 ;
        RECT 2000.565 1700.000 2000.845 1704.000 ;
        RECT 2000.700 21.070 2000.840 1700.000 ;
        RECT 2000.640 20.750 2000.900 21.070 ;
        RECT 2256.400 20.750 2256.660 21.070 ;
        RECT 2256.460 2.400 2256.600 20.750 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2007.510 28.120 2007.830 28.180 ;
        RECT 2274.310 28.120 2274.630 28.180 ;
        RECT 2007.510 27.980 2274.630 28.120 ;
        RECT 2007.510 27.920 2007.830 27.980 ;
        RECT 2274.310 27.920 2274.630 27.980 ;
      LAYER via ;
        RECT 2007.540 27.920 2007.800 28.180 ;
        RECT 2274.340 27.920 2274.600 28.180 ;
      LAYER met2 ;
        RECT 2007.465 1700.000 2007.745 1704.000 ;
        RECT 2007.600 28.210 2007.740 1700.000 ;
        RECT 2007.540 27.890 2007.800 28.210 ;
        RECT 2274.340 27.890 2274.600 28.210 ;
        RECT 2274.400 2.400 2274.540 27.890 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2014.410 28.460 2014.730 28.520 ;
        RECT 2292.250 28.460 2292.570 28.520 ;
        RECT 2014.410 28.320 2292.570 28.460 ;
        RECT 2014.410 28.260 2014.730 28.320 ;
        RECT 2292.250 28.260 2292.570 28.320 ;
      LAYER via ;
        RECT 2014.440 28.260 2014.700 28.520 ;
        RECT 2292.280 28.260 2292.540 28.520 ;
      LAYER met2 ;
        RECT 2013.905 1700.410 2014.185 1704.000 ;
        RECT 2013.905 1700.270 2014.640 1700.410 ;
        RECT 2013.905 1700.000 2014.185 1700.270 ;
        RECT 2014.500 28.550 2014.640 1700.270 ;
        RECT 2014.440 28.230 2014.700 28.550 ;
        RECT 2292.280 28.230 2292.540 28.550 ;
        RECT 2292.340 2.400 2292.480 28.230 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2021.310 28.800 2021.630 28.860 ;
        RECT 2310.190 28.800 2310.510 28.860 ;
        RECT 2021.310 28.660 2310.510 28.800 ;
        RECT 2021.310 28.600 2021.630 28.660 ;
        RECT 2310.190 28.600 2310.510 28.660 ;
      LAYER via ;
        RECT 2021.340 28.600 2021.600 28.860 ;
        RECT 2310.220 28.600 2310.480 28.860 ;
      LAYER met2 ;
        RECT 2020.805 1700.410 2021.085 1704.000 ;
        RECT 2020.805 1700.270 2021.540 1700.410 ;
        RECT 2020.805 1700.000 2021.085 1700.270 ;
        RECT 2021.400 28.890 2021.540 1700.270 ;
        RECT 2021.340 28.570 2021.600 28.890 ;
        RECT 2310.220 28.570 2310.480 28.890 ;
        RECT 2310.280 2.400 2310.420 28.570 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2028.210 29.140 2028.530 29.200 ;
        RECT 2328.130 29.140 2328.450 29.200 ;
        RECT 2028.210 29.000 2328.450 29.140 ;
        RECT 2028.210 28.940 2028.530 29.000 ;
        RECT 2328.130 28.940 2328.450 29.000 ;
      LAYER via ;
        RECT 2028.240 28.940 2028.500 29.200 ;
        RECT 2328.160 28.940 2328.420 29.200 ;
      LAYER met2 ;
        RECT 2027.245 1700.410 2027.525 1704.000 ;
        RECT 2027.245 1700.270 2028.440 1700.410 ;
        RECT 2027.245 1700.000 2027.525 1700.270 ;
        RECT 2028.300 29.230 2028.440 1700.270 ;
        RECT 2028.240 28.910 2028.500 29.230 ;
        RECT 2328.160 28.910 2328.420 29.230 ;
        RECT 2328.220 2.400 2328.360 28.910 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2035.110 29.480 2035.430 29.540 ;
        RECT 2345.610 29.480 2345.930 29.540 ;
        RECT 2035.110 29.340 2345.930 29.480 ;
        RECT 2035.110 29.280 2035.430 29.340 ;
        RECT 2345.610 29.280 2345.930 29.340 ;
      LAYER via ;
        RECT 2035.140 29.280 2035.400 29.540 ;
        RECT 2345.640 29.280 2345.900 29.540 ;
      LAYER met2 ;
        RECT 2034.145 1700.410 2034.425 1704.000 ;
        RECT 2034.145 1700.270 2035.340 1700.410 ;
        RECT 2034.145 1700.000 2034.425 1700.270 ;
        RECT 2035.200 29.570 2035.340 1700.270 ;
        RECT 2035.140 29.250 2035.400 29.570 ;
        RECT 2345.640 29.250 2345.900 29.570 ;
        RECT 2345.700 2.400 2345.840 29.250 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 29.820 2042.330 29.880 ;
        RECT 2363.550 29.820 2363.870 29.880 ;
        RECT 2042.010 29.680 2363.870 29.820 ;
        RECT 2042.010 29.620 2042.330 29.680 ;
        RECT 2363.550 29.620 2363.870 29.680 ;
      LAYER via ;
        RECT 2042.040 29.620 2042.300 29.880 ;
        RECT 2363.580 29.620 2363.840 29.880 ;
      LAYER met2 ;
        RECT 2041.045 1700.410 2041.325 1704.000 ;
        RECT 2041.045 1700.270 2042.240 1700.410 ;
        RECT 2041.045 1700.000 2041.325 1700.270 ;
        RECT 2042.100 29.910 2042.240 1700.270 ;
        RECT 2042.040 29.590 2042.300 29.910 ;
        RECT 2363.580 29.590 2363.840 29.910 ;
        RECT 2363.640 2.400 2363.780 29.590 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.910 30.160 2049.230 30.220 ;
        RECT 2381.490 30.160 2381.810 30.220 ;
        RECT 2048.910 30.020 2381.810 30.160 ;
        RECT 2048.910 29.960 2049.230 30.020 ;
        RECT 2381.490 29.960 2381.810 30.020 ;
      LAYER via ;
        RECT 2048.940 29.960 2049.200 30.220 ;
        RECT 2381.520 29.960 2381.780 30.220 ;
      LAYER met2 ;
        RECT 2047.485 1700.410 2047.765 1704.000 ;
        RECT 2047.485 1700.270 2049.140 1700.410 ;
        RECT 2047.485 1700.000 2047.765 1700.270 ;
        RECT 2049.000 30.250 2049.140 1700.270 ;
        RECT 2048.940 29.930 2049.200 30.250 ;
        RECT 2381.520 29.930 2381.780 30.250 ;
        RECT 2381.580 2.400 2381.720 29.930 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.810 30.500 2056.130 30.560 ;
        RECT 2399.430 30.500 2399.750 30.560 ;
        RECT 2055.810 30.360 2399.750 30.500 ;
        RECT 2055.810 30.300 2056.130 30.360 ;
        RECT 2399.430 30.300 2399.750 30.360 ;
      LAYER via ;
        RECT 2055.840 30.300 2056.100 30.560 ;
        RECT 2399.460 30.300 2399.720 30.560 ;
      LAYER met2 ;
        RECT 2054.385 1700.410 2054.665 1704.000 ;
        RECT 2054.385 1700.270 2056.040 1700.410 ;
        RECT 2054.385 1700.000 2054.665 1700.270 ;
        RECT 2055.900 30.590 2056.040 1700.270 ;
        RECT 2055.840 30.270 2056.100 30.590 ;
        RECT 2399.460 30.270 2399.720 30.590 ;
        RECT 2399.520 2.400 2399.660 30.270 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1443.625 1414.145 1443.795 1448.655 ;
        RECT 1443.625 1317.585 1443.795 1352.095 ;
        RECT 1443.625 1159.145 1443.795 1200.455 ;
        RECT 1443.625 1062.585 1443.795 1076.695 ;
        RECT 1444.085 1014.305 1444.255 1028.415 ;
        RECT 1443.625 966.025 1443.795 980.135 ;
        RECT 1444.085 917.745 1444.255 931.855 ;
        RECT 1443.625 769.165 1443.795 807.075 ;
        RECT 1444.085 697.425 1444.255 745.195 ;
        RECT 1443.625 524.365 1443.795 572.475 ;
        RECT 1443.165 430.525 1443.335 497.335 ;
        RECT 1443.625 289.765 1443.795 369.155 ;
      LAYER mcon ;
        RECT 1443.625 1448.485 1443.795 1448.655 ;
        RECT 1443.625 1351.925 1443.795 1352.095 ;
        RECT 1443.625 1200.285 1443.795 1200.455 ;
        RECT 1443.625 1076.525 1443.795 1076.695 ;
        RECT 1444.085 1028.245 1444.255 1028.415 ;
        RECT 1443.625 979.965 1443.795 980.135 ;
        RECT 1444.085 931.685 1444.255 931.855 ;
        RECT 1443.625 806.905 1443.795 807.075 ;
        RECT 1444.085 745.025 1444.255 745.195 ;
        RECT 1443.625 572.305 1443.795 572.475 ;
        RECT 1443.165 497.165 1443.335 497.335 ;
        RECT 1443.625 368.985 1443.795 369.155 ;
      LAYER met1 ;
        RECT 1444.010 1642.440 1444.330 1642.500 ;
        RECT 1447.690 1642.440 1448.010 1642.500 ;
        RECT 1444.010 1642.300 1448.010 1642.440 ;
        RECT 1444.010 1642.240 1444.330 1642.300 ;
        RECT 1447.690 1642.240 1448.010 1642.300 ;
        RECT 1443.550 1511.340 1443.870 1511.600 ;
        RECT 1443.640 1510.920 1443.780 1511.340 ;
        RECT 1443.550 1510.660 1443.870 1510.920 ;
        RECT 1443.550 1449.320 1443.870 1449.380 ;
        RECT 1444.930 1449.320 1445.250 1449.380 ;
        RECT 1443.550 1449.180 1445.250 1449.320 ;
        RECT 1443.550 1449.120 1443.870 1449.180 ;
        RECT 1444.930 1449.120 1445.250 1449.180 ;
        RECT 1443.550 1448.640 1443.870 1448.700 ;
        RECT 1443.355 1448.500 1443.870 1448.640 ;
        RECT 1443.550 1448.440 1443.870 1448.500 ;
        RECT 1443.550 1414.300 1443.870 1414.360 ;
        RECT 1443.355 1414.160 1443.870 1414.300 ;
        RECT 1443.550 1414.100 1443.870 1414.160 ;
        RECT 1443.090 1352.760 1443.410 1352.820 ;
        RECT 1443.550 1352.760 1443.870 1352.820 ;
        RECT 1443.090 1352.620 1443.870 1352.760 ;
        RECT 1443.090 1352.560 1443.410 1352.620 ;
        RECT 1443.550 1352.560 1443.870 1352.620 ;
        RECT 1443.550 1352.080 1443.870 1352.140 ;
        RECT 1443.355 1351.940 1443.870 1352.080 ;
        RECT 1443.550 1351.880 1443.870 1351.940 ;
        RECT 1443.550 1317.740 1443.870 1317.800 ;
        RECT 1443.355 1317.600 1443.870 1317.740 ;
        RECT 1443.550 1317.540 1443.870 1317.600 ;
        RECT 1443.090 1256.200 1443.410 1256.260 ;
        RECT 1443.550 1256.200 1443.870 1256.260 ;
        RECT 1443.090 1256.060 1443.870 1256.200 ;
        RECT 1443.090 1256.000 1443.410 1256.060 ;
        RECT 1443.550 1256.000 1443.870 1256.060 ;
        RECT 1443.550 1221.320 1443.870 1221.580 ;
        RECT 1443.640 1220.840 1443.780 1221.320 ;
        RECT 1444.010 1220.840 1444.330 1220.900 ;
        RECT 1443.640 1220.700 1444.330 1220.840 ;
        RECT 1444.010 1220.640 1444.330 1220.700 ;
        RECT 1443.550 1200.440 1443.870 1200.500 ;
        RECT 1443.355 1200.300 1443.870 1200.440 ;
        RECT 1443.550 1200.240 1443.870 1200.300 ;
        RECT 1443.565 1159.300 1443.855 1159.345 ;
        RECT 1444.010 1159.300 1444.330 1159.360 ;
        RECT 1443.565 1159.160 1444.330 1159.300 ;
        RECT 1443.565 1159.115 1443.855 1159.160 ;
        RECT 1444.010 1159.100 1444.330 1159.160 ;
        RECT 1444.010 1124.760 1444.330 1125.020 ;
        RECT 1444.100 1124.340 1444.240 1124.760 ;
        RECT 1444.010 1124.080 1444.330 1124.340 ;
        RECT 1443.550 1076.680 1443.870 1076.740 ;
        RECT 1443.355 1076.540 1443.870 1076.680 ;
        RECT 1443.550 1076.480 1443.870 1076.540 ;
        RECT 1443.565 1062.740 1443.855 1062.785 ;
        RECT 1444.010 1062.740 1444.330 1062.800 ;
        RECT 1443.565 1062.600 1444.330 1062.740 ;
        RECT 1443.565 1062.555 1443.855 1062.600 ;
        RECT 1444.010 1062.540 1444.330 1062.600 ;
        RECT 1444.010 1028.400 1444.330 1028.460 ;
        RECT 1443.815 1028.260 1444.330 1028.400 ;
        RECT 1444.010 1028.200 1444.330 1028.260 ;
        RECT 1444.010 1014.460 1444.330 1014.520 ;
        RECT 1443.815 1014.320 1444.330 1014.460 ;
        RECT 1444.010 1014.260 1444.330 1014.320 ;
        RECT 1443.550 980.120 1443.870 980.180 ;
        RECT 1443.355 979.980 1443.870 980.120 ;
        RECT 1443.550 979.920 1443.870 979.980 ;
        RECT 1443.565 966.180 1443.855 966.225 ;
        RECT 1444.010 966.180 1444.330 966.240 ;
        RECT 1443.565 966.040 1444.330 966.180 ;
        RECT 1443.565 965.995 1443.855 966.040 ;
        RECT 1444.010 965.980 1444.330 966.040 ;
        RECT 1444.010 931.840 1444.330 931.900 ;
        RECT 1443.815 931.700 1444.330 931.840 ;
        RECT 1444.010 931.640 1444.330 931.700 ;
        RECT 1444.010 917.900 1444.330 917.960 ;
        RECT 1443.815 917.760 1444.330 917.900 ;
        RECT 1444.010 917.700 1444.330 917.760 ;
        RECT 1444.010 883.700 1444.330 883.960 ;
        RECT 1444.100 883.280 1444.240 883.700 ;
        RECT 1444.010 883.020 1444.330 883.280 ;
        RECT 1443.550 814.200 1443.870 814.260 ;
        RECT 1444.010 814.200 1444.330 814.260 ;
        RECT 1443.550 814.060 1444.330 814.200 ;
        RECT 1443.550 814.000 1443.870 814.060 ;
        RECT 1444.010 814.000 1444.330 814.060 ;
        RECT 1443.550 807.060 1443.870 807.120 ;
        RECT 1443.355 806.920 1443.870 807.060 ;
        RECT 1443.550 806.860 1443.870 806.920 ;
        RECT 1443.565 769.320 1443.855 769.365 ;
        RECT 1444.010 769.320 1444.330 769.380 ;
        RECT 1443.565 769.180 1444.330 769.320 ;
        RECT 1443.565 769.135 1443.855 769.180 ;
        RECT 1444.010 769.120 1444.330 769.180 ;
        RECT 1444.010 745.180 1444.330 745.240 ;
        RECT 1443.815 745.040 1444.330 745.180 ;
        RECT 1444.010 744.980 1444.330 745.040 ;
        RECT 1444.010 697.580 1444.330 697.640 ;
        RECT 1443.815 697.440 1444.330 697.580 ;
        RECT 1444.010 697.380 1444.330 697.440 ;
        RECT 1444.010 696.900 1444.330 696.960 ;
        RECT 1444.470 696.900 1444.790 696.960 ;
        RECT 1444.010 696.760 1444.790 696.900 ;
        RECT 1444.010 696.700 1444.330 696.760 ;
        RECT 1444.470 696.700 1444.790 696.760 ;
        RECT 1443.550 572.460 1443.870 572.520 ;
        RECT 1443.355 572.320 1443.870 572.460 ;
        RECT 1443.550 572.260 1443.870 572.320 ;
        RECT 1443.565 524.520 1443.855 524.565 ;
        RECT 1444.010 524.520 1444.330 524.580 ;
        RECT 1443.565 524.380 1444.330 524.520 ;
        RECT 1443.565 524.335 1443.855 524.380 ;
        RECT 1444.010 524.320 1444.330 524.380 ;
        RECT 1443.105 497.320 1443.395 497.365 ;
        RECT 1444.010 497.320 1444.330 497.380 ;
        RECT 1443.105 497.180 1444.330 497.320 ;
        RECT 1443.105 497.135 1443.395 497.180 ;
        RECT 1444.010 497.120 1444.330 497.180 ;
        RECT 1443.090 430.680 1443.410 430.740 ;
        RECT 1442.895 430.540 1443.410 430.680 ;
        RECT 1443.090 430.480 1443.410 430.540 ;
        RECT 1443.090 369.140 1443.410 369.200 ;
        RECT 1443.565 369.140 1443.855 369.185 ;
        RECT 1443.090 369.000 1443.855 369.140 ;
        RECT 1443.090 368.940 1443.410 369.000 ;
        RECT 1443.565 368.955 1443.855 369.000 ;
        RECT 1443.550 289.920 1443.870 289.980 ;
        RECT 1443.355 289.780 1443.870 289.920 ;
        RECT 1443.550 289.720 1443.870 289.780 ;
        RECT 1443.090 241.300 1443.410 241.360 ;
        RECT 1444.010 241.300 1444.330 241.360 ;
        RECT 1443.090 241.160 1444.330 241.300 ;
        RECT 1443.090 241.100 1443.410 241.160 ;
        RECT 1444.010 241.100 1444.330 241.160 ;
        RECT 1443.550 96.800 1443.870 96.860 ;
        RECT 1444.930 96.800 1445.250 96.860 ;
        RECT 1443.550 96.660 1445.250 96.800 ;
        RECT 1443.550 96.600 1443.870 96.660 ;
        RECT 1444.930 96.600 1445.250 96.660 ;
        RECT 800.010 66.880 800.330 66.940 ;
        RECT 1443.550 66.880 1443.870 66.940 ;
        RECT 800.010 66.740 1443.870 66.880 ;
        RECT 800.010 66.680 800.330 66.740 ;
        RECT 1443.550 66.680 1443.870 66.740 ;
        RECT 793.570 35.600 793.890 35.660 ;
        RECT 800.010 35.600 800.330 35.660 ;
        RECT 793.570 35.460 800.330 35.600 ;
        RECT 793.570 35.400 793.890 35.460 ;
        RECT 800.010 35.400 800.330 35.460 ;
      LAYER via ;
        RECT 1444.040 1642.240 1444.300 1642.500 ;
        RECT 1447.720 1642.240 1447.980 1642.500 ;
        RECT 1443.580 1511.340 1443.840 1511.600 ;
        RECT 1443.580 1510.660 1443.840 1510.920 ;
        RECT 1443.580 1449.120 1443.840 1449.380 ;
        RECT 1444.960 1449.120 1445.220 1449.380 ;
        RECT 1443.580 1448.440 1443.840 1448.700 ;
        RECT 1443.580 1414.100 1443.840 1414.360 ;
        RECT 1443.120 1352.560 1443.380 1352.820 ;
        RECT 1443.580 1352.560 1443.840 1352.820 ;
        RECT 1443.580 1351.880 1443.840 1352.140 ;
        RECT 1443.580 1317.540 1443.840 1317.800 ;
        RECT 1443.120 1256.000 1443.380 1256.260 ;
        RECT 1443.580 1256.000 1443.840 1256.260 ;
        RECT 1443.580 1221.320 1443.840 1221.580 ;
        RECT 1444.040 1220.640 1444.300 1220.900 ;
        RECT 1443.580 1200.240 1443.840 1200.500 ;
        RECT 1444.040 1159.100 1444.300 1159.360 ;
        RECT 1444.040 1124.760 1444.300 1125.020 ;
        RECT 1444.040 1124.080 1444.300 1124.340 ;
        RECT 1443.580 1076.480 1443.840 1076.740 ;
        RECT 1444.040 1062.540 1444.300 1062.800 ;
        RECT 1444.040 1028.200 1444.300 1028.460 ;
        RECT 1444.040 1014.260 1444.300 1014.520 ;
        RECT 1443.580 979.920 1443.840 980.180 ;
        RECT 1444.040 965.980 1444.300 966.240 ;
        RECT 1444.040 931.640 1444.300 931.900 ;
        RECT 1444.040 917.700 1444.300 917.960 ;
        RECT 1444.040 883.700 1444.300 883.960 ;
        RECT 1444.040 883.020 1444.300 883.280 ;
        RECT 1443.580 814.000 1443.840 814.260 ;
        RECT 1444.040 814.000 1444.300 814.260 ;
        RECT 1443.580 806.860 1443.840 807.120 ;
        RECT 1444.040 769.120 1444.300 769.380 ;
        RECT 1444.040 744.980 1444.300 745.240 ;
        RECT 1444.040 697.380 1444.300 697.640 ;
        RECT 1444.040 696.700 1444.300 696.960 ;
        RECT 1444.500 696.700 1444.760 696.960 ;
        RECT 1443.580 572.260 1443.840 572.520 ;
        RECT 1444.040 524.320 1444.300 524.580 ;
        RECT 1444.040 497.120 1444.300 497.380 ;
        RECT 1443.120 430.480 1443.380 430.740 ;
        RECT 1443.120 368.940 1443.380 369.200 ;
        RECT 1443.580 289.720 1443.840 289.980 ;
        RECT 1443.120 241.100 1443.380 241.360 ;
        RECT 1444.040 241.100 1444.300 241.360 ;
        RECT 1443.580 96.600 1443.840 96.860 ;
        RECT 1444.960 96.600 1445.220 96.860 ;
        RECT 800.040 66.680 800.300 66.940 ;
        RECT 1443.580 66.680 1443.840 66.940 ;
        RECT 793.600 35.400 793.860 35.660 ;
        RECT 800.040 35.400 800.300 35.660 ;
      LAYER met2 ;
        RECT 1448.105 1700.410 1448.385 1704.000 ;
        RECT 1447.780 1700.270 1448.385 1700.410 ;
        RECT 1447.780 1642.530 1447.920 1700.270 ;
        RECT 1448.105 1700.000 1448.385 1700.270 ;
        RECT 1444.040 1642.210 1444.300 1642.530 ;
        RECT 1447.720 1642.210 1447.980 1642.530 ;
        RECT 1444.100 1559.650 1444.240 1642.210 ;
        RECT 1443.640 1559.510 1444.240 1559.650 ;
        RECT 1443.640 1511.630 1443.780 1559.510 ;
        RECT 1443.580 1511.310 1443.840 1511.630 ;
        RECT 1443.580 1510.630 1443.840 1510.950 ;
        RECT 1443.640 1497.600 1443.780 1510.630 ;
        RECT 1443.640 1497.460 1444.240 1497.600 ;
        RECT 1444.100 1497.205 1444.240 1497.460 ;
        RECT 1444.030 1496.835 1444.310 1497.205 ;
        RECT 1444.950 1496.835 1445.230 1497.205 ;
        RECT 1445.020 1449.410 1445.160 1496.835 ;
        RECT 1443.580 1449.090 1443.840 1449.410 ;
        RECT 1444.960 1449.090 1445.220 1449.410 ;
        RECT 1443.640 1448.730 1443.780 1449.090 ;
        RECT 1443.580 1448.410 1443.840 1448.730 ;
        RECT 1443.580 1414.070 1443.840 1414.390 ;
        RECT 1443.640 1401.210 1443.780 1414.070 ;
        RECT 1443.640 1401.070 1444.240 1401.210 ;
        RECT 1444.100 1400.700 1444.240 1401.070 ;
        RECT 1443.640 1400.560 1444.240 1400.700 ;
        RECT 1443.640 1366.530 1443.780 1400.560 ;
        RECT 1443.180 1366.390 1443.780 1366.530 ;
        RECT 1443.180 1352.850 1443.320 1366.390 ;
        RECT 1443.120 1352.530 1443.380 1352.850 ;
        RECT 1443.580 1352.530 1443.840 1352.850 ;
        RECT 1443.640 1352.170 1443.780 1352.530 ;
        RECT 1443.580 1351.850 1443.840 1352.170 ;
        RECT 1443.580 1317.510 1443.840 1317.830 ;
        RECT 1443.640 1304.650 1443.780 1317.510 ;
        RECT 1443.640 1304.510 1444.240 1304.650 ;
        RECT 1444.100 1304.140 1444.240 1304.510 ;
        RECT 1443.640 1304.000 1444.240 1304.140 ;
        RECT 1443.640 1269.970 1443.780 1304.000 ;
        RECT 1443.180 1269.830 1443.780 1269.970 ;
        RECT 1443.180 1256.290 1443.320 1269.830 ;
        RECT 1443.120 1255.970 1443.380 1256.290 ;
        RECT 1443.580 1255.970 1443.840 1256.290 ;
        RECT 1443.640 1221.610 1443.780 1255.970 ;
        RECT 1443.580 1221.290 1443.840 1221.610 ;
        RECT 1444.040 1220.610 1444.300 1220.930 ;
        RECT 1444.100 1207.410 1444.240 1220.610 ;
        RECT 1443.640 1207.270 1444.240 1207.410 ;
        RECT 1443.640 1200.530 1443.780 1207.270 ;
        RECT 1443.580 1200.210 1443.840 1200.530 ;
        RECT 1444.040 1159.070 1444.300 1159.390 ;
        RECT 1444.100 1125.050 1444.240 1159.070 ;
        RECT 1444.040 1124.730 1444.300 1125.050 ;
        RECT 1444.040 1124.050 1444.300 1124.370 ;
        RECT 1444.100 1110.850 1444.240 1124.050 ;
        RECT 1443.640 1110.710 1444.240 1110.850 ;
        RECT 1443.640 1076.770 1443.780 1110.710 ;
        RECT 1443.580 1076.450 1443.840 1076.770 ;
        RECT 1444.040 1062.510 1444.300 1062.830 ;
        RECT 1444.100 1028.490 1444.240 1062.510 ;
        RECT 1444.040 1028.170 1444.300 1028.490 ;
        RECT 1444.100 1014.550 1444.240 1014.705 ;
        RECT 1444.040 1014.290 1444.300 1014.550 ;
        RECT 1443.640 1014.230 1444.300 1014.290 ;
        RECT 1443.640 1014.150 1444.240 1014.230 ;
        RECT 1443.640 980.210 1443.780 1014.150 ;
        RECT 1443.580 979.890 1443.840 980.210 ;
        RECT 1444.040 965.950 1444.300 966.270 ;
        RECT 1444.100 931.930 1444.240 965.950 ;
        RECT 1444.040 931.610 1444.300 931.930 ;
        RECT 1444.040 917.670 1444.300 917.990 ;
        RECT 1444.100 883.990 1444.240 917.670 ;
        RECT 1444.040 883.670 1444.300 883.990 ;
        RECT 1444.040 882.990 1444.300 883.310 ;
        RECT 1444.100 814.290 1444.240 882.990 ;
        RECT 1443.580 813.970 1443.840 814.290 ;
        RECT 1444.040 813.970 1444.300 814.290 ;
        RECT 1443.640 807.150 1443.780 813.970 ;
        RECT 1443.580 806.830 1443.840 807.150 ;
        RECT 1444.040 769.090 1444.300 769.410 ;
        RECT 1444.100 745.270 1444.240 769.090 ;
        RECT 1444.040 744.950 1444.300 745.270 ;
        RECT 1444.040 697.350 1444.300 697.670 ;
        RECT 1444.100 696.990 1444.240 697.350 ;
        RECT 1444.040 696.670 1444.300 696.990 ;
        RECT 1444.500 696.670 1444.760 696.990 ;
        RECT 1444.560 640.970 1444.700 696.670 ;
        RECT 1444.100 640.830 1444.700 640.970 ;
        RECT 1444.100 572.970 1444.240 640.830 ;
        RECT 1443.640 572.830 1444.240 572.970 ;
        RECT 1443.640 572.550 1443.780 572.830 ;
        RECT 1443.580 572.230 1443.840 572.550 ;
        RECT 1444.040 524.290 1444.300 524.610 ;
        RECT 1444.100 497.410 1444.240 524.290 ;
        RECT 1444.040 497.090 1444.300 497.410 ;
        RECT 1443.120 430.450 1443.380 430.770 ;
        RECT 1443.180 369.230 1443.320 430.450 ;
        RECT 1443.120 368.910 1443.380 369.230 ;
        RECT 1443.580 289.690 1443.840 290.010 ;
        RECT 1443.640 265.610 1443.780 289.690 ;
        RECT 1443.640 265.470 1444.700 265.610 ;
        RECT 1444.560 254.730 1444.700 265.470 ;
        RECT 1444.100 254.590 1444.700 254.730 ;
        RECT 1444.100 241.390 1444.240 254.590 ;
        RECT 1443.120 241.070 1443.380 241.390 ;
        RECT 1444.040 241.070 1444.300 241.390 ;
        RECT 1443.180 193.530 1443.320 241.070 ;
        RECT 1443.180 193.390 1443.780 193.530 ;
        RECT 1443.640 169.050 1443.780 193.390 ;
        RECT 1443.640 168.910 1445.160 169.050 ;
        RECT 1445.020 96.890 1445.160 168.910 ;
        RECT 1443.580 96.570 1443.840 96.890 ;
        RECT 1444.960 96.570 1445.220 96.890 ;
        RECT 1443.640 66.970 1443.780 96.570 ;
        RECT 800.040 66.650 800.300 66.970 ;
        RECT 1443.580 66.650 1443.840 66.970 ;
        RECT 800.100 35.690 800.240 66.650 ;
        RECT 793.600 35.370 793.860 35.690 ;
        RECT 800.040 35.370 800.300 35.690 ;
        RECT 793.660 2.400 793.800 35.370 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 1444.030 1496.880 1444.310 1497.160 ;
        RECT 1444.950 1496.880 1445.230 1497.160 ;
      LAYER met3 ;
        RECT 1444.005 1497.170 1444.335 1497.185 ;
        RECT 1444.925 1497.170 1445.255 1497.185 ;
        RECT 1444.005 1496.870 1445.255 1497.170 ;
        RECT 1444.005 1496.855 1444.335 1496.870 ;
        RECT 1444.925 1496.855 1445.255 1496.870 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1387.430 1678.140 1387.750 1678.200 ;
        RECT 1388.350 1678.140 1388.670 1678.200 ;
        RECT 1387.430 1678.000 1388.670 1678.140 ;
        RECT 1387.430 1677.940 1387.750 1678.000 ;
        RECT 1388.350 1677.940 1388.670 1678.000 ;
        RECT 641.310 59.400 641.630 59.460 ;
        RECT 1387.430 59.400 1387.750 59.460 ;
        RECT 641.310 59.260 1387.750 59.400 ;
        RECT 641.310 59.200 641.630 59.260 ;
        RECT 1387.430 59.200 1387.750 59.260 ;
      LAYER via ;
        RECT 1387.460 1677.940 1387.720 1678.200 ;
        RECT 1388.380 1677.940 1388.640 1678.200 ;
        RECT 641.340 59.200 641.600 59.460 ;
        RECT 1387.460 59.200 1387.720 59.460 ;
      LAYER met2 ;
        RECT 1390.145 1700.410 1390.425 1704.000 ;
        RECT 1388.440 1700.270 1390.425 1700.410 ;
        RECT 1388.440 1678.230 1388.580 1700.270 ;
        RECT 1390.145 1700.000 1390.425 1700.270 ;
        RECT 1387.460 1677.910 1387.720 1678.230 ;
        RECT 1388.380 1677.910 1388.640 1678.230 ;
        RECT 1387.520 59.490 1387.660 1677.910 ;
        RECT 641.340 59.170 641.600 59.490 ;
        RECT 1387.460 59.170 1387.720 59.490 ;
        RECT 641.400 17.410 641.540 59.170 ;
        RECT 639.100 17.270 641.540 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2063.170 1688.340 2063.490 1688.400 ;
        RECT 2069.610 1688.340 2069.930 1688.400 ;
        RECT 2063.170 1688.200 2069.930 1688.340 ;
        RECT 2063.170 1688.140 2063.490 1688.200 ;
        RECT 2069.610 1688.140 2069.930 1688.200 ;
        RECT 2069.610 34.240 2069.930 34.300 ;
        RECT 2422.890 34.240 2423.210 34.300 ;
        RECT 2069.610 34.100 2423.210 34.240 ;
        RECT 2069.610 34.040 2069.930 34.100 ;
        RECT 2422.890 34.040 2423.210 34.100 ;
      LAYER via ;
        RECT 2063.200 1688.140 2063.460 1688.400 ;
        RECT 2069.640 1688.140 2069.900 1688.400 ;
        RECT 2069.640 34.040 2069.900 34.300 ;
        RECT 2422.920 34.040 2423.180 34.300 ;
      LAYER met2 ;
        RECT 2063.125 1700.000 2063.405 1704.000 ;
        RECT 2063.260 1688.430 2063.400 1700.000 ;
        RECT 2063.200 1688.110 2063.460 1688.430 ;
        RECT 2069.640 1688.110 2069.900 1688.430 ;
        RECT 2069.700 34.330 2069.840 1688.110 ;
        RECT 2069.640 34.010 2069.900 34.330 ;
        RECT 2422.920 34.010 2423.180 34.330 ;
        RECT 2422.980 2.400 2423.120 34.010 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2070.070 1688.680 2070.390 1688.740 ;
        RECT 2076.510 1688.680 2076.830 1688.740 ;
        RECT 2070.070 1688.540 2076.830 1688.680 ;
        RECT 2070.070 1688.480 2070.390 1688.540 ;
        RECT 2076.510 1688.480 2076.830 1688.540 ;
        RECT 2076.510 33.900 2076.830 33.960 ;
        RECT 2440.830 33.900 2441.150 33.960 ;
        RECT 2076.510 33.760 2441.150 33.900 ;
        RECT 2076.510 33.700 2076.830 33.760 ;
        RECT 2440.830 33.700 2441.150 33.760 ;
      LAYER via ;
        RECT 2070.100 1688.480 2070.360 1688.740 ;
        RECT 2076.540 1688.480 2076.800 1688.740 ;
        RECT 2076.540 33.700 2076.800 33.960 ;
        RECT 2440.860 33.700 2441.120 33.960 ;
      LAYER met2 ;
        RECT 2070.025 1700.000 2070.305 1704.000 ;
        RECT 2070.160 1688.770 2070.300 1700.000 ;
        RECT 2070.100 1688.450 2070.360 1688.770 ;
        RECT 2076.540 1688.450 2076.800 1688.770 ;
        RECT 2076.600 33.990 2076.740 1688.450 ;
        RECT 2076.540 33.670 2076.800 33.990 ;
        RECT 2440.860 33.670 2441.120 33.990 ;
        RECT 2440.920 2.400 2441.060 33.670 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2076.970 1687.320 2077.290 1687.380 ;
        RECT 2082.950 1687.320 2083.270 1687.380 ;
        RECT 2076.970 1687.180 2083.270 1687.320 ;
        RECT 2076.970 1687.120 2077.290 1687.180 ;
        RECT 2082.950 1687.120 2083.270 1687.180 ;
        RECT 2082.950 33.560 2083.270 33.620 ;
        RECT 2458.770 33.560 2459.090 33.620 ;
        RECT 2082.950 33.420 2459.090 33.560 ;
        RECT 2082.950 33.360 2083.270 33.420 ;
        RECT 2458.770 33.360 2459.090 33.420 ;
      LAYER via ;
        RECT 2077.000 1687.120 2077.260 1687.380 ;
        RECT 2082.980 1687.120 2083.240 1687.380 ;
        RECT 2082.980 33.360 2083.240 33.620 ;
        RECT 2458.800 33.360 2459.060 33.620 ;
      LAYER met2 ;
        RECT 2076.925 1700.000 2077.205 1704.000 ;
        RECT 2077.060 1687.410 2077.200 1700.000 ;
        RECT 2077.000 1687.090 2077.260 1687.410 ;
        RECT 2082.980 1687.090 2083.240 1687.410 ;
        RECT 2083.040 33.650 2083.180 1687.090 ;
        RECT 2082.980 33.330 2083.240 33.650 ;
        RECT 2458.800 33.330 2459.060 33.650 ;
        RECT 2458.860 2.400 2459.000 33.330 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2083.410 33.220 2083.730 33.280 ;
        RECT 2476.710 33.220 2477.030 33.280 ;
        RECT 2083.410 33.080 2477.030 33.220 ;
        RECT 2083.410 33.020 2083.730 33.080 ;
        RECT 2476.710 33.020 2477.030 33.080 ;
      LAYER via ;
        RECT 2083.440 33.020 2083.700 33.280 ;
        RECT 2476.740 33.020 2477.000 33.280 ;
      LAYER met2 ;
        RECT 2083.365 1700.000 2083.645 1704.000 ;
        RECT 2083.500 33.310 2083.640 1700.000 ;
        RECT 2083.440 32.990 2083.700 33.310 ;
        RECT 2476.740 32.990 2477.000 33.310 ;
        RECT 2476.800 2.400 2476.940 32.990 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2090.310 32.880 2090.630 32.940 ;
        RECT 2494.650 32.880 2494.970 32.940 ;
        RECT 2090.310 32.740 2494.970 32.880 ;
        RECT 2090.310 32.680 2090.630 32.740 ;
        RECT 2494.650 32.680 2494.970 32.740 ;
      LAYER via ;
        RECT 2090.340 32.680 2090.600 32.940 ;
        RECT 2494.680 32.680 2494.940 32.940 ;
      LAYER met2 ;
        RECT 2090.265 1700.000 2090.545 1704.000 ;
        RECT 2090.400 32.970 2090.540 1700.000 ;
        RECT 2090.340 32.650 2090.600 32.970 ;
        RECT 2494.680 32.650 2494.940 32.970 ;
        RECT 2494.740 2.400 2494.880 32.650 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2097.210 32.540 2097.530 32.600 ;
        RECT 2512.130 32.540 2512.450 32.600 ;
        RECT 2097.210 32.400 2512.450 32.540 ;
        RECT 2097.210 32.340 2097.530 32.400 ;
        RECT 2512.130 32.340 2512.450 32.400 ;
      LAYER via ;
        RECT 2097.240 32.340 2097.500 32.600 ;
        RECT 2512.160 32.340 2512.420 32.600 ;
      LAYER met2 ;
        RECT 2097.165 1700.000 2097.445 1704.000 ;
        RECT 2097.300 32.630 2097.440 1700.000 ;
        RECT 2097.240 32.310 2097.500 32.630 ;
        RECT 2512.160 32.310 2512.420 32.630 ;
        RECT 2512.220 2.400 2512.360 32.310 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2104.110 32.200 2104.430 32.260 ;
        RECT 2530.070 32.200 2530.390 32.260 ;
        RECT 2104.110 32.060 2530.390 32.200 ;
        RECT 2104.110 32.000 2104.430 32.060 ;
        RECT 2530.070 32.000 2530.390 32.060 ;
      LAYER via ;
        RECT 2104.140 32.000 2104.400 32.260 ;
        RECT 2530.100 32.000 2530.360 32.260 ;
      LAYER met2 ;
        RECT 2103.605 1700.410 2103.885 1704.000 ;
        RECT 2103.605 1700.270 2104.340 1700.410 ;
        RECT 2103.605 1700.000 2103.885 1700.270 ;
        RECT 2104.200 32.290 2104.340 1700.270 ;
        RECT 2104.140 31.970 2104.400 32.290 ;
        RECT 2530.100 31.970 2530.360 32.290 ;
        RECT 2530.160 2.400 2530.300 31.970 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2111.010 31.860 2111.330 31.920 ;
        RECT 2548.010 31.860 2548.330 31.920 ;
        RECT 2111.010 31.720 2548.330 31.860 ;
        RECT 2111.010 31.660 2111.330 31.720 ;
        RECT 2548.010 31.660 2548.330 31.720 ;
      LAYER via ;
        RECT 2111.040 31.660 2111.300 31.920 ;
        RECT 2548.040 31.660 2548.300 31.920 ;
      LAYER met2 ;
        RECT 2110.505 1700.410 2110.785 1704.000 ;
        RECT 2110.505 1700.270 2111.240 1700.410 ;
        RECT 2110.505 1700.000 2110.785 1700.270 ;
        RECT 2111.100 31.950 2111.240 1700.270 ;
        RECT 2111.040 31.630 2111.300 31.950 ;
        RECT 2548.040 31.630 2548.300 31.950 ;
        RECT 2548.100 2.400 2548.240 31.630 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2117.450 31.520 2117.770 31.580 ;
        RECT 2565.950 31.520 2566.270 31.580 ;
        RECT 2117.450 31.380 2566.270 31.520 ;
        RECT 2117.450 31.320 2117.770 31.380 ;
        RECT 2565.950 31.320 2566.270 31.380 ;
      LAYER via ;
        RECT 2117.480 31.320 2117.740 31.580 ;
        RECT 2565.980 31.320 2566.240 31.580 ;
      LAYER met2 ;
        RECT 2117.405 1700.000 2117.685 1704.000 ;
        RECT 2117.540 31.610 2117.680 1700.000 ;
        RECT 2117.480 31.290 2117.740 31.610 ;
        RECT 2565.980 31.290 2566.240 31.610 ;
        RECT 2566.040 2.400 2566.180 31.290 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.350 31.180 2124.670 31.240 ;
        RECT 2583.890 31.180 2584.210 31.240 ;
        RECT 2124.350 31.040 2584.210 31.180 ;
        RECT 2124.350 30.980 2124.670 31.040 ;
        RECT 2583.890 30.980 2584.210 31.040 ;
      LAYER via ;
        RECT 2124.380 30.980 2124.640 31.240 ;
        RECT 2583.920 30.980 2584.180 31.240 ;
      LAYER met2 ;
        RECT 2123.845 1700.410 2124.125 1704.000 ;
        RECT 2123.845 1700.270 2124.580 1700.410 ;
        RECT 2123.845 1700.000 2124.125 1700.270 ;
        RECT 2124.440 31.270 2124.580 1700.270 ;
        RECT 2124.380 30.950 2124.640 31.270 ;
        RECT 2583.920 30.950 2584.180 31.270 ;
        RECT 2583.980 2.400 2584.120 30.950 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 33.220 817.810 33.280 ;
        RECT 1455.970 33.220 1456.290 33.280 ;
        RECT 817.490 33.080 1456.290 33.220 ;
        RECT 817.490 33.020 817.810 33.080 ;
        RECT 1455.970 33.020 1456.290 33.080 ;
      LAYER via ;
        RECT 817.520 33.020 817.780 33.280 ;
        RECT 1456.000 33.020 1456.260 33.280 ;
      LAYER met2 ;
        RECT 1457.305 1700.410 1457.585 1704.000 ;
        RECT 1456.060 1700.270 1457.585 1700.410 ;
        RECT 1456.060 33.310 1456.200 1700.270 ;
        RECT 1457.305 1700.000 1457.585 1700.270 ;
        RECT 817.520 32.990 817.780 33.310 ;
        RECT 1456.000 32.990 1456.260 33.310 ;
        RECT 817.580 2.400 817.720 32.990 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2131.250 30.840 2131.570 30.900 ;
        RECT 2601.370 30.840 2601.690 30.900 ;
        RECT 2131.250 30.700 2601.690 30.840 ;
        RECT 2131.250 30.640 2131.570 30.700 ;
        RECT 2601.370 30.640 2601.690 30.700 ;
      LAYER via ;
        RECT 2131.280 30.640 2131.540 30.900 ;
        RECT 2601.400 30.640 2601.660 30.900 ;
      LAYER met2 ;
        RECT 2130.745 1700.410 2131.025 1704.000 ;
        RECT 2130.745 1700.270 2131.480 1700.410 ;
        RECT 2130.745 1700.000 2131.025 1700.270 ;
        RECT 2131.340 30.930 2131.480 1700.270 ;
        RECT 2131.280 30.610 2131.540 30.930 ;
        RECT 2601.400 30.610 2601.660 30.930 ;
        RECT 2601.460 2.400 2601.600 30.610 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.150 40.700 2138.470 40.760 ;
        RECT 2619.310 40.700 2619.630 40.760 ;
        RECT 2138.150 40.560 2619.630 40.700 ;
        RECT 2138.150 40.500 2138.470 40.560 ;
        RECT 2619.310 40.500 2619.630 40.560 ;
      LAYER via ;
        RECT 2138.180 40.500 2138.440 40.760 ;
        RECT 2619.340 40.500 2619.600 40.760 ;
      LAYER met2 ;
        RECT 2137.645 1700.410 2137.925 1704.000 ;
        RECT 2137.645 1700.270 2138.380 1700.410 ;
        RECT 2137.645 1700.000 2137.925 1700.270 ;
        RECT 2138.240 40.790 2138.380 1700.270 ;
        RECT 2138.180 40.470 2138.440 40.790 ;
        RECT 2619.340 40.470 2619.600 40.790 ;
        RECT 2619.400 2.400 2619.540 40.470 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2145.050 40.360 2145.370 40.420 ;
        RECT 2637.250 40.360 2637.570 40.420 ;
        RECT 2145.050 40.220 2637.570 40.360 ;
        RECT 2145.050 40.160 2145.370 40.220 ;
        RECT 2637.250 40.160 2637.570 40.220 ;
      LAYER via ;
        RECT 2145.080 40.160 2145.340 40.420 ;
        RECT 2637.280 40.160 2637.540 40.420 ;
      LAYER met2 ;
        RECT 2144.085 1700.410 2144.365 1704.000 ;
        RECT 2144.085 1700.270 2145.280 1700.410 ;
        RECT 2144.085 1700.000 2144.365 1700.270 ;
        RECT 2145.140 40.450 2145.280 1700.270 ;
        RECT 2145.080 40.130 2145.340 40.450 ;
        RECT 2637.280 40.130 2637.540 40.450 ;
        RECT 2637.340 2.400 2637.480 40.130 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2151.950 40.020 2152.270 40.080 ;
        RECT 2655.190 40.020 2655.510 40.080 ;
        RECT 2151.950 39.880 2655.510 40.020 ;
        RECT 2151.950 39.820 2152.270 39.880 ;
        RECT 2655.190 39.820 2655.510 39.880 ;
      LAYER via ;
        RECT 2151.980 39.820 2152.240 40.080 ;
        RECT 2655.220 39.820 2655.480 40.080 ;
      LAYER met2 ;
        RECT 2150.985 1700.410 2151.265 1704.000 ;
        RECT 2150.985 1700.270 2152.180 1700.410 ;
        RECT 2150.985 1700.000 2151.265 1700.270 ;
        RECT 2152.040 40.110 2152.180 1700.270 ;
        RECT 2151.980 39.790 2152.240 40.110 ;
        RECT 2655.220 39.790 2655.480 40.110 ;
        RECT 2655.280 2.400 2655.420 39.790 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2158.850 39.680 2159.170 39.740 ;
        RECT 2672.670 39.680 2672.990 39.740 ;
        RECT 2158.850 39.540 2672.990 39.680 ;
        RECT 2158.850 39.480 2159.170 39.540 ;
        RECT 2672.670 39.480 2672.990 39.540 ;
      LAYER via ;
        RECT 2158.880 39.480 2159.140 39.740 ;
        RECT 2672.700 39.480 2672.960 39.740 ;
      LAYER met2 ;
        RECT 2157.425 1700.410 2157.705 1704.000 ;
        RECT 2157.425 1700.270 2159.080 1700.410 ;
        RECT 2157.425 1700.000 2157.705 1700.270 ;
        RECT 2158.940 39.770 2159.080 1700.270 ;
        RECT 2158.880 39.450 2159.140 39.770 ;
        RECT 2672.700 39.450 2672.960 39.770 ;
        RECT 2672.760 2.400 2672.900 39.450 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2165.750 39.340 2166.070 39.400 ;
        RECT 2690.610 39.340 2690.930 39.400 ;
        RECT 2165.750 39.200 2690.930 39.340 ;
        RECT 2165.750 39.140 2166.070 39.200 ;
        RECT 2690.610 39.140 2690.930 39.200 ;
      LAYER via ;
        RECT 2165.780 39.140 2166.040 39.400 ;
        RECT 2690.640 39.140 2690.900 39.400 ;
      LAYER met2 ;
        RECT 2164.325 1700.410 2164.605 1704.000 ;
        RECT 2164.325 1700.270 2165.980 1700.410 ;
        RECT 2164.325 1700.000 2164.605 1700.270 ;
        RECT 2165.840 39.430 2165.980 1700.270 ;
        RECT 2165.780 39.110 2166.040 39.430 ;
        RECT 2690.640 39.110 2690.900 39.430 ;
        RECT 2690.700 2.400 2690.840 39.110 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2171.345 1497.445 2171.515 1545.555 ;
        RECT 2171.345 1400.885 2171.515 1448.995 ;
        RECT 2171.345 1304.325 2171.515 1352.435 ;
        RECT 2171.345 1207.425 2171.515 1255.875 ;
        RECT 2171.345 1076.185 2171.515 1103.895 ;
        RECT 2172.265 966.025 2172.435 980.135 ;
        RECT 2172.265 772.905 2172.435 795.855 ;
        RECT 2172.265 689.605 2172.435 717.655 ;
        RECT 2171.805 476.085 2171.975 524.195 ;
        RECT 2171.805 435.625 2171.975 458.915 ;
        RECT 2171.345 331.585 2171.515 379.355 ;
        RECT 2172.265 145.265 2172.435 175.355 ;
        RECT 2173.185 89.845 2173.355 137.955 ;
      LAYER mcon ;
        RECT 2171.345 1545.385 2171.515 1545.555 ;
        RECT 2171.345 1448.825 2171.515 1448.995 ;
        RECT 2171.345 1352.265 2171.515 1352.435 ;
        RECT 2171.345 1255.705 2171.515 1255.875 ;
        RECT 2171.345 1103.725 2171.515 1103.895 ;
        RECT 2172.265 979.965 2172.435 980.135 ;
        RECT 2172.265 795.685 2172.435 795.855 ;
        RECT 2172.265 717.485 2172.435 717.655 ;
        RECT 2171.805 524.025 2171.975 524.195 ;
        RECT 2171.805 458.745 2171.975 458.915 ;
        RECT 2171.345 379.185 2171.515 379.355 ;
        RECT 2172.265 175.185 2172.435 175.355 ;
        RECT 2173.185 137.785 2173.355 137.955 ;
      LAYER met1 ;
        RECT 2171.730 1594.160 2172.050 1594.220 ;
        RECT 2172.190 1594.160 2172.510 1594.220 ;
        RECT 2171.730 1594.020 2172.510 1594.160 ;
        RECT 2171.730 1593.960 2172.050 1594.020 ;
        RECT 2172.190 1593.960 2172.510 1594.020 ;
        RECT 2171.285 1545.540 2171.575 1545.585 ;
        RECT 2172.650 1545.540 2172.970 1545.600 ;
        RECT 2171.285 1545.400 2172.970 1545.540 ;
        RECT 2171.285 1545.355 2171.575 1545.400 ;
        RECT 2172.650 1545.340 2172.970 1545.400 ;
        RECT 2171.270 1497.600 2171.590 1497.660 ;
        RECT 2171.075 1497.460 2171.590 1497.600 ;
        RECT 2171.270 1497.400 2171.590 1497.460 ;
        RECT 2171.285 1448.980 2171.575 1449.025 ;
        RECT 2171.730 1448.980 2172.050 1449.040 ;
        RECT 2171.285 1448.840 2172.050 1448.980 ;
        RECT 2171.285 1448.795 2171.575 1448.840 ;
        RECT 2171.730 1448.780 2172.050 1448.840 ;
        RECT 2171.270 1401.040 2171.590 1401.100 ;
        RECT 2171.075 1400.900 2171.590 1401.040 ;
        RECT 2171.270 1400.840 2171.590 1400.900 ;
        RECT 2171.285 1352.420 2171.575 1352.465 ;
        RECT 2171.730 1352.420 2172.050 1352.480 ;
        RECT 2171.285 1352.280 2172.050 1352.420 ;
        RECT 2171.285 1352.235 2171.575 1352.280 ;
        RECT 2171.730 1352.220 2172.050 1352.280 ;
        RECT 2171.270 1304.480 2171.590 1304.540 ;
        RECT 2171.075 1304.340 2171.590 1304.480 ;
        RECT 2171.270 1304.280 2171.590 1304.340 ;
        RECT 2171.285 1255.860 2171.575 1255.905 ;
        RECT 2171.730 1255.860 2172.050 1255.920 ;
        RECT 2171.285 1255.720 2172.050 1255.860 ;
        RECT 2171.285 1255.675 2171.575 1255.720 ;
        RECT 2171.730 1255.660 2172.050 1255.720 ;
        RECT 2171.270 1207.580 2171.590 1207.640 ;
        RECT 2171.075 1207.440 2171.590 1207.580 ;
        RECT 2171.270 1207.380 2171.590 1207.440 ;
        RECT 2171.270 1173.040 2171.590 1173.300 ;
        RECT 2171.360 1172.560 2171.500 1173.040 ;
        RECT 2171.730 1172.560 2172.050 1172.620 ;
        RECT 2171.360 1172.420 2172.050 1172.560 ;
        RECT 2171.730 1172.360 2172.050 1172.420 ;
        RECT 2171.730 1125.300 2172.050 1125.360 ;
        RECT 2171.360 1125.160 2172.050 1125.300 ;
        RECT 2171.360 1124.680 2171.500 1125.160 ;
        RECT 2171.730 1125.100 2172.050 1125.160 ;
        RECT 2171.270 1124.420 2171.590 1124.680 ;
        RECT 2171.270 1103.880 2171.590 1103.940 ;
        RECT 2171.075 1103.740 2171.590 1103.880 ;
        RECT 2171.270 1103.680 2171.590 1103.740 ;
        RECT 2171.270 1076.340 2171.590 1076.400 ;
        RECT 2171.075 1076.200 2171.590 1076.340 ;
        RECT 2171.270 1076.140 2171.590 1076.200 ;
        RECT 2171.730 1014.460 2172.050 1014.520 ;
        RECT 2172.650 1014.460 2172.970 1014.520 ;
        RECT 2171.730 1014.320 2172.970 1014.460 ;
        RECT 2171.730 1014.260 2172.050 1014.320 ;
        RECT 2172.650 1014.260 2172.970 1014.320 ;
        RECT 2172.190 980.120 2172.510 980.180 ;
        RECT 2171.995 979.980 2172.510 980.120 ;
        RECT 2172.190 979.920 2172.510 979.980 ;
        RECT 2172.190 966.180 2172.510 966.240 ;
        RECT 2171.995 966.040 2172.510 966.180 ;
        RECT 2172.190 965.980 2172.510 966.040 ;
        RECT 2172.190 918.240 2172.510 918.300 ;
        RECT 2171.360 918.100 2172.510 918.240 ;
        RECT 2171.360 917.960 2171.500 918.100 ;
        RECT 2172.190 918.040 2172.510 918.100 ;
        RECT 2171.270 917.700 2171.590 917.960 ;
        RECT 2172.190 795.840 2172.510 795.900 ;
        RECT 2171.995 795.700 2172.510 795.840 ;
        RECT 2172.190 795.640 2172.510 795.700 ;
        RECT 2172.190 773.060 2172.510 773.120 ;
        RECT 2171.995 772.920 2172.510 773.060 ;
        RECT 2172.190 772.860 2172.510 772.920 ;
        RECT 2172.190 738.040 2172.510 738.100 ;
        RECT 2173.570 738.040 2173.890 738.100 ;
        RECT 2172.190 737.900 2173.890 738.040 ;
        RECT 2172.190 737.840 2172.510 737.900 ;
        RECT 2173.570 737.840 2173.890 737.900 ;
        RECT 2172.190 717.640 2172.510 717.700 ;
        RECT 2171.995 717.500 2172.510 717.640 ;
        RECT 2172.190 717.440 2172.510 717.500 ;
        RECT 2172.205 689.760 2172.495 689.805 ;
        RECT 2172.650 689.760 2172.970 689.820 ;
        RECT 2172.205 689.620 2172.970 689.760 ;
        RECT 2172.205 689.575 2172.495 689.620 ;
        RECT 2172.650 689.560 2172.970 689.620 ;
        RECT 2171.730 545.060 2172.050 545.320 ;
        RECT 2171.820 544.920 2171.960 545.060 ;
        RECT 2172.190 544.920 2172.510 544.980 ;
        RECT 2171.820 544.780 2172.510 544.920 ;
        RECT 2172.190 544.720 2172.510 544.780 ;
        RECT 2171.745 524.180 2172.035 524.225 ;
        RECT 2172.190 524.180 2172.510 524.240 ;
        RECT 2171.745 524.040 2172.510 524.180 ;
        RECT 2171.745 523.995 2172.035 524.040 ;
        RECT 2172.190 523.980 2172.510 524.040 ;
        RECT 2171.730 476.240 2172.050 476.300 ;
        RECT 2171.535 476.100 2172.050 476.240 ;
        RECT 2171.730 476.040 2172.050 476.100 ;
        RECT 2171.730 458.900 2172.050 458.960 ;
        RECT 2171.535 458.760 2172.050 458.900 ;
        RECT 2171.730 458.700 2172.050 458.760 ;
        RECT 2171.745 435.780 2172.035 435.825 ;
        RECT 2172.650 435.780 2172.970 435.840 ;
        RECT 2171.745 435.640 2172.970 435.780 ;
        RECT 2171.745 435.595 2172.035 435.640 ;
        RECT 2172.650 435.580 2172.970 435.640 ;
        RECT 2171.285 379.340 2171.575 379.385 ;
        RECT 2171.730 379.340 2172.050 379.400 ;
        RECT 2171.285 379.200 2172.050 379.340 ;
        RECT 2171.285 379.155 2171.575 379.200 ;
        RECT 2171.730 379.140 2172.050 379.200 ;
        RECT 2171.270 331.740 2171.590 331.800 ;
        RECT 2171.075 331.600 2171.590 331.740 ;
        RECT 2171.270 331.540 2171.590 331.600 ;
        RECT 2171.270 330.860 2171.590 331.120 ;
        RECT 2171.360 330.720 2171.500 330.860 ;
        RECT 2172.190 330.720 2172.510 330.780 ;
        RECT 2171.360 330.580 2172.510 330.720 ;
        RECT 2172.190 330.520 2172.510 330.580 ;
        RECT 2171.730 255.580 2172.050 255.640 ;
        RECT 2171.360 255.440 2172.050 255.580 ;
        RECT 2171.360 255.300 2171.500 255.440 ;
        RECT 2171.730 255.380 2172.050 255.440 ;
        RECT 2171.270 255.040 2171.590 255.300 ;
        RECT 2172.190 175.340 2172.510 175.400 ;
        RECT 2171.995 175.200 2172.510 175.340 ;
        RECT 2172.190 175.140 2172.510 175.200 ;
        RECT 2172.205 145.420 2172.495 145.465 ;
        RECT 2172.650 145.420 2172.970 145.480 ;
        RECT 2172.205 145.280 2172.970 145.420 ;
        RECT 2172.205 145.235 2172.495 145.280 ;
        RECT 2172.650 145.220 2172.970 145.280 ;
        RECT 2172.650 137.940 2172.970 138.000 ;
        RECT 2173.125 137.940 2173.415 137.985 ;
        RECT 2172.650 137.800 2173.415 137.940 ;
        RECT 2172.650 137.740 2172.970 137.800 ;
        RECT 2173.125 137.755 2173.415 137.800 ;
        RECT 2172.650 90.000 2172.970 90.060 ;
        RECT 2173.125 90.000 2173.415 90.045 ;
        RECT 2172.650 89.860 2173.415 90.000 ;
        RECT 2172.650 89.800 2172.970 89.860 ;
        RECT 2173.125 89.815 2173.415 89.860 ;
        RECT 2172.650 85.040 2172.970 85.300 ;
        RECT 2172.740 84.280 2172.880 85.040 ;
        RECT 2172.650 84.020 2172.970 84.280 ;
        RECT 2172.650 39.000 2172.970 39.060 ;
        RECT 2708.550 39.000 2708.870 39.060 ;
        RECT 2172.650 38.860 2708.870 39.000 ;
        RECT 2172.650 38.800 2172.970 38.860 ;
        RECT 2708.550 38.800 2708.870 38.860 ;
      LAYER via ;
        RECT 2171.760 1593.960 2172.020 1594.220 ;
        RECT 2172.220 1593.960 2172.480 1594.220 ;
        RECT 2172.680 1545.340 2172.940 1545.600 ;
        RECT 2171.300 1497.400 2171.560 1497.660 ;
        RECT 2171.760 1448.780 2172.020 1449.040 ;
        RECT 2171.300 1400.840 2171.560 1401.100 ;
        RECT 2171.760 1352.220 2172.020 1352.480 ;
        RECT 2171.300 1304.280 2171.560 1304.540 ;
        RECT 2171.760 1255.660 2172.020 1255.920 ;
        RECT 2171.300 1207.380 2171.560 1207.640 ;
        RECT 2171.300 1173.040 2171.560 1173.300 ;
        RECT 2171.760 1172.360 2172.020 1172.620 ;
        RECT 2171.760 1125.100 2172.020 1125.360 ;
        RECT 2171.300 1124.420 2171.560 1124.680 ;
        RECT 2171.300 1103.680 2171.560 1103.940 ;
        RECT 2171.300 1076.140 2171.560 1076.400 ;
        RECT 2171.760 1014.260 2172.020 1014.520 ;
        RECT 2172.680 1014.260 2172.940 1014.520 ;
        RECT 2172.220 979.920 2172.480 980.180 ;
        RECT 2172.220 965.980 2172.480 966.240 ;
        RECT 2172.220 918.040 2172.480 918.300 ;
        RECT 2171.300 917.700 2171.560 917.960 ;
        RECT 2172.220 795.640 2172.480 795.900 ;
        RECT 2172.220 772.860 2172.480 773.120 ;
        RECT 2172.220 737.840 2172.480 738.100 ;
        RECT 2173.600 737.840 2173.860 738.100 ;
        RECT 2172.220 717.440 2172.480 717.700 ;
        RECT 2172.680 689.560 2172.940 689.820 ;
        RECT 2171.760 545.060 2172.020 545.320 ;
        RECT 2172.220 544.720 2172.480 544.980 ;
        RECT 2172.220 523.980 2172.480 524.240 ;
        RECT 2171.760 476.040 2172.020 476.300 ;
        RECT 2171.760 458.700 2172.020 458.960 ;
        RECT 2172.680 435.580 2172.940 435.840 ;
        RECT 2171.760 379.140 2172.020 379.400 ;
        RECT 2171.300 331.540 2171.560 331.800 ;
        RECT 2171.300 330.860 2171.560 331.120 ;
        RECT 2172.220 330.520 2172.480 330.780 ;
        RECT 2171.760 255.380 2172.020 255.640 ;
        RECT 2171.300 255.040 2171.560 255.300 ;
        RECT 2172.220 175.140 2172.480 175.400 ;
        RECT 2172.680 145.220 2172.940 145.480 ;
        RECT 2172.680 137.740 2172.940 138.000 ;
        RECT 2172.680 89.800 2172.940 90.060 ;
        RECT 2172.680 85.040 2172.940 85.300 ;
        RECT 2172.680 84.020 2172.940 84.280 ;
        RECT 2172.680 38.800 2172.940 39.060 ;
        RECT 2708.580 38.800 2708.840 39.060 ;
      LAYER met2 ;
        RECT 2171.225 1700.410 2171.505 1704.000 ;
        RECT 2171.225 1700.270 2172.420 1700.410 ;
        RECT 2171.225 1700.000 2171.505 1700.270 ;
        RECT 2172.280 1594.250 2172.420 1700.270 ;
        RECT 2171.760 1593.930 2172.020 1594.250 ;
        RECT 2172.220 1593.930 2172.480 1594.250 ;
        RECT 2171.820 1559.650 2171.960 1593.930 ;
        RECT 2171.820 1559.510 2172.880 1559.650 ;
        RECT 2172.740 1545.630 2172.880 1559.510 ;
        RECT 2172.680 1545.310 2172.940 1545.630 ;
        RECT 2171.300 1497.370 2171.560 1497.690 ;
        RECT 2171.360 1497.090 2171.500 1497.370 ;
        RECT 2171.750 1497.090 2172.030 1497.205 ;
        RECT 2171.360 1496.950 2172.030 1497.090 ;
        RECT 2171.750 1496.835 2172.030 1496.950 ;
        RECT 2171.750 1449.235 2172.030 1449.605 ;
        RECT 2171.820 1449.070 2171.960 1449.235 ;
        RECT 2171.760 1448.750 2172.020 1449.070 ;
        RECT 2171.300 1400.810 2171.560 1401.130 ;
        RECT 2171.360 1400.530 2171.500 1400.810 ;
        RECT 2171.750 1400.530 2172.030 1400.645 ;
        RECT 2171.360 1400.390 2172.030 1400.530 ;
        RECT 2171.750 1400.275 2172.030 1400.390 ;
        RECT 2171.750 1352.675 2172.030 1353.045 ;
        RECT 2171.820 1352.510 2171.960 1352.675 ;
        RECT 2171.760 1352.190 2172.020 1352.510 ;
        RECT 2171.300 1304.250 2171.560 1304.570 ;
        RECT 2171.360 1303.970 2171.500 1304.250 ;
        RECT 2171.750 1303.970 2172.030 1304.085 ;
        RECT 2171.360 1303.830 2172.030 1303.970 ;
        RECT 2171.750 1303.715 2172.030 1303.830 ;
        RECT 2171.750 1256.115 2172.030 1256.485 ;
        RECT 2171.820 1255.950 2171.960 1256.115 ;
        RECT 2171.760 1255.630 2172.020 1255.950 ;
        RECT 2171.300 1207.350 2171.560 1207.670 ;
        RECT 2171.360 1173.330 2171.500 1207.350 ;
        RECT 2171.300 1173.010 2171.560 1173.330 ;
        RECT 2171.760 1172.330 2172.020 1172.650 ;
        RECT 2171.820 1125.390 2171.960 1172.330 ;
        RECT 2171.760 1125.070 2172.020 1125.390 ;
        RECT 2171.300 1124.390 2171.560 1124.710 ;
        RECT 2171.360 1103.970 2171.500 1124.390 ;
        RECT 2171.300 1103.650 2171.560 1103.970 ;
        RECT 2171.300 1076.110 2171.560 1076.430 ;
        RECT 2171.360 1055.770 2171.500 1076.110 ;
        RECT 2171.360 1055.630 2171.960 1055.770 ;
        RECT 2171.820 1014.550 2171.960 1055.630 ;
        RECT 2172.740 1014.550 2172.880 1014.705 ;
        RECT 2171.760 1014.230 2172.020 1014.550 ;
        RECT 2172.680 1014.290 2172.940 1014.550 ;
        RECT 2172.280 1014.230 2172.940 1014.290 ;
        RECT 2172.280 1014.150 2172.880 1014.230 ;
        RECT 2172.280 980.210 2172.420 1014.150 ;
        RECT 2172.220 979.890 2172.480 980.210 ;
        RECT 2172.220 965.950 2172.480 966.270 ;
        RECT 2172.280 918.330 2172.420 965.950 ;
        RECT 2172.220 918.010 2172.480 918.330 ;
        RECT 2171.300 917.670 2171.560 917.990 ;
        RECT 2171.360 869.450 2171.500 917.670 ;
        RECT 2171.750 869.450 2172.030 869.565 ;
        RECT 2171.360 869.310 2172.030 869.450 ;
        RECT 2171.750 869.195 2172.030 869.310 ;
        RECT 2172.210 820.915 2172.490 821.285 ;
        RECT 2172.280 795.930 2172.420 820.915 ;
        RECT 2172.220 795.610 2172.480 795.930 ;
        RECT 2172.220 772.830 2172.480 773.150 ;
        RECT 2172.280 738.130 2172.420 772.830 ;
        RECT 2172.220 737.810 2172.480 738.130 ;
        RECT 2173.600 737.810 2173.860 738.130 ;
        RECT 2173.660 717.925 2173.800 737.810 ;
        RECT 2172.670 717.810 2172.950 717.925 ;
        RECT 2172.280 717.730 2172.950 717.810 ;
        RECT 2172.220 717.670 2172.950 717.730 ;
        RECT 2172.220 717.410 2172.480 717.670 ;
        RECT 2172.670 717.555 2172.950 717.670 ;
        RECT 2173.590 717.555 2173.870 717.925 ;
        RECT 2172.680 689.530 2172.940 689.850 ;
        RECT 2172.740 643.010 2172.880 689.530 ;
        RECT 2172.280 642.870 2172.880 643.010 ;
        RECT 2172.280 603.570 2172.420 642.870 ;
        RECT 2171.820 603.430 2172.420 603.570 ;
        RECT 2171.820 545.350 2171.960 603.430 ;
        RECT 2171.760 545.030 2172.020 545.350 ;
        RECT 2172.220 544.690 2172.480 545.010 ;
        RECT 2172.280 524.270 2172.420 544.690 ;
        RECT 2172.220 523.950 2172.480 524.270 ;
        RECT 2171.760 476.010 2172.020 476.330 ;
        RECT 2171.820 458.990 2171.960 476.010 ;
        RECT 2171.760 458.670 2172.020 458.990 ;
        RECT 2172.680 435.550 2172.940 435.870 ;
        RECT 2172.740 400.250 2172.880 435.550 ;
        RECT 2171.820 400.110 2172.880 400.250 ;
        RECT 2171.820 379.430 2171.960 400.110 ;
        RECT 2171.760 379.110 2172.020 379.430 ;
        RECT 2171.300 331.510 2171.560 331.830 ;
        RECT 2171.360 331.150 2171.500 331.510 ;
        RECT 2171.300 330.830 2171.560 331.150 ;
        RECT 2172.220 330.490 2172.480 330.810 ;
        RECT 2172.280 303.010 2172.420 330.490 ;
        RECT 2171.820 302.870 2172.420 303.010 ;
        RECT 2171.820 255.670 2171.960 302.870 ;
        RECT 2171.760 255.350 2172.020 255.670 ;
        RECT 2171.300 255.010 2171.560 255.330 ;
        RECT 2171.360 241.245 2171.500 255.010 ;
        RECT 2171.290 240.875 2171.570 241.245 ;
        RECT 2172.210 206.195 2172.490 206.565 ;
        RECT 2172.280 175.430 2172.420 206.195 ;
        RECT 2172.220 175.110 2172.480 175.430 ;
        RECT 2172.680 145.190 2172.940 145.510 ;
        RECT 2172.740 138.030 2172.880 145.190 ;
        RECT 2172.680 137.710 2172.940 138.030 ;
        RECT 2172.680 89.770 2172.940 90.090 ;
        RECT 2172.740 85.330 2172.880 89.770 ;
        RECT 2172.680 85.010 2172.940 85.330 ;
        RECT 2172.680 83.990 2172.940 84.310 ;
        RECT 2172.740 39.090 2172.880 83.990 ;
        RECT 2172.680 38.770 2172.940 39.090 ;
        RECT 2708.580 38.770 2708.840 39.090 ;
        RECT 2708.640 2.400 2708.780 38.770 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
      LAYER via2 ;
        RECT 2171.750 1496.880 2172.030 1497.160 ;
        RECT 2171.750 1449.280 2172.030 1449.560 ;
        RECT 2171.750 1400.320 2172.030 1400.600 ;
        RECT 2171.750 1352.720 2172.030 1353.000 ;
        RECT 2171.750 1303.760 2172.030 1304.040 ;
        RECT 2171.750 1256.160 2172.030 1256.440 ;
        RECT 2171.750 869.240 2172.030 869.520 ;
        RECT 2172.210 820.960 2172.490 821.240 ;
        RECT 2172.670 717.600 2172.950 717.880 ;
        RECT 2173.590 717.600 2173.870 717.880 ;
        RECT 2171.290 240.920 2171.570 241.200 ;
        RECT 2172.210 206.240 2172.490 206.520 ;
      LAYER met3 ;
        RECT 2171.725 1497.170 2172.055 1497.185 ;
        RECT 2172.390 1497.170 2172.770 1497.180 ;
        RECT 2171.725 1496.870 2172.770 1497.170 ;
        RECT 2171.725 1496.855 2172.055 1496.870 ;
        RECT 2172.390 1496.860 2172.770 1496.870 ;
        RECT 2171.725 1449.570 2172.055 1449.585 ;
        RECT 2172.390 1449.570 2172.770 1449.580 ;
        RECT 2171.725 1449.270 2172.770 1449.570 ;
        RECT 2171.725 1449.255 2172.055 1449.270 ;
        RECT 2172.390 1449.260 2172.770 1449.270 ;
        RECT 2171.725 1400.610 2172.055 1400.625 ;
        RECT 2172.390 1400.610 2172.770 1400.620 ;
        RECT 2171.725 1400.310 2172.770 1400.610 ;
        RECT 2171.725 1400.295 2172.055 1400.310 ;
        RECT 2172.390 1400.300 2172.770 1400.310 ;
        RECT 2171.725 1353.010 2172.055 1353.025 ;
        RECT 2172.390 1353.010 2172.770 1353.020 ;
        RECT 2171.725 1352.710 2172.770 1353.010 ;
        RECT 2171.725 1352.695 2172.055 1352.710 ;
        RECT 2172.390 1352.700 2172.770 1352.710 ;
        RECT 2171.725 1304.050 2172.055 1304.065 ;
        RECT 2172.390 1304.050 2172.770 1304.060 ;
        RECT 2171.725 1303.750 2172.770 1304.050 ;
        RECT 2171.725 1303.735 2172.055 1303.750 ;
        RECT 2172.390 1303.740 2172.770 1303.750 ;
        RECT 2171.725 1256.450 2172.055 1256.465 ;
        RECT 2172.390 1256.450 2172.770 1256.460 ;
        RECT 2171.725 1256.150 2172.770 1256.450 ;
        RECT 2171.725 1256.135 2172.055 1256.150 ;
        RECT 2172.390 1256.140 2172.770 1256.150 ;
        RECT 2171.725 869.540 2172.055 869.545 ;
        RECT 2171.470 869.530 2172.055 869.540 ;
        RECT 2171.470 869.230 2172.280 869.530 ;
        RECT 2171.470 869.220 2172.055 869.230 ;
        RECT 2171.725 869.215 2172.055 869.220 ;
        RECT 2171.470 821.250 2171.850 821.260 ;
        RECT 2172.185 821.250 2172.515 821.265 ;
        RECT 2171.470 820.950 2172.515 821.250 ;
        RECT 2171.470 820.940 2171.850 820.950 ;
        RECT 2172.185 820.935 2172.515 820.950 ;
        RECT 2172.645 717.890 2172.975 717.905 ;
        RECT 2173.565 717.890 2173.895 717.905 ;
        RECT 2172.645 717.590 2173.895 717.890 ;
        RECT 2172.645 717.575 2172.975 717.590 ;
        RECT 2173.565 717.575 2173.895 717.590 ;
        RECT 2171.265 241.220 2171.595 241.225 ;
        RECT 2171.265 241.210 2171.850 241.220 ;
        RECT 2171.265 240.910 2172.050 241.210 ;
        RECT 2171.265 240.900 2171.850 240.910 ;
        RECT 2171.265 240.895 2171.595 240.900 ;
        RECT 2171.470 206.530 2171.850 206.540 ;
        RECT 2172.185 206.530 2172.515 206.545 ;
        RECT 2171.470 206.230 2172.515 206.530 ;
        RECT 2171.470 206.220 2171.850 206.230 ;
        RECT 2172.185 206.215 2172.515 206.230 ;
      LAYER via3 ;
        RECT 2172.420 1496.860 2172.740 1497.180 ;
        RECT 2172.420 1449.260 2172.740 1449.580 ;
        RECT 2172.420 1400.300 2172.740 1400.620 ;
        RECT 2172.420 1352.700 2172.740 1353.020 ;
        RECT 2172.420 1303.740 2172.740 1304.060 ;
        RECT 2172.420 1256.140 2172.740 1256.460 ;
        RECT 2171.500 869.220 2171.820 869.540 ;
        RECT 2171.500 820.940 2171.820 821.260 ;
        RECT 2171.500 240.900 2171.820 241.220 ;
        RECT 2171.500 206.220 2171.820 206.540 ;
      LAYER met4 ;
        RECT 2172.415 1496.855 2172.745 1497.185 ;
        RECT 2172.430 1449.585 2172.730 1496.855 ;
        RECT 2172.415 1449.255 2172.745 1449.585 ;
        RECT 2172.415 1400.295 2172.745 1400.625 ;
        RECT 2172.430 1353.025 2172.730 1400.295 ;
        RECT 2172.415 1352.695 2172.745 1353.025 ;
        RECT 2172.415 1303.735 2172.745 1304.065 ;
        RECT 2172.430 1256.465 2172.730 1303.735 ;
        RECT 2172.415 1256.135 2172.745 1256.465 ;
        RECT 2171.495 869.215 2171.825 869.545 ;
        RECT 2171.510 821.265 2171.810 869.215 ;
        RECT 2171.495 820.935 2171.825 821.265 ;
        RECT 2171.495 240.895 2171.825 241.225 ;
        RECT 2171.510 206.545 2171.810 240.895 ;
        RECT 2171.495 206.215 2171.825 206.545 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2179.550 38.660 2179.870 38.720 ;
        RECT 2726.490 38.660 2726.810 38.720 ;
        RECT 2179.550 38.520 2726.810 38.660 ;
        RECT 2179.550 38.460 2179.870 38.520 ;
        RECT 2726.490 38.460 2726.810 38.520 ;
      LAYER via ;
        RECT 2179.580 38.460 2179.840 38.720 ;
        RECT 2726.520 38.460 2726.780 38.720 ;
      LAYER met2 ;
        RECT 2177.665 1700.410 2177.945 1704.000 ;
        RECT 2177.665 1700.270 2179.780 1700.410 ;
        RECT 2177.665 1700.000 2177.945 1700.270 ;
        RECT 2179.640 38.750 2179.780 1700.270 ;
        RECT 2179.580 38.430 2179.840 38.750 ;
        RECT 2726.520 38.430 2726.780 38.750 ;
        RECT 2726.580 2.400 2726.720 38.430 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2186.450 38.320 2186.770 38.380 ;
        RECT 2744.430 38.320 2744.750 38.380 ;
        RECT 2186.450 38.180 2744.750 38.320 ;
        RECT 2186.450 38.120 2186.770 38.180 ;
        RECT 2744.430 38.120 2744.750 38.180 ;
      LAYER via ;
        RECT 2186.480 38.120 2186.740 38.380 ;
        RECT 2744.460 38.120 2744.720 38.380 ;
      LAYER met2 ;
        RECT 2184.565 1700.410 2184.845 1704.000 ;
        RECT 2184.565 1700.270 2186.680 1700.410 ;
        RECT 2184.565 1700.000 2184.845 1700.270 ;
        RECT 2186.540 38.410 2186.680 1700.270 ;
        RECT 2186.480 38.090 2186.740 38.410 ;
        RECT 2744.460 38.090 2744.720 38.410 ;
        RECT 2744.520 2.400 2744.660 38.090 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2193.350 37.980 2193.670 38.040 ;
        RECT 2761.910 37.980 2762.230 38.040 ;
        RECT 2193.350 37.840 2762.230 37.980 ;
        RECT 2193.350 37.780 2193.670 37.840 ;
        RECT 2761.910 37.780 2762.230 37.840 ;
      LAYER via ;
        RECT 2193.380 37.780 2193.640 38.040 ;
        RECT 2761.940 37.780 2762.200 38.040 ;
      LAYER met2 ;
        RECT 2191.465 1700.410 2191.745 1704.000 ;
        RECT 2191.465 1700.270 2193.580 1700.410 ;
        RECT 2191.465 1700.000 2191.745 1700.270 ;
        RECT 2193.440 38.070 2193.580 1700.270 ;
        RECT 2193.380 37.750 2193.640 38.070 ;
        RECT 2761.940 37.750 2762.200 38.070 ;
        RECT 2762.000 2.400 2762.140 37.750 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 835.430 33.560 835.750 33.620 ;
        RECT 1462.870 33.560 1463.190 33.620 ;
        RECT 835.430 33.420 1463.190 33.560 ;
        RECT 835.430 33.360 835.750 33.420 ;
        RECT 1462.870 33.360 1463.190 33.420 ;
      LAYER via ;
        RECT 835.460 33.360 835.720 33.620 ;
        RECT 1462.900 33.360 1463.160 33.620 ;
      LAYER met2 ;
        RECT 1464.205 1700.410 1464.485 1704.000 ;
        RECT 1462.960 1700.270 1464.485 1700.410 ;
        RECT 1462.960 33.650 1463.100 1700.270 ;
        RECT 1464.205 1700.000 1464.485 1700.270 ;
        RECT 835.460 33.330 835.720 33.650 ;
        RECT 1462.900 33.330 1463.160 33.650 ;
        RECT 835.520 2.400 835.660 33.330 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2199.790 47.160 2200.110 47.220 ;
        RECT 2779.850 47.160 2780.170 47.220 ;
        RECT 2199.790 47.020 2780.170 47.160 ;
        RECT 2199.790 46.960 2200.110 47.020 ;
        RECT 2779.850 46.960 2780.170 47.020 ;
      LAYER via ;
        RECT 2199.820 46.960 2200.080 47.220 ;
        RECT 2779.880 46.960 2780.140 47.220 ;
      LAYER met2 ;
        RECT 2197.905 1700.410 2198.185 1704.000 ;
        RECT 2197.905 1700.270 2200.020 1700.410 ;
        RECT 2197.905 1700.000 2198.185 1700.270 ;
        RECT 2199.880 47.250 2200.020 1700.270 ;
        RECT 2199.820 46.930 2200.080 47.250 ;
        RECT 2779.880 46.930 2780.140 47.250 ;
        RECT 2779.940 2.400 2780.080 46.930 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2207.150 46.820 2207.470 46.880 ;
        RECT 2797.790 46.820 2798.110 46.880 ;
        RECT 2207.150 46.680 2798.110 46.820 ;
        RECT 2207.150 46.620 2207.470 46.680 ;
        RECT 2797.790 46.620 2798.110 46.680 ;
      LAYER via ;
        RECT 2207.180 46.620 2207.440 46.880 ;
        RECT 2797.820 46.620 2798.080 46.880 ;
      LAYER met2 ;
        RECT 2204.805 1700.410 2205.085 1704.000 ;
        RECT 2204.805 1700.270 2206.460 1700.410 ;
        RECT 2204.805 1700.000 2205.085 1700.270 ;
        RECT 2206.320 1677.970 2206.460 1700.270 ;
        RECT 2206.320 1677.830 2207.380 1677.970 ;
        RECT 2207.240 46.910 2207.380 1677.830 ;
        RECT 2207.180 46.590 2207.440 46.910 ;
        RECT 2797.820 46.590 2798.080 46.910 ;
        RECT 2797.880 2.400 2798.020 46.590 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2213.590 46.480 2213.910 46.540 ;
        RECT 2815.730 46.480 2816.050 46.540 ;
        RECT 2213.590 46.340 2816.050 46.480 ;
        RECT 2213.590 46.280 2213.910 46.340 ;
        RECT 2815.730 46.280 2816.050 46.340 ;
      LAYER via ;
        RECT 2213.620 46.280 2213.880 46.540 ;
        RECT 2815.760 46.280 2816.020 46.540 ;
      LAYER met2 ;
        RECT 2211.705 1700.410 2211.985 1704.000 ;
        RECT 2211.705 1700.270 2212.900 1700.410 ;
        RECT 2211.705 1700.000 2211.985 1700.270 ;
        RECT 2212.760 1666.410 2212.900 1700.270 ;
        RECT 2212.760 1666.270 2213.820 1666.410 ;
        RECT 2213.680 46.570 2213.820 1666.270 ;
        RECT 2213.620 46.250 2213.880 46.570 ;
        RECT 2815.760 46.250 2816.020 46.570 ;
        RECT 2815.820 2.400 2815.960 46.250 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2220.565 786.505 2220.735 821.015 ;
        RECT 2220.565 724.965 2220.735 772.735 ;
        RECT 2220.565 641.325 2220.735 717.655 ;
        RECT 2221.025 593.045 2221.195 627.895 ;
        RECT 2220.565 496.485 2220.735 531.335 ;
        RECT 2220.565 386.325 2220.735 434.775 ;
        RECT 2220.565 193.205 2220.735 241.315 ;
        RECT 2220.565 144.925 2220.735 159.375 ;
      LAYER mcon ;
        RECT 2220.565 820.845 2220.735 821.015 ;
        RECT 2220.565 772.565 2220.735 772.735 ;
        RECT 2220.565 717.485 2220.735 717.655 ;
        RECT 2221.025 627.725 2221.195 627.895 ;
        RECT 2220.565 531.165 2220.735 531.335 ;
        RECT 2220.565 434.605 2220.735 434.775 ;
        RECT 2220.565 241.145 2220.735 241.315 ;
        RECT 2220.565 159.205 2220.735 159.375 ;
      LAYER met1 ;
        RECT 2220.490 1594.160 2220.810 1594.220 ;
        RECT 2220.950 1594.160 2221.270 1594.220 ;
        RECT 2220.490 1594.020 2221.270 1594.160 ;
        RECT 2220.490 1593.960 2220.810 1594.020 ;
        RECT 2220.950 1593.960 2221.270 1594.020 ;
        RECT 2220.490 1559.820 2220.810 1559.880 ;
        RECT 2220.950 1559.820 2221.270 1559.880 ;
        RECT 2220.490 1559.680 2221.270 1559.820 ;
        RECT 2220.490 1559.620 2220.810 1559.680 ;
        RECT 2220.950 1559.620 2221.270 1559.680 ;
        RECT 2220.030 1511.200 2220.350 1511.260 ;
        RECT 2220.950 1511.200 2221.270 1511.260 ;
        RECT 2220.030 1511.060 2221.270 1511.200 ;
        RECT 2220.030 1511.000 2220.350 1511.060 ;
        RECT 2220.950 1511.000 2221.270 1511.060 ;
        RECT 2220.030 1414.640 2220.350 1414.700 ;
        RECT 2220.950 1414.640 2221.270 1414.700 ;
        RECT 2220.030 1414.500 2221.270 1414.640 ;
        RECT 2220.030 1414.440 2220.350 1414.500 ;
        RECT 2220.950 1414.440 2221.270 1414.500 ;
        RECT 2220.030 1318.080 2220.350 1318.140 ;
        RECT 2220.950 1318.080 2221.270 1318.140 ;
        RECT 2220.030 1317.940 2221.270 1318.080 ;
        RECT 2220.030 1317.880 2220.350 1317.940 ;
        RECT 2220.950 1317.880 2221.270 1317.940 ;
        RECT 2220.030 1221.520 2220.350 1221.580 ;
        RECT 2220.950 1221.520 2221.270 1221.580 ;
        RECT 2220.030 1221.380 2221.270 1221.520 ;
        RECT 2220.030 1221.320 2220.350 1221.380 ;
        RECT 2220.950 1221.320 2221.270 1221.380 ;
        RECT 2220.030 1124.960 2220.350 1125.020 ;
        RECT 2220.950 1124.960 2221.270 1125.020 ;
        RECT 2220.030 1124.820 2221.270 1124.960 ;
        RECT 2220.030 1124.760 2220.350 1124.820 ;
        RECT 2220.950 1124.760 2221.270 1124.820 ;
        RECT 2220.030 1028.400 2220.350 1028.460 ;
        RECT 2220.950 1028.400 2221.270 1028.460 ;
        RECT 2220.030 1028.260 2221.270 1028.400 ;
        RECT 2220.030 1028.200 2220.350 1028.260 ;
        RECT 2220.950 1028.200 2221.270 1028.260 ;
        RECT 2220.030 931.840 2220.350 931.900 ;
        RECT 2220.950 931.840 2221.270 931.900 ;
        RECT 2220.030 931.700 2221.270 931.840 ;
        RECT 2220.030 931.640 2220.350 931.700 ;
        RECT 2220.950 931.640 2221.270 931.700 ;
        RECT 2219.570 869.620 2219.890 869.680 ;
        RECT 2220.490 869.620 2220.810 869.680 ;
        RECT 2219.570 869.480 2220.810 869.620 ;
        RECT 2219.570 869.420 2219.890 869.480 ;
        RECT 2220.490 869.420 2220.810 869.480 ;
        RECT 2220.490 821.000 2220.810 821.060 ;
        RECT 2220.295 820.860 2220.810 821.000 ;
        RECT 2220.490 820.800 2220.810 820.860 ;
        RECT 2220.490 786.660 2220.810 786.720 ;
        RECT 2220.295 786.520 2220.810 786.660 ;
        RECT 2220.490 786.460 2220.810 786.520 ;
        RECT 2220.505 772.720 2220.795 772.765 ;
        RECT 2220.950 772.720 2221.270 772.780 ;
        RECT 2220.505 772.580 2221.270 772.720 ;
        RECT 2220.505 772.535 2220.795 772.580 ;
        RECT 2220.950 772.520 2221.270 772.580 ;
        RECT 2220.490 725.120 2220.810 725.180 ;
        RECT 2220.295 724.980 2220.810 725.120 ;
        RECT 2220.490 724.920 2220.810 724.980 ;
        RECT 2220.490 717.640 2220.810 717.700 ;
        RECT 2220.295 717.500 2220.810 717.640 ;
        RECT 2220.490 717.440 2220.810 717.500 ;
        RECT 2220.490 641.480 2220.810 641.540 ;
        RECT 2220.295 641.340 2220.810 641.480 ;
        RECT 2220.490 641.280 2220.810 641.340 ;
        RECT 2220.490 627.880 2220.810 627.940 ;
        RECT 2220.965 627.880 2221.255 627.925 ;
        RECT 2220.490 627.740 2221.255 627.880 ;
        RECT 2220.490 627.680 2220.810 627.740 ;
        RECT 2220.965 627.695 2221.255 627.740 ;
        RECT 2220.950 593.200 2221.270 593.260 ;
        RECT 2220.755 593.060 2221.270 593.200 ;
        RECT 2220.950 593.000 2221.270 593.060 ;
        RECT 2220.030 545.260 2220.350 545.320 ;
        RECT 2220.950 545.260 2221.270 545.320 ;
        RECT 2220.030 545.120 2221.270 545.260 ;
        RECT 2220.030 545.060 2220.350 545.120 ;
        RECT 2220.950 545.060 2221.270 545.120 ;
        RECT 2220.490 531.320 2220.810 531.380 ;
        RECT 2220.295 531.180 2220.810 531.320 ;
        RECT 2220.490 531.120 2220.810 531.180 ;
        RECT 2220.490 496.640 2220.810 496.700 ;
        RECT 2220.295 496.500 2220.810 496.640 ;
        RECT 2220.490 496.440 2220.810 496.500 ;
        RECT 2220.030 448.700 2220.350 448.760 ;
        RECT 2220.950 448.700 2221.270 448.760 ;
        RECT 2220.030 448.560 2221.270 448.700 ;
        RECT 2220.030 448.500 2220.350 448.560 ;
        RECT 2220.950 448.500 2221.270 448.560 ;
        RECT 2220.490 434.760 2220.810 434.820 ;
        RECT 2220.295 434.620 2220.810 434.760 ;
        RECT 2220.490 434.560 2220.810 434.620 ;
        RECT 2220.505 386.480 2220.795 386.525 ;
        RECT 2220.950 386.480 2221.270 386.540 ;
        RECT 2220.505 386.340 2221.270 386.480 ;
        RECT 2220.505 386.295 2220.795 386.340 ;
        RECT 2220.950 386.280 2221.270 386.340 ;
        RECT 2220.490 338.200 2220.810 338.260 ;
        RECT 2220.950 338.200 2221.270 338.260 ;
        RECT 2220.490 338.060 2221.270 338.200 ;
        RECT 2220.490 338.000 2220.810 338.060 ;
        RECT 2220.950 338.000 2221.270 338.060 ;
        RECT 2220.490 304.200 2220.810 304.260 ;
        RECT 2220.120 304.060 2220.810 304.200 ;
        RECT 2220.120 303.580 2220.260 304.060 ;
        RECT 2220.490 304.000 2220.810 304.060 ;
        RECT 2220.030 303.320 2220.350 303.580 ;
        RECT 2220.030 255.240 2220.350 255.300 ;
        RECT 2220.950 255.240 2221.270 255.300 ;
        RECT 2220.030 255.100 2221.270 255.240 ;
        RECT 2220.030 255.040 2220.350 255.100 ;
        RECT 2220.950 255.040 2221.270 255.100 ;
        RECT 2220.505 241.300 2220.795 241.345 ;
        RECT 2220.950 241.300 2221.270 241.360 ;
        RECT 2220.505 241.160 2221.270 241.300 ;
        RECT 2220.505 241.115 2220.795 241.160 ;
        RECT 2220.950 241.100 2221.270 241.160 ;
        RECT 2220.490 193.360 2220.810 193.420 ;
        RECT 2220.295 193.220 2220.810 193.360 ;
        RECT 2220.490 193.160 2220.810 193.220 ;
        RECT 2220.490 159.360 2220.810 159.420 ;
        RECT 2220.295 159.220 2220.810 159.360 ;
        RECT 2220.490 159.160 2220.810 159.220 ;
        RECT 2220.490 145.080 2220.810 145.140 ;
        RECT 2220.295 144.940 2220.810 145.080 ;
        RECT 2220.490 144.880 2220.810 144.940 ;
        RECT 2220.030 46.140 2220.350 46.200 ;
        RECT 2833.670 46.140 2833.990 46.200 ;
        RECT 2220.030 46.000 2833.990 46.140 ;
        RECT 2220.030 45.940 2220.350 46.000 ;
        RECT 2833.670 45.940 2833.990 46.000 ;
      LAYER via ;
        RECT 2220.520 1593.960 2220.780 1594.220 ;
        RECT 2220.980 1593.960 2221.240 1594.220 ;
        RECT 2220.520 1559.620 2220.780 1559.880 ;
        RECT 2220.980 1559.620 2221.240 1559.880 ;
        RECT 2220.060 1511.000 2220.320 1511.260 ;
        RECT 2220.980 1511.000 2221.240 1511.260 ;
        RECT 2220.060 1414.440 2220.320 1414.700 ;
        RECT 2220.980 1414.440 2221.240 1414.700 ;
        RECT 2220.060 1317.880 2220.320 1318.140 ;
        RECT 2220.980 1317.880 2221.240 1318.140 ;
        RECT 2220.060 1221.320 2220.320 1221.580 ;
        RECT 2220.980 1221.320 2221.240 1221.580 ;
        RECT 2220.060 1124.760 2220.320 1125.020 ;
        RECT 2220.980 1124.760 2221.240 1125.020 ;
        RECT 2220.060 1028.200 2220.320 1028.460 ;
        RECT 2220.980 1028.200 2221.240 1028.460 ;
        RECT 2220.060 931.640 2220.320 931.900 ;
        RECT 2220.980 931.640 2221.240 931.900 ;
        RECT 2219.600 869.420 2219.860 869.680 ;
        RECT 2220.520 869.420 2220.780 869.680 ;
        RECT 2220.520 820.800 2220.780 821.060 ;
        RECT 2220.520 786.460 2220.780 786.720 ;
        RECT 2220.980 772.520 2221.240 772.780 ;
        RECT 2220.520 724.920 2220.780 725.180 ;
        RECT 2220.520 717.440 2220.780 717.700 ;
        RECT 2220.520 641.280 2220.780 641.540 ;
        RECT 2220.520 627.680 2220.780 627.940 ;
        RECT 2220.980 593.000 2221.240 593.260 ;
        RECT 2220.060 545.060 2220.320 545.320 ;
        RECT 2220.980 545.060 2221.240 545.320 ;
        RECT 2220.520 531.120 2220.780 531.380 ;
        RECT 2220.520 496.440 2220.780 496.700 ;
        RECT 2220.060 448.500 2220.320 448.760 ;
        RECT 2220.980 448.500 2221.240 448.760 ;
        RECT 2220.520 434.560 2220.780 434.820 ;
        RECT 2220.980 386.280 2221.240 386.540 ;
        RECT 2220.520 338.000 2220.780 338.260 ;
        RECT 2220.980 338.000 2221.240 338.260 ;
        RECT 2220.520 304.000 2220.780 304.260 ;
        RECT 2220.060 303.320 2220.320 303.580 ;
        RECT 2220.060 255.040 2220.320 255.300 ;
        RECT 2220.980 255.040 2221.240 255.300 ;
        RECT 2220.980 241.100 2221.240 241.360 ;
        RECT 2220.520 193.160 2220.780 193.420 ;
        RECT 2220.520 159.160 2220.780 159.420 ;
        RECT 2220.520 144.880 2220.780 145.140 ;
        RECT 2220.060 45.940 2220.320 46.200 ;
        RECT 2833.700 45.940 2833.960 46.200 ;
      LAYER met2 ;
        RECT 2218.145 1700.410 2218.425 1704.000 ;
        RECT 2218.145 1700.270 2219.800 1700.410 ;
        RECT 2218.145 1700.000 2218.425 1700.270 ;
        RECT 2219.660 1677.970 2219.800 1700.270 ;
        RECT 2219.660 1677.830 2221.180 1677.970 ;
        RECT 2221.040 1594.250 2221.180 1677.830 ;
        RECT 2220.520 1593.930 2220.780 1594.250 ;
        RECT 2220.980 1593.930 2221.240 1594.250 ;
        RECT 2220.580 1559.910 2220.720 1593.930 ;
        RECT 2220.520 1559.590 2220.780 1559.910 ;
        RECT 2220.980 1559.590 2221.240 1559.910 ;
        RECT 2221.040 1511.290 2221.180 1559.590 ;
        RECT 2220.060 1510.970 2220.320 1511.290 ;
        RECT 2220.980 1510.970 2221.240 1511.290 ;
        RECT 2220.120 1510.690 2220.260 1510.970 ;
        RECT 2220.120 1510.550 2220.720 1510.690 ;
        RECT 2220.580 1463.090 2220.720 1510.550 ;
        RECT 2220.580 1462.950 2221.180 1463.090 ;
        RECT 2221.040 1414.730 2221.180 1462.950 ;
        RECT 2220.060 1414.410 2220.320 1414.730 ;
        RECT 2220.980 1414.410 2221.240 1414.730 ;
        RECT 2220.120 1414.130 2220.260 1414.410 ;
        RECT 2220.120 1413.990 2220.720 1414.130 ;
        RECT 2220.580 1366.530 2220.720 1413.990 ;
        RECT 2220.580 1366.390 2221.180 1366.530 ;
        RECT 2221.040 1318.170 2221.180 1366.390 ;
        RECT 2220.060 1317.850 2220.320 1318.170 ;
        RECT 2220.980 1317.850 2221.240 1318.170 ;
        RECT 2220.120 1317.570 2220.260 1317.850 ;
        RECT 2220.120 1317.430 2220.720 1317.570 ;
        RECT 2220.580 1269.970 2220.720 1317.430 ;
        RECT 2220.580 1269.830 2221.180 1269.970 ;
        RECT 2221.040 1221.610 2221.180 1269.830 ;
        RECT 2220.060 1221.290 2220.320 1221.610 ;
        RECT 2220.980 1221.290 2221.240 1221.610 ;
        RECT 2220.120 1221.010 2220.260 1221.290 ;
        RECT 2220.120 1220.870 2220.720 1221.010 ;
        RECT 2220.580 1173.410 2220.720 1220.870 ;
        RECT 2220.580 1173.270 2221.180 1173.410 ;
        RECT 2221.040 1125.050 2221.180 1173.270 ;
        RECT 2220.060 1124.730 2220.320 1125.050 ;
        RECT 2220.980 1124.730 2221.240 1125.050 ;
        RECT 2220.120 1124.450 2220.260 1124.730 ;
        RECT 2220.120 1124.310 2220.720 1124.450 ;
        RECT 2220.580 1076.850 2220.720 1124.310 ;
        RECT 2220.580 1076.710 2221.180 1076.850 ;
        RECT 2221.040 1028.490 2221.180 1076.710 ;
        RECT 2220.060 1028.170 2220.320 1028.490 ;
        RECT 2220.980 1028.170 2221.240 1028.490 ;
        RECT 2220.120 1027.890 2220.260 1028.170 ;
        RECT 2220.120 1027.750 2220.720 1027.890 ;
        RECT 2220.580 980.290 2220.720 1027.750 ;
        RECT 2220.580 980.150 2221.180 980.290 ;
        RECT 2221.040 931.930 2221.180 980.150 ;
        RECT 2220.060 931.610 2220.320 931.930 ;
        RECT 2220.980 931.610 2221.240 931.930 ;
        RECT 2220.120 931.330 2220.260 931.610 ;
        RECT 2220.120 931.190 2220.720 931.330 ;
        RECT 2220.580 917.845 2220.720 931.190 ;
        RECT 2219.590 917.475 2219.870 917.845 ;
        RECT 2220.510 917.475 2220.790 917.845 ;
        RECT 2219.660 869.710 2219.800 917.475 ;
        RECT 2219.600 869.390 2219.860 869.710 ;
        RECT 2220.520 869.390 2220.780 869.710 ;
        RECT 2220.580 835.450 2220.720 869.390 ;
        RECT 2220.120 835.310 2220.720 835.450 ;
        RECT 2220.120 834.770 2220.260 835.310 ;
        RECT 2220.120 834.630 2220.720 834.770 ;
        RECT 2220.580 821.090 2220.720 834.630 ;
        RECT 2220.520 820.770 2220.780 821.090 ;
        RECT 2220.520 786.430 2220.780 786.750 ;
        RECT 2220.580 772.890 2220.720 786.430 ;
        RECT 2220.580 772.810 2221.180 772.890 ;
        RECT 2220.580 772.750 2221.240 772.810 ;
        RECT 2220.980 772.490 2221.240 772.750 ;
        RECT 2221.040 772.335 2221.180 772.490 ;
        RECT 2220.520 724.890 2220.780 725.210 ;
        RECT 2220.580 717.730 2220.720 724.890 ;
        RECT 2220.520 717.410 2220.780 717.730 ;
        RECT 2220.520 641.250 2220.780 641.570 ;
        RECT 2220.580 627.970 2220.720 641.250 ;
        RECT 2220.520 627.650 2220.780 627.970 ;
        RECT 2220.980 592.970 2221.240 593.290 ;
        RECT 2221.040 545.350 2221.180 592.970 ;
        RECT 2220.060 545.090 2220.320 545.350 ;
        RECT 2220.060 545.030 2220.720 545.090 ;
        RECT 2220.980 545.030 2221.240 545.350 ;
        RECT 2220.120 544.950 2220.720 545.030 ;
        RECT 2220.580 531.410 2220.720 544.950 ;
        RECT 2220.520 531.090 2220.780 531.410 ;
        RECT 2220.520 496.410 2220.780 496.730 ;
        RECT 2220.580 483.210 2220.720 496.410 ;
        RECT 2220.580 483.070 2221.180 483.210 ;
        RECT 2221.040 448.790 2221.180 483.070 ;
        RECT 2220.060 448.530 2220.320 448.790 ;
        RECT 2220.060 448.470 2220.720 448.530 ;
        RECT 2220.980 448.470 2221.240 448.790 ;
        RECT 2220.120 448.390 2220.720 448.470 ;
        RECT 2220.580 434.850 2220.720 448.390 ;
        RECT 2220.520 434.530 2220.780 434.850 ;
        RECT 2220.980 386.250 2221.240 386.570 ;
        RECT 2221.040 338.290 2221.180 386.250 ;
        RECT 2220.520 337.970 2220.780 338.290 ;
        RECT 2220.980 337.970 2221.240 338.290 ;
        RECT 2220.580 304.290 2220.720 337.970 ;
        RECT 2220.520 303.970 2220.780 304.290 ;
        RECT 2220.060 303.290 2220.320 303.610 ;
        RECT 2220.120 255.330 2220.260 303.290 ;
        RECT 2220.060 255.010 2220.320 255.330 ;
        RECT 2220.980 255.010 2221.240 255.330 ;
        RECT 2221.040 241.390 2221.180 255.010 ;
        RECT 2220.980 241.070 2221.240 241.390 ;
        RECT 2220.520 193.130 2220.780 193.450 ;
        RECT 2220.580 159.450 2220.720 193.130 ;
        RECT 2220.520 159.130 2220.780 159.450 ;
        RECT 2220.520 144.850 2220.780 145.170 ;
        RECT 2220.580 110.570 2220.720 144.850 ;
        RECT 2220.580 110.430 2221.180 110.570 ;
        RECT 2221.040 62.290 2221.180 110.430 ;
        RECT 2220.120 62.150 2221.180 62.290 ;
        RECT 2220.120 46.230 2220.260 62.150 ;
        RECT 2220.060 45.910 2220.320 46.230 ;
        RECT 2833.700 45.910 2833.960 46.230 ;
        RECT 2833.760 2.400 2833.900 45.910 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
      LAYER via2 ;
        RECT 2219.590 917.520 2219.870 917.800 ;
        RECT 2220.510 917.520 2220.790 917.800 ;
      LAYER met3 ;
        RECT 2219.565 917.810 2219.895 917.825 ;
        RECT 2220.485 917.810 2220.815 917.825 ;
        RECT 2219.565 917.510 2220.815 917.810 ;
        RECT 2219.565 917.495 2219.895 917.510 ;
        RECT 2220.485 917.495 2220.815 917.510 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2227.390 45.800 2227.710 45.860 ;
        RECT 2851.150 45.800 2851.470 45.860 ;
        RECT 2227.390 45.660 2851.470 45.800 ;
        RECT 2227.390 45.600 2227.710 45.660 ;
        RECT 2851.150 45.600 2851.470 45.660 ;
      LAYER via ;
        RECT 2227.420 45.600 2227.680 45.860 ;
        RECT 2851.180 45.600 2851.440 45.860 ;
      LAYER met2 ;
        RECT 2225.045 1700.410 2225.325 1704.000 ;
        RECT 2225.045 1700.270 2226.700 1700.410 ;
        RECT 2225.045 1700.000 2225.325 1700.270 ;
        RECT 2226.560 1659.610 2226.700 1700.270 ;
        RECT 2226.560 1659.470 2227.620 1659.610 ;
        RECT 2227.480 45.890 2227.620 1659.470 ;
        RECT 2227.420 45.570 2227.680 45.890 ;
        RECT 2851.180 45.570 2851.440 45.890 ;
        RECT 2851.240 2.400 2851.380 45.570 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2234.750 45.460 2235.070 45.520 ;
        RECT 2869.090 45.460 2869.410 45.520 ;
        RECT 2234.750 45.320 2869.410 45.460 ;
        RECT 2234.750 45.260 2235.070 45.320 ;
        RECT 2869.090 45.260 2869.410 45.320 ;
      LAYER via ;
        RECT 2234.780 45.260 2235.040 45.520 ;
        RECT 2869.120 45.260 2869.380 45.520 ;
      LAYER met2 ;
        RECT 2231.485 1700.410 2231.765 1704.000 ;
        RECT 2231.485 1700.270 2233.140 1700.410 ;
        RECT 2231.485 1700.000 2231.765 1700.270 ;
        RECT 2233.000 1677.970 2233.140 1700.270 ;
        RECT 2233.000 1677.830 2234.980 1677.970 ;
        RECT 2234.840 45.550 2234.980 1677.830 ;
        RECT 2234.780 45.230 2235.040 45.550 ;
        RECT 2869.120 45.230 2869.380 45.550 ;
        RECT 2869.180 2.400 2869.320 45.230 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2241.650 45.120 2241.970 45.180 ;
        RECT 2887.030 45.120 2887.350 45.180 ;
        RECT 2241.650 44.980 2887.350 45.120 ;
        RECT 2241.650 44.920 2241.970 44.980 ;
        RECT 2887.030 44.920 2887.350 44.980 ;
      LAYER via ;
        RECT 2241.680 44.920 2241.940 45.180 ;
        RECT 2887.060 44.920 2887.320 45.180 ;
      LAYER met2 ;
        RECT 2238.385 1701.090 2238.665 1704.000 ;
        RECT 2238.385 1700.950 2240.500 1701.090 ;
        RECT 2238.385 1700.000 2238.665 1700.950 ;
        RECT 2240.360 1688.340 2240.500 1700.950 ;
        RECT 2240.360 1688.200 2241.880 1688.340 ;
        RECT 2241.740 45.210 2241.880 1688.200 ;
        RECT 2241.680 44.890 2241.940 45.210 ;
        RECT 2887.060 44.890 2887.320 45.210 ;
        RECT 2887.120 2.400 2887.260 44.890 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2248.550 44.780 2248.870 44.840 ;
        RECT 2904.970 44.780 2905.290 44.840 ;
        RECT 2248.550 44.640 2905.290 44.780 ;
        RECT 2248.550 44.580 2248.870 44.640 ;
        RECT 2904.970 44.580 2905.290 44.640 ;
      LAYER via ;
        RECT 2248.580 44.580 2248.840 44.840 ;
        RECT 2905.000 44.580 2905.260 44.840 ;
      LAYER met2 ;
        RECT 2245.285 1700.410 2245.565 1704.000 ;
        RECT 2245.285 1700.270 2246.940 1700.410 ;
        RECT 2245.285 1700.000 2245.565 1700.270 ;
        RECT 2246.800 1686.130 2246.940 1700.270 ;
        RECT 2246.800 1685.990 2248.780 1686.130 ;
        RECT 2248.640 44.870 2248.780 1685.990 ;
        RECT 2248.580 44.550 2248.840 44.870 ;
        RECT 2905.000 44.550 2905.260 44.870 ;
        RECT 2905.060 2.400 2905.200 44.550 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 852.910 33.900 853.230 33.960 ;
        RECT 1469.770 33.900 1470.090 33.960 ;
        RECT 852.910 33.760 1470.090 33.900 ;
        RECT 852.910 33.700 853.230 33.760 ;
        RECT 1469.770 33.700 1470.090 33.760 ;
      LAYER via ;
        RECT 852.940 33.700 853.200 33.960 ;
        RECT 1469.800 33.700 1470.060 33.960 ;
      LAYER met2 ;
        RECT 1470.645 1700.410 1470.925 1704.000 ;
        RECT 1469.860 1700.270 1470.925 1700.410 ;
        RECT 1469.860 33.990 1470.000 1700.270 ;
        RECT 1470.645 1700.000 1470.925 1700.270 ;
        RECT 852.940 33.670 853.200 33.990 ;
        RECT 1469.800 33.670 1470.060 33.990 ;
        RECT 853.000 2.400 853.140 33.670 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 34.240 871.170 34.300 ;
        RECT 1476.670 34.240 1476.990 34.300 ;
        RECT 870.850 34.100 1476.990 34.240 ;
        RECT 870.850 34.040 871.170 34.100 ;
        RECT 1476.670 34.040 1476.990 34.100 ;
      LAYER via ;
        RECT 870.880 34.040 871.140 34.300 ;
        RECT 1476.700 34.040 1476.960 34.300 ;
      LAYER met2 ;
        RECT 1477.545 1700.410 1477.825 1704.000 ;
        RECT 1476.760 1700.270 1477.825 1700.410 ;
        RECT 1476.760 34.330 1476.900 1700.270 ;
        RECT 1477.545 1700.000 1477.825 1700.270 ;
        RECT 870.880 34.010 871.140 34.330 ;
        RECT 1476.700 34.010 1476.960 34.330 ;
        RECT 870.940 2.400 871.080 34.010 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 888.790 30.500 889.110 30.560 ;
        RECT 1483.570 30.500 1483.890 30.560 ;
        RECT 888.790 30.360 1483.890 30.500 ;
        RECT 888.790 30.300 889.110 30.360 ;
        RECT 1483.570 30.300 1483.890 30.360 ;
      LAYER via ;
        RECT 888.820 30.300 889.080 30.560 ;
        RECT 1483.600 30.300 1483.860 30.560 ;
      LAYER met2 ;
        RECT 1484.445 1700.410 1484.725 1704.000 ;
        RECT 1483.660 1700.270 1484.725 1700.410 ;
        RECT 1483.660 30.590 1483.800 1700.270 ;
        RECT 1484.445 1700.000 1484.725 1700.270 ;
        RECT 888.820 30.270 889.080 30.590 ;
        RECT 1483.600 30.270 1483.860 30.590 ;
        RECT 888.880 2.400 889.020 30.270 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 906.730 30.160 907.050 30.220 ;
        RECT 1490.470 30.160 1490.790 30.220 ;
        RECT 906.730 30.020 1490.790 30.160 ;
        RECT 906.730 29.960 907.050 30.020 ;
        RECT 1490.470 29.960 1490.790 30.020 ;
      LAYER via ;
        RECT 906.760 29.960 907.020 30.220 ;
        RECT 1490.500 29.960 1490.760 30.220 ;
      LAYER met2 ;
        RECT 1490.885 1700.410 1491.165 1704.000 ;
        RECT 1490.560 1700.270 1491.165 1700.410 ;
        RECT 1490.560 30.250 1490.700 1700.270 ;
        RECT 1490.885 1700.000 1491.165 1700.270 ;
        RECT 906.760 29.930 907.020 30.250 ;
        RECT 1490.500 29.930 1490.760 30.250 ;
        RECT 906.820 2.400 906.960 29.930 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 29.820 924.530 29.880 ;
        RECT 1497.370 29.820 1497.690 29.880 ;
        RECT 924.210 29.680 1497.690 29.820 ;
        RECT 924.210 29.620 924.530 29.680 ;
        RECT 1497.370 29.620 1497.690 29.680 ;
      LAYER via ;
        RECT 924.240 29.620 924.500 29.880 ;
        RECT 1497.400 29.620 1497.660 29.880 ;
      LAYER met2 ;
        RECT 1497.785 1700.410 1498.065 1704.000 ;
        RECT 1497.460 1700.270 1498.065 1700.410 ;
        RECT 1497.460 29.910 1497.600 1700.270 ;
        RECT 1497.785 1700.000 1498.065 1700.270 ;
        RECT 924.240 29.590 924.500 29.910 ;
        RECT 1497.400 29.590 1497.660 29.910 ;
        RECT 924.300 2.400 924.440 29.590 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 942.150 29.480 942.470 29.540 ;
        RECT 1504.270 29.480 1504.590 29.540 ;
        RECT 942.150 29.340 1504.590 29.480 ;
        RECT 942.150 29.280 942.470 29.340 ;
        RECT 1504.270 29.280 1504.590 29.340 ;
      LAYER via ;
        RECT 942.180 29.280 942.440 29.540 ;
        RECT 1504.300 29.280 1504.560 29.540 ;
      LAYER met2 ;
        RECT 1504.225 1700.000 1504.505 1704.000 ;
        RECT 1504.360 29.570 1504.500 1700.000 ;
        RECT 942.180 29.250 942.440 29.570 ;
        RECT 1504.300 29.250 1504.560 29.570 ;
        RECT 942.240 2.400 942.380 29.250 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 29.140 960.410 29.200 ;
        RECT 1511.170 29.140 1511.490 29.200 ;
        RECT 960.090 29.000 1511.490 29.140 ;
        RECT 960.090 28.940 960.410 29.000 ;
        RECT 1511.170 28.940 1511.490 29.000 ;
      LAYER via ;
        RECT 960.120 28.940 960.380 29.200 ;
        RECT 1511.200 28.940 1511.460 29.200 ;
      LAYER met2 ;
        RECT 1511.125 1700.000 1511.405 1704.000 ;
        RECT 1511.260 29.230 1511.400 1700.000 ;
        RECT 960.120 28.910 960.380 29.230 ;
        RECT 1511.200 28.910 1511.460 29.230 ;
        RECT 960.180 2.400 960.320 28.910 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.030 28.800 978.350 28.860 ;
        RECT 1518.070 28.800 1518.390 28.860 ;
        RECT 978.030 28.660 1518.390 28.800 ;
        RECT 978.030 28.600 978.350 28.660 ;
        RECT 1518.070 28.600 1518.390 28.660 ;
      LAYER via ;
        RECT 978.060 28.600 978.320 28.860 ;
        RECT 1518.100 28.600 1518.360 28.860 ;
      LAYER met2 ;
        RECT 1518.025 1700.000 1518.305 1704.000 ;
        RECT 1518.160 28.890 1518.300 1700.000 ;
        RECT 978.060 28.570 978.320 28.890 ;
        RECT 1518.100 28.570 1518.360 28.890 ;
        RECT 978.120 2.400 978.260 28.570 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 32.880 657.270 32.940 ;
        RECT 1395.250 32.880 1395.570 32.940 ;
        RECT 656.950 32.740 1395.570 32.880 ;
        RECT 656.950 32.680 657.270 32.740 ;
        RECT 1395.250 32.680 1395.570 32.740 ;
      LAYER via ;
        RECT 656.980 32.680 657.240 32.940 ;
        RECT 1395.280 32.680 1395.540 32.940 ;
      LAYER met2 ;
        RECT 1396.585 1700.410 1396.865 1704.000 ;
        RECT 1395.340 1700.270 1396.865 1700.410 ;
        RECT 1395.340 32.970 1395.480 1700.270 ;
        RECT 1396.585 1700.000 1396.865 1700.270 ;
        RECT 656.980 32.650 657.240 32.970 ;
        RECT 1395.280 32.650 1395.540 32.970 ;
        RECT 657.040 2.400 657.180 32.650 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1518.530 1678.480 1518.850 1678.540 ;
        RECT 1523.130 1678.480 1523.450 1678.540 ;
        RECT 1518.530 1678.340 1523.450 1678.480 ;
        RECT 1518.530 1678.280 1518.850 1678.340 ;
        RECT 1523.130 1678.280 1523.450 1678.340 ;
        RECT 995.970 28.460 996.290 28.520 ;
        RECT 1518.530 28.460 1518.850 28.520 ;
        RECT 995.970 28.320 1518.850 28.460 ;
        RECT 995.970 28.260 996.290 28.320 ;
        RECT 1518.530 28.260 1518.850 28.320 ;
      LAYER via ;
        RECT 1518.560 1678.280 1518.820 1678.540 ;
        RECT 1523.160 1678.280 1523.420 1678.540 ;
        RECT 996.000 28.260 996.260 28.520 ;
        RECT 1518.560 28.260 1518.820 28.520 ;
      LAYER met2 ;
        RECT 1524.465 1700.410 1524.745 1704.000 ;
        RECT 1523.220 1700.270 1524.745 1700.410 ;
        RECT 1523.220 1678.570 1523.360 1700.270 ;
        RECT 1524.465 1700.000 1524.745 1700.270 ;
        RECT 1518.560 1678.250 1518.820 1678.570 ;
        RECT 1523.160 1678.250 1523.420 1678.570 ;
        RECT 1518.620 28.550 1518.760 1678.250 ;
        RECT 996.000 28.230 996.260 28.550 ;
        RECT 1518.560 28.230 1518.820 28.550 ;
        RECT 996.060 2.400 996.200 28.230 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1527.345 1490.645 1527.515 1538.755 ;
        RECT 1525.965 1207.425 1526.135 1255.875 ;
        RECT 1526.425 1014.305 1526.595 1028.415 ;
        RECT 1526.425 979.625 1526.595 1007.335 ;
        RECT 1526.425 766.105 1526.595 814.215 ;
        RECT 1526.425 710.685 1526.595 765.595 ;
        RECT 1526.885 614.125 1527.055 662.235 ;
        RECT 1526.425 510.765 1526.595 531.335 ;
        RECT 1526.425 324.445 1526.595 372.215 ;
        RECT 1526.885 124.185 1527.055 179.435 ;
      LAYER mcon ;
        RECT 1527.345 1538.585 1527.515 1538.755 ;
        RECT 1525.965 1255.705 1526.135 1255.875 ;
        RECT 1526.425 1028.245 1526.595 1028.415 ;
        RECT 1526.425 1007.165 1526.595 1007.335 ;
        RECT 1526.425 814.045 1526.595 814.215 ;
        RECT 1526.425 765.425 1526.595 765.595 ;
        RECT 1526.885 662.065 1527.055 662.235 ;
        RECT 1526.425 531.165 1526.595 531.335 ;
        RECT 1526.425 372.045 1526.595 372.215 ;
        RECT 1526.885 179.265 1527.055 179.435 ;
      LAYER met1 ;
        RECT 1526.810 1642.440 1527.130 1642.500 ;
        RECT 1530.490 1642.440 1530.810 1642.500 ;
        RECT 1526.810 1642.300 1530.810 1642.440 ;
        RECT 1526.810 1642.240 1527.130 1642.300 ;
        RECT 1530.490 1642.240 1530.810 1642.300 ;
        RECT 1526.810 1563.900 1527.130 1563.960 ;
        RECT 1528.190 1563.900 1528.510 1563.960 ;
        RECT 1526.810 1563.760 1528.510 1563.900 ;
        RECT 1526.810 1563.700 1527.130 1563.760 ;
        RECT 1528.190 1563.700 1528.510 1563.760 ;
        RECT 1527.285 1538.740 1527.575 1538.785 ;
        RECT 1527.730 1538.740 1528.050 1538.800 ;
        RECT 1527.285 1538.600 1528.050 1538.740 ;
        RECT 1527.285 1538.555 1527.575 1538.600 ;
        RECT 1527.730 1538.540 1528.050 1538.600 ;
        RECT 1527.270 1490.800 1527.590 1490.860 ;
        RECT 1527.075 1490.660 1527.590 1490.800 ;
        RECT 1527.270 1490.600 1527.590 1490.660 ;
        RECT 1527.270 1449.120 1527.590 1449.380 ;
        RECT 1527.360 1448.700 1527.500 1449.120 ;
        RECT 1527.270 1448.440 1527.590 1448.700 ;
        RECT 1527.270 1400.700 1527.590 1400.760 ;
        RECT 1526.440 1400.560 1527.590 1400.700 ;
        RECT 1526.440 1400.420 1526.580 1400.560 ;
        RECT 1527.270 1400.500 1527.590 1400.560 ;
        RECT 1526.350 1400.160 1526.670 1400.420 ;
        RECT 1525.905 1255.860 1526.195 1255.905 ;
        RECT 1526.350 1255.860 1526.670 1255.920 ;
        RECT 1525.905 1255.720 1526.670 1255.860 ;
        RECT 1525.905 1255.675 1526.195 1255.720 ;
        RECT 1526.350 1255.660 1526.670 1255.720 ;
        RECT 1525.890 1207.580 1526.210 1207.640 ;
        RECT 1525.695 1207.440 1526.210 1207.580 ;
        RECT 1525.890 1207.380 1526.210 1207.440 ;
        RECT 1525.890 1159.300 1526.210 1159.360 ;
        RECT 1526.350 1159.300 1526.670 1159.360 ;
        RECT 1525.890 1159.160 1526.670 1159.300 ;
        RECT 1525.890 1159.100 1526.210 1159.160 ;
        RECT 1526.350 1159.100 1526.670 1159.160 ;
        RECT 1526.810 1076.680 1527.130 1076.740 ;
        RECT 1526.440 1076.540 1527.130 1076.680 ;
        RECT 1526.440 1076.400 1526.580 1076.540 ;
        RECT 1526.810 1076.480 1527.130 1076.540 ;
        RECT 1526.350 1076.140 1526.670 1076.400 ;
        RECT 1526.350 1028.400 1526.670 1028.460 ;
        RECT 1526.155 1028.260 1526.670 1028.400 ;
        RECT 1526.350 1028.200 1526.670 1028.260 ;
        RECT 1526.350 1014.460 1526.670 1014.520 ;
        RECT 1526.155 1014.320 1526.670 1014.460 ;
        RECT 1526.350 1014.260 1526.670 1014.320 ;
        RECT 1526.350 1007.320 1526.670 1007.380 ;
        RECT 1526.155 1007.180 1526.670 1007.320 ;
        RECT 1526.350 1007.120 1526.670 1007.180 ;
        RECT 1526.350 979.780 1526.670 979.840 ;
        RECT 1526.155 979.640 1526.670 979.780 ;
        RECT 1526.350 979.580 1526.670 979.640 ;
        RECT 1525.890 917.900 1526.210 917.960 ;
        RECT 1527.270 917.900 1527.590 917.960 ;
        RECT 1525.890 917.760 1527.590 917.900 ;
        RECT 1525.890 917.700 1526.210 917.760 ;
        RECT 1527.270 917.700 1527.590 917.760 ;
        RECT 1526.810 869.620 1527.130 869.680 ;
        RECT 1527.270 869.620 1527.590 869.680 ;
        RECT 1526.810 869.480 1527.590 869.620 ;
        RECT 1526.810 869.420 1527.130 869.480 ;
        RECT 1527.270 869.420 1527.590 869.480 ;
        RECT 1526.365 814.200 1526.655 814.245 ;
        RECT 1526.810 814.200 1527.130 814.260 ;
        RECT 1526.365 814.060 1527.130 814.200 ;
        RECT 1526.365 814.015 1526.655 814.060 ;
        RECT 1526.810 814.000 1527.130 814.060 ;
        RECT 1526.350 766.260 1526.670 766.320 ;
        RECT 1526.155 766.120 1526.670 766.260 ;
        RECT 1526.350 766.060 1526.670 766.120 ;
        RECT 1526.350 765.580 1526.670 765.640 ;
        RECT 1526.155 765.440 1526.670 765.580 ;
        RECT 1526.350 765.380 1526.670 765.440 ;
        RECT 1526.365 710.840 1526.655 710.885 ;
        RECT 1526.810 710.840 1527.130 710.900 ;
        RECT 1526.365 710.700 1527.130 710.840 ;
        RECT 1526.365 710.655 1526.655 710.700 ;
        RECT 1526.810 710.640 1527.130 710.700 ;
        RECT 1526.810 662.220 1527.130 662.280 ;
        RECT 1526.615 662.080 1527.130 662.220 ;
        RECT 1526.810 662.020 1527.130 662.080 ;
        RECT 1526.810 614.280 1527.130 614.340 ;
        RECT 1526.615 614.140 1527.130 614.280 ;
        RECT 1526.810 614.080 1527.130 614.140 ;
        RECT 1524.970 593.880 1525.290 593.940 ;
        RECT 1526.810 593.880 1527.130 593.940 ;
        RECT 1524.970 593.740 1527.130 593.880 ;
        RECT 1524.970 593.680 1525.290 593.740 ;
        RECT 1526.810 593.680 1527.130 593.740 ;
        RECT 1526.350 531.320 1526.670 531.380 ;
        RECT 1526.155 531.180 1526.670 531.320 ;
        RECT 1526.350 531.120 1526.670 531.180 ;
        RECT 1526.350 510.920 1526.670 510.980 ;
        RECT 1526.155 510.780 1526.670 510.920 ;
        RECT 1526.350 510.720 1526.670 510.780 ;
        RECT 1527.730 435.100 1528.050 435.160 ;
        RECT 1527.360 434.960 1528.050 435.100 ;
        RECT 1527.360 434.820 1527.500 434.960 ;
        RECT 1527.730 434.900 1528.050 434.960 ;
        RECT 1527.270 434.560 1527.590 434.820 ;
        RECT 1526.350 372.880 1526.670 372.940 ;
        RECT 1527.270 372.880 1527.590 372.940 ;
        RECT 1526.350 372.740 1527.590 372.880 ;
        RECT 1526.350 372.680 1526.670 372.740 ;
        RECT 1527.270 372.680 1527.590 372.740 ;
        RECT 1526.350 372.200 1526.670 372.260 ;
        RECT 1526.155 372.060 1526.670 372.200 ;
        RECT 1526.350 372.000 1526.670 372.060 ;
        RECT 1526.365 324.600 1526.655 324.645 ;
        RECT 1526.810 324.600 1527.130 324.660 ;
        RECT 1526.365 324.460 1527.130 324.600 ;
        RECT 1526.365 324.415 1526.655 324.460 ;
        RECT 1526.810 324.400 1527.130 324.460 ;
        RECT 1526.810 179.420 1527.130 179.480 ;
        RECT 1526.615 179.280 1527.130 179.420 ;
        RECT 1526.810 179.220 1527.130 179.280 ;
        RECT 1526.810 124.340 1527.130 124.400 ;
        RECT 1526.615 124.200 1527.130 124.340 ;
        RECT 1526.810 124.140 1527.130 124.200 ;
        RECT 1013.450 28.120 1013.770 28.180 ;
        RECT 1525.890 28.120 1526.210 28.180 ;
        RECT 1013.450 27.980 1526.210 28.120 ;
        RECT 1013.450 27.920 1013.770 27.980 ;
        RECT 1525.890 27.920 1526.210 27.980 ;
      LAYER via ;
        RECT 1526.840 1642.240 1527.100 1642.500 ;
        RECT 1530.520 1642.240 1530.780 1642.500 ;
        RECT 1526.840 1563.700 1527.100 1563.960 ;
        RECT 1528.220 1563.700 1528.480 1563.960 ;
        RECT 1527.760 1538.540 1528.020 1538.800 ;
        RECT 1527.300 1490.600 1527.560 1490.860 ;
        RECT 1527.300 1449.120 1527.560 1449.380 ;
        RECT 1527.300 1448.440 1527.560 1448.700 ;
        RECT 1527.300 1400.500 1527.560 1400.760 ;
        RECT 1526.380 1400.160 1526.640 1400.420 ;
        RECT 1526.380 1255.660 1526.640 1255.920 ;
        RECT 1525.920 1207.380 1526.180 1207.640 ;
        RECT 1525.920 1159.100 1526.180 1159.360 ;
        RECT 1526.380 1159.100 1526.640 1159.360 ;
        RECT 1526.840 1076.480 1527.100 1076.740 ;
        RECT 1526.380 1076.140 1526.640 1076.400 ;
        RECT 1526.380 1028.200 1526.640 1028.460 ;
        RECT 1526.380 1014.260 1526.640 1014.520 ;
        RECT 1526.380 1007.120 1526.640 1007.380 ;
        RECT 1526.380 979.580 1526.640 979.840 ;
        RECT 1525.920 917.700 1526.180 917.960 ;
        RECT 1527.300 917.700 1527.560 917.960 ;
        RECT 1526.840 869.420 1527.100 869.680 ;
        RECT 1527.300 869.420 1527.560 869.680 ;
        RECT 1526.840 814.000 1527.100 814.260 ;
        RECT 1526.380 766.060 1526.640 766.320 ;
        RECT 1526.380 765.380 1526.640 765.640 ;
        RECT 1526.840 710.640 1527.100 710.900 ;
        RECT 1526.840 662.020 1527.100 662.280 ;
        RECT 1526.840 614.080 1527.100 614.340 ;
        RECT 1525.000 593.680 1525.260 593.940 ;
        RECT 1526.840 593.680 1527.100 593.940 ;
        RECT 1526.380 531.120 1526.640 531.380 ;
        RECT 1526.380 510.720 1526.640 510.980 ;
        RECT 1527.760 434.900 1528.020 435.160 ;
        RECT 1527.300 434.560 1527.560 434.820 ;
        RECT 1526.380 372.680 1526.640 372.940 ;
        RECT 1527.300 372.680 1527.560 372.940 ;
        RECT 1526.380 372.000 1526.640 372.260 ;
        RECT 1526.840 324.400 1527.100 324.660 ;
        RECT 1526.840 179.220 1527.100 179.480 ;
        RECT 1526.840 124.140 1527.100 124.400 ;
        RECT 1013.480 27.920 1013.740 28.180 ;
        RECT 1525.920 27.920 1526.180 28.180 ;
      LAYER met2 ;
        RECT 1531.365 1700.410 1531.645 1704.000 ;
        RECT 1530.580 1700.270 1531.645 1700.410 ;
        RECT 1530.580 1642.530 1530.720 1700.270 ;
        RECT 1531.365 1700.000 1531.645 1700.270 ;
        RECT 1526.840 1642.210 1527.100 1642.530 ;
        RECT 1530.520 1642.210 1530.780 1642.530 ;
        RECT 1526.900 1563.990 1527.040 1642.210 ;
        RECT 1526.840 1563.670 1527.100 1563.990 ;
        RECT 1528.220 1563.670 1528.480 1563.990 ;
        RECT 1528.280 1539.250 1528.420 1563.670 ;
        RECT 1527.820 1539.110 1528.420 1539.250 ;
        RECT 1527.820 1538.830 1527.960 1539.110 ;
        RECT 1527.760 1538.510 1528.020 1538.830 ;
        RECT 1527.300 1490.570 1527.560 1490.890 ;
        RECT 1527.360 1449.410 1527.500 1490.570 ;
        RECT 1527.300 1449.090 1527.560 1449.410 ;
        RECT 1527.300 1448.410 1527.560 1448.730 ;
        RECT 1527.360 1400.790 1527.500 1448.410 ;
        RECT 1527.300 1400.470 1527.560 1400.790 ;
        RECT 1526.380 1400.130 1526.640 1400.450 ;
        RECT 1526.440 1393.845 1526.580 1400.130 ;
        RECT 1526.370 1393.475 1526.650 1393.845 ;
        RECT 1527.750 1393.475 1528.030 1393.845 ;
        RECT 1527.820 1268.610 1527.960 1393.475 ;
        RECT 1526.440 1268.470 1527.960 1268.610 ;
        RECT 1526.440 1255.950 1526.580 1268.470 ;
        RECT 1526.380 1255.630 1526.640 1255.950 ;
        RECT 1525.920 1207.350 1526.180 1207.670 ;
        RECT 1525.980 1159.390 1526.120 1207.350 ;
        RECT 1525.920 1159.070 1526.180 1159.390 ;
        RECT 1526.380 1159.070 1526.640 1159.390 ;
        RECT 1526.440 1104.050 1526.580 1159.070 ;
        RECT 1526.440 1103.910 1527.040 1104.050 ;
        RECT 1526.900 1076.770 1527.040 1103.910 ;
        RECT 1526.840 1076.450 1527.100 1076.770 ;
        RECT 1526.380 1076.110 1526.640 1076.430 ;
        RECT 1526.440 1028.490 1526.580 1076.110 ;
        RECT 1526.380 1028.170 1526.640 1028.490 ;
        RECT 1526.380 1014.230 1526.640 1014.550 ;
        RECT 1526.440 1007.410 1526.580 1014.230 ;
        RECT 1526.380 1007.090 1526.640 1007.410 ;
        RECT 1526.380 979.550 1526.640 979.870 ;
        RECT 1526.440 942.210 1526.580 979.550 ;
        RECT 1525.980 942.070 1526.580 942.210 ;
        RECT 1525.980 917.990 1526.120 942.070 ;
        RECT 1525.920 917.670 1526.180 917.990 ;
        RECT 1527.300 917.670 1527.560 917.990 ;
        RECT 1527.360 869.710 1527.500 917.670 ;
        RECT 1526.840 869.390 1527.100 869.710 ;
        RECT 1527.300 869.390 1527.560 869.710 ;
        RECT 1526.900 814.290 1527.040 869.390 ;
        RECT 1526.840 813.970 1527.100 814.290 ;
        RECT 1526.380 766.030 1526.640 766.350 ;
        RECT 1526.440 765.670 1526.580 766.030 ;
        RECT 1526.380 765.350 1526.640 765.670 ;
        RECT 1526.840 710.610 1527.100 710.930 ;
        RECT 1526.900 662.310 1527.040 710.610 ;
        RECT 1526.840 661.990 1527.100 662.310 ;
        RECT 1526.840 614.050 1527.100 614.370 ;
        RECT 1526.900 593.970 1527.040 614.050 ;
        RECT 1525.000 593.650 1525.260 593.970 ;
        RECT 1526.840 593.650 1527.100 593.970 ;
        RECT 1525.060 566.285 1525.200 593.650 ;
        RECT 1524.990 565.915 1525.270 566.285 ;
        RECT 1526.370 565.915 1526.650 566.285 ;
        RECT 1526.440 531.410 1526.580 565.915 ;
        RECT 1526.380 531.090 1526.640 531.410 ;
        RECT 1526.380 510.690 1526.640 511.010 ;
        RECT 1526.440 486.610 1526.580 510.690 ;
        RECT 1526.440 486.470 1527.960 486.610 ;
        RECT 1527.820 435.190 1527.960 486.470 ;
        RECT 1527.760 434.870 1528.020 435.190 ;
        RECT 1527.300 434.530 1527.560 434.850 ;
        RECT 1527.360 372.970 1527.500 434.530 ;
        RECT 1526.380 372.650 1526.640 372.970 ;
        RECT 1527.300 372.650 1527.560 372.970 ;
        RECT 1526.440 372.290 1526.580 372.650 ;
        RECT 1526.380 371.970 1526.640 372.290 ;
        RECT 1526.840 324.370 1527.100 324.690 ;
        RECT 1526.900 265.610 1527.040 324.370 ;
        RECT 1526.900 265.470 1527.500 265.610 ;
        RECT 1527.360 203.730 1527.500 265.470 ;
        RECT 1526.900 203.590 1527.500 203.730 ;
        RECT 1526.900 179.510 1527.040 203.590 ;
        RECT 1526.840 179.190 1527.100 179.510 ;
        RECT 1526.840 124.110 1527.100 124.430 ;
        RECT 1526.900 76.005 1527.040 124.110 ;
        RECT 1525.910 75.635 1526.190 76.005 ;
        RECT 1526.830 75.635 1527.110 76.005 ;
        RECT 1525.980 28.210 1526.120 75.635 ;
        RECT 1013.480 27.890 1013.740 28.210 ;
        RECT 1525.920 27.890 1526.180 28.210 ;
        RECT 1013.540 2.400 1013.680 27.890 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
      LAYER via2 ;
        RECT 1526.370 1393.520 1526.650 1393.800 ;
        RECT 1527.750 1393.520 1528.030 1393.800 ;
        RECT 1524.990 565.960 1525.270 566.240 ;
        RECT 1526.370 565.960 1526.650 566.240 ;
        RECT 1525.910 75.680 1526.190 75.960 ;
        RECT 1526.830 75.680 1527.110 75.960 ;
      LAYER met3 ;
        RECT 1526.345 1393.810 1526.675 1393.825 ;
        RECT 1527.725 1393.810 1528.055 1393.825 ;
        RECT 1526.345 1393.510 1528.055 1393.810 ;
        RECT 1526.345 1393.495 1526.675 1393.510 ;
        RECT 1527.725 1393.495 1528.055 1393.510 ;
        RECT 1524.965 566.250 1525.295 566.265 ;
        RECT 1526.345 566.250 1526.675 566.265 ;
        RECT 1524.965 565.950 1526.675 566.250 ;
        RECT 1524.965 565.935 1525.295 565.950 ;
        RECT 1526.345 565.935 1526.675 565.950 ;
        RECT 1525.885 75.970 1526.215 75.985 ;
        RECT 1526.805 75.970 1527.135 75.985 ;
        RECT 1525.885 75.670 1527.135 75.970 ;
        RECT 1525.885 75.655 1526.215 75.670 ;
        RECT 1526.805 75.655 1527.135 75.670 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1532.330 1678.480 1532.650 1678.540 ;
        RECT 1536.470 1678.480 1536.790 1678.540 ;
        RECT 1532.330 1678.340 1536.790 1678.480 ;
        RECT 1532.330 1678.280 1532.650 1678.340 ;
        RECT 1536.470 1678.280 1536.790 1678.340 ;
        RECT 1031.390 27.780 1031.710 27.840 ;
        RECT 1532.330 27.780 1532.650 27.840 ;
        RECT 1031.390 27.640 1532.650 27.780 ;
        RECT 1031.390 27.580 1031.710 27.640 ;
        RECT 1532.330 27.580 1532.650 27.640 ;
      LAYER via ;
        RECT 1532.360 1678.280 1532.620 1678.540 ;
        RECT 1536.500 1678.280 1536.760 1678.540 ;
        RECT 1031.420 27.580 1031.680 27.840 ;
        RECT 1532.360 27.580 1532.620 27.840 ;
      LAYER met2 ;
        RECT 1538.265 1700.410 1538.545 1704.000 ;
        RECT 1536.560 1700.270 1538.545 1700.410 ;
        RECT 1536.560 1678.570 1536.700 1700.270 ;
        RECT 1538.265 1700.000 1538.545 1700.270 ;
        RECT 1532.360 1678.250 1532.620 1678.570 ;
        RECT 1536.500 1678.250 1536.760 1678.570 ;
        RECT 1532.420 27.870 1532.560 1678.250 ;
        RECT 1031.420 27.550 1031.680 27.870 ;
        RECT 1532.360 27.550 1532.620 27.870 ;
        RECT 1031.480 2.400 1031.620 27.550 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1539.765 1290.385 1539.935 1352.435 ;
        RECT 1539.765 1221.025 1539.935 1255.875 ;
        RECT 1540.225 1062.585 1540.395 1087.235 ;
        RECT 1540.225 966.025 1540.395 980.135 ;
        RECT 1540.225 758.965 1540.395 807.075 ;
        RECT 1539.765 372.725 1539.935 420.835 ;
        RECT 1540.225 324.445 1540.395 331.415 ;
        RECT 1540.685 64.685 1540.855 97.495 ;
      LAYER mcon ;
        RECT 1539.765 1352.265 1539.935 1352.435 ;
        RECT 1539.765 1255.705 1539.935 1255.875 ;
        RECT 1540.225 1087.065 1540.395 1087.235 ;
        RECT 1540.225 979.965 1540.395 980.135 ;
        RECT 1540.225 806.905 1540.395 807.075 ;
        RECT 1539.765 420.665 1539.935 420.835 ;
        RECT 1540.225 331.245 1540.395 331.415 ;
        RECT 1540.685 97.325 1540.855 97.495 ;
      LAYER met1 ;
        RECT 1540.610 1642.440 1540.930 1642.500 ;
        RECT 1543.370 1642.440 1543.690 1642.500 ;
        RECT 1540.610 1642.300 1543.690 1642.440 ;
        RECT 1540.610 1642.240 1540.930 1642.300 ;
        RECT 1543.370 1642.240 1543.690 1642.300 ;
        RECT 1540.150 1545.540 1540.470 1545.600 ;
        RECT 1541.070 1545.540 1541.390 1545.600 ;
        RECT 1540.150 1545.400 1541.390 1545.540 ;
        RECT 1540.150 1545.340 1540.470 1545.400 ;
        RECT 1541.070 1545.340 1541.390 1545.400 ;
        RECT 1540.610 1490.460 1540.930 1490.520 ;
        RECT 1541.070 1490.460 1541.390 1490.520 ;
        RECT 1540.610 1490.320 1541.390 1490.460 ;
        RECT 1540.610 1490.260 1540.930 1490.320 ;
        RECT 1541.070 1490.260 1541.390 1490.320 ;
        RECT 1539.690 1393.900 1540.010 1393.960 ;
        RECT 1541.070 1393.900 1541.390 1393.960 ;
        RECT 1539.690 1393.760 1541.390 1393.900 ;
        RECT 1539.690 1393.700 1540.010 1393.760 ;
        RECT 1541.070 1393.700 1541.390 1393.760 ;
        RECT 1539.690 1352.420 1540.010 1352.480 ;
        RECT 1539.495 1352.280 1540.010 1352.420 ;
        RECT 1539.690 1352.220 1540.010 1352.280 ;
        RECT 1539.690 1290.540 1540.010 1290.600 ;
        RECT 1539.495 1290.400 1540.010 1290.540 ;
        RECT 1539.690 1290.340 1540.010 1290.400 ;
        RECT 1539.690 1255.860 1540.010 1255.920 ;
        RECT 1539.495 1255.720 1540.010 1255.860 ;
        RECT 1539.690 1255.660 1540.010 1255.720 ;
        RECT 1539.705 1221.180 1539.995 1221.225 ;
        RECT 1540.150 1221.180 1540.470 1221.240 ;
        RECT 1539.705 1221.040 1540.470 1221.180 ;
        RECT 1539.705 1220.995 1539.995 1221.040 ;
        RECT 1540.150 1220.980 1540.470 1221.040 ;
        RECT 1540.150 1159.780 1540.470 1160.040 ;
        RECT 1540.240 1159.360 1540.380 1159.780 ;
        RECT 1540.150 1159.100 1540.470 1159.360 ;
        RECT 1540.150 1087.220 1540.470 1087.280 ;
        RECT 1539.955 1087.080 1540.470 1087.220 ;
        RECT 1540.150 1087.020 1540.470 1087.080 ;
        RECT 1540.150 1062.740 1540.470 1062.800 ;
        RECT 1539.955 1062.600 1540.470 1062.740 ;
        RECT 1540.150 1062.540 1540.470 1062.600 ;
        RECT 1540.150 1027.720 1540.470 1027.780 ;
        RECT 1541.070 1027.720 1541.390 1027.780 ;
        RECT 1540.150 1027.580 1541.390 1027.720 ;
        RECT 1540.150 1027.520 1540.470 1027.580 ;
        RECT 1541.070 1027.520 1541.390 1027.580 ;
        RECT 1540.150 980.120 1540.470 980.180 ;
        RECT 1539.955 979.980 1540.470 980.120 ;
        RECT 1540.150 979.920 1540.470 979.980 ;
        RECT 1540.150 966.180 1540.470 966.240 ;
        RECT 1539.955 966.040 1540.470 966.180 ;
        RECT 1540.150 965.980 1540.470 966.040 ;
        RECT 1540.610 917.900 1540.930 917.960 ;
        RECT 1541.530 917.900 1541.850 917.960 ;
        RECT 1540.610 917.760 1541.850 917.900 ;
        RECT 1540.610 917.700 1540.930 917.760 ;
        RECT 1541.530 917.700 1541.850 917.760 ;
        RECT 1540.150 869.620 1540.470 869.680 ;
        RECT 1541.070 869.620 1541.390 869.680 ;
        RECT 1540.150 869.480 1541.390 869.620 ;
        RECT 1540.150 869.420 1540.470 869.480 ;
        RECT 1541.070 869.420 1541.390 869.480 ;
        RECT 1540.165 807.060 1540.455 807.105 ;
        RECT 1540.610 807.060 1540.930 807.120 ;
        RECT 1540.165 806.920 1540.930 807.060 ;
        RECT 1540.165 806.875 1540.455 806.920 ;
        RECT 1540.610 806.860 1540.930 806.920 ;
        RECT 1540.150 759.120 1540.470 759.180 ;
        RECT 1539.955 758.980 1540.470 759.120 ;
        RECT 1540.150 758.920 1540.470 758.980 ;
        RECT 1540.610 669.700 1540.930 669.760 ;
        RECT 1541.070 669.700 1541.390 669.760 ;
        RECT 1540.610 669.560 1541.390 669.700 ;
        RECT 1540.610 669.500 1540.930 669.560 ;
        RECT 1541.070 669.500 1541.390 669.560 ;
        RECT 1540.150 517.380 1540.470 517.440 ;
        RECT 1540.610 517.380 1540.930 517.440 ;
        RECT 1540.150 517.240 1540.930 517.380 ;
        RECT 1540.150 517.180 1540.470 517.240 ;
        RECT 1540.610 517.180 1540.930 517.240 ;
        RECT 1539.690 420.820 1540.010 420.880 ;
        RECT 1539.495 420.680 1540.010 420.820 ;
        RECT 1539.690 420.620 1540.010 420.680 ;
        RECT 1539.705 372.880 1539.995 372.925 ;
        RECT 1540.610 372.880 1540.930 372.940 ;
        RECT 1539.705 372.740 1540.930 372.880 ;
        RECT 1539.705 372.695 1539.995 372.740 ;
        RECT 1540.610 372.680 1540.930 372.740 ;
        RECT 1540.150 331.400 1540.470 331.460 ;
        RECT 1539.955 331.260 1540.470 331.400 ;
        RECT 1540.150 331.200 1540.470 331.260 ;
        RECT 1540.150 324.600 1540.470 324.660 ;
        RECT 1539.955 324.460 1540.470 324.600 ;
        RECT 1540.150 324.400 1540.470 324.460 ;
        RECT 1539.690 172.620 1540.010 172.680 ;
        RECT 1540.610 172.620 1540.930 172.680 ;
        RECT 1539.690 172.480 1540.930 172.620 ;
        RECT 1539.690 172.420 1540.010 172.480 ;
        RECT 1540.610 172.420 1540.930 172.480 ;
        RECT 1540.610 97.480 1540.930 97.540 ;
        RECT 1540.415 97.340 1540.930 97.480 ;
        RECT 1540.610 97.280 1540.930 97.340 ;
        RECT 1055.310 64.840 1055.630 64.900 ;
        RECT 1540.625 64.840 1540.915 64.885 ;
        RECT 1055.310 64.700 1540.915 64.840 ;
        RECT 1055.310 64.640 1055.630 64.700 ;
        RECT 1540.625 64.655 1540.915 64.700 ;
        RECT 1049.330 34.580 1049.650 34.640 ;
        RECT 1055.310 34.580 1055.630 34.640 ;
        RECT 1049.330 34.440 1055.630 34.580 ;
        RECT 1049.330 34.380 1049.650 34.440 ;
        RECT 1055.310 34.380 1055.630 34.440 ;
      LAYER via ;
        RECT 1540.640 1642.240 1540.900 1642.500 ;
        RECT 1543.400 1642.240 1543.660 1642.500 ;
        RECT 1540.180 1545.340 1540.440 1545.600 ;
        RECT 1541.100 1545.340 1541.360 1545.600 ;
        RECT 1540.640 1490.260 1540.900 1490.520 ;
        RECT 1541.100 1490.260 1541.360 1490.520 ;
        RECT 1539.720 1393.700 1539.980 1393.960 ;
        RECT 1541.100 1393.700 1541.360 1393.960 ;
        RECT 1539.720 1352.220 1539.980 1352.480 ;
        RECT 1539.720 1290.340 1539.980 1290.600 ;
        RECT 1539.720 1255.660 1539.980 1255.920 ;
        RECT 1540.180 1220.980 1540.440 1221.240 ;
        RECT 1540.180 1159.780 1540.440 1160.040 ;
        RECT 1540.180 1159.100 1540.440 1159.360 ;
        RECT 1540.180 1087.020 1540.440 1087.280 ;
        RECT 1540.180 1062.540 1540.440 1062.800 ;
        RECT 1540.180 1027.520 1540.440 1027.780 ;
        RECT 1541.100 1027.520 1541.360 1027.780 ;
        RECT 1540.180 979.920 1540.440 980.180 ;
        RECT 1540.180 965.980 1540.440 966.240 ;
        RECT 1540.640 917.700 1540.900 917.960 ;
        RECT 1541.560 917.700 1541.820 917.960 ;
        RECT 1540.180 869.420 1540.440 869.680 ;
        RECT 1541.100 869.420 1541.360 869.680 ;
        RECT 1540.640 806.860 1540.900 807.120 ;
        RECT 1540.180 758.920 1540.440 759.180 ;
        RECT 1540.640 669.500 1540.900 669.760 ;
        RECT 1541.100 669.500 1541.360 669.760 ;
        RECT 1540.180 517.180 1540.440 517.440 ;
        RECT 1540.640 517.180 1540.900 517.440 ;
        RECT 1539.720 420.620 1539.980 420.880 ;
        RECT 1540.640 372.680 1540.900 372.940 ;
        RECT 1540.180 331.200 1540.440 331.460 ;
        RECT 1540.180 324.400 1540.440 324.660 ;
        RECT 1539.720 172.420 1539.980 172.680 ;
        RECT 1540.640 172.420 1540.900 172.680 ;
        RECT 1540.640 97.280 1540.900 97.540 ;
        RECT 1055.340 64.640 1055.600 64.900 ;
        RECT 1049.360 34.380 1049.620 34.640 ;
        RECT 1055.340 34.380 1055.600 34.640 ;
      LAYER met2 ;
        RECT 1544.705 1700.410 1544.985 1704.000 ;
        RECT 1543.460 1700.270 1544.985 1700.410 ;
        RECT 1543.460 1642.530 1543.600 1700.270 ;
        RECT 1544.705 1700.000 1544.985 1700.270 ;
        RECT 1540.640 1642.210 1540.900 1642.530 ;
        RECT 1543.400 1642.210 1543.660 1642.530 ;
        RECT 1540.700 1559.650 1540.840 1642.210 ;
        RECT 1540.240 1559.510 1540.840 1559.650 ;
        RECT 1540.240 1545.630 1540.380 1559.510 ;
        RECT 1540.180 1545.310 1540.440 1545.630 ;
        RECT 1541.100 1545.310 1541.360 1545.630 ;
        RECT 1541.160 1514.770 1541.300 1545.310 ;
        RECT 1540.700 1514.630 1541.300 1514.770 ;
        RECT 1540.700 1490.550 1540.840 1514.630 ;
        RECT 1540.640 1490.230 1540.900 1490.550 ;
        RECT 1541.100 1490.230 1541.360 1490.550 ;
        RECT 1541.160 1393.990 1541.300 1490.230 ;
        RECT 1539.720 1393.670 1539.980 1393.990 ;
        RECT 1541.100 1393.670 1541.360 1393.990 ;
        RECT 1539.780 1352.510 1539.920 1393.670 ;
        RECT 1539.720 1352.190 1539.980 1352.510 ;
        RECT 1539.720 1290.310 1539.980 1290.630 ;
        RECT 1539.780 1255.950 1539.920 1290.310 ;
        RECT 1539.720 1255.630 1539.980 1255.950 ;
        RECT 1540.180 1220.950 1540.440 1221.270 ;
        RECT 1540.240 1160.070 1540.380 1220.950 ;
        RECT 1540.180 1159.750 1540.440 1160.070 ;
        RECT 1540.180 1159.070 1540.440 1159.390 ;
        RECT 1540.240 1087.310 1540.380 1159.070 ;
        RECT 1540.180 1086.990 1540.440 1087.310 ;
        RECT 1540.180 1062.685 1540.440 1062.830 ;
        RECT 1540.170 1062.315 1540.450 1062.685 ;
        RECT 1541.090 1062.315 1541.370 1062.685 ;
        RECT 1541.160 1027.810 1541.300 1062.315 ;
        RECT 1540.180 1027.490 1540.440 1027.810 ;
        RECT 1541.100 1027.490 1541.360 1027.810 ;
        RECT 1540.240 980.210 1540.380 1027.490 ;
        RECT 1540.180 979.890 1540.440 980.210 ;
        RECT 1540.180 966.125 1540.440 966.270 ;
        RECT 1540.170 965.755 1540.450 966.125 ;
        RECT 1541.550 965.755 1541.830 966.125 ;
        RECT 1541.620 917.990 1541.760 965.755 ;
        RECT 1540.640 917.670 1540.900 917.990 ;
        RECT 1541.560 917.670 1541.820 917.990 ;
        RECT 1540.700 893.930 1540.840 917.670 ;
        RECT 1540.700 893.790 1541.300 893.930 ;
        RECT 1541.160 869.710 1541.300 893.790 ;
        RECT 1540.180 869.390 1540.440 869.710 ;
        RECT 1541.100 869.390 1541.360 869.710 ;
        RECT 1540.240 814.370 1540.380 869.390 ;
        RECT 1540.240 814.230 1540.840 814.370 ;
        RECT 1540.700 807.150 1540.840 814.230 ;
        RECT 1540.640 806.830 1540.900 807.150 ;
        RECT 1540.180 758.890 1540.440 759.210 ;
        RECT 1540.240 741.610 1540.380 758.890 ;
        RECT 1540.240 741.470 1541.300 741.610 ;
        RECT 1541.160 669.790 1541.300 741.470 ;
        RECT 1540.640 669.470 1540.900 669.790 ;
        RECT 1541.100 669.470 1541.360 669.790 ;
        RECT 1540.700 621.250 1540.840 669.470 ;
        RECT 1540.240 621.110 1540.840 621.250 ;
        RECT 1540.240 541.690 1540.380 621.110 ;
        RECT 1540.240 541.550 1541.300 541.690 ;
        RECT 1541.160 524.010 1541.300 541.550 ;
        RECT 1540.700 523.870 1541.300 524.010 ;
        RECT 1540.700 517.470 1540.840 523.870 ;
        RECT 1540.180 517.150 1540.440 517.470 ;
        RECT 1540.640 517.150 1540.900 517.470 ;
        RECT 1540.240 492.730 1540.380 517.150 ;
        RECT 1540.240 492.590 1540.840 492.730 ;
        RECT 1540.700 435.045 1540.840 492.590 ;
        RECT 1539.710 434.675 1539.990 435.045 ;
        RECT 1540.630 434.675 1540.910 435.045 ;
        RECT 1539.780 420.910 1539.920 434.675 ;
        RECT 1539.720 420.590 1539.980 420.910 ;
        RECT 1540.640 372.650 1540.900 372.970 ;
        RECT 1540.700 372.370 1540.840 372.650 ;
        RECT 1540.240 372.230 1540.840 372.370 ;
        RECT 1540.240 331.490 1540.380 372.230 ;
        RECT 1540.180 331.170 1540.440 331.490 ;
        RECT 1540.180 324.370 1540.440 324.690 ;
        RECT 1540.240 324.090 1540.380 324.370 ;
        RECT 1540.240 323.950 1541.300 324.090 ;
        RECT 1541.160 282.610 1541.300 323.950 ;
        RECT 1540.700 282.470 1541.300 282.610 ;
        RECT 1540.700 252.010 1540.840 282.470 ;
        RECT 1540.700 251.870 1541.300 252.010 ;
        RECT 1541.160 220.845 1541.300 251.870 ;
        RECT 1539.710 220.475 1539.990 220.845 ;
        RECT 1541.090 220.475 1541.370 220.845 ;
        RECT 1539.780 172.710 1539.920 220.475 ;
        RECT 1539.720 172.390 1539.980 172.710 ;
        RECT 1540.640 172.390 1540.900 172.710 ;
        RECT 1540.700 97.570 1540.840 172.390 ;
        RECT 1540.640 97.250 1540.900 97.570 ;
        RECT 1055.340 64.610 1055.600 64.930 ;
        RECT 1055.400 34.670 1055.540 64.610 ;
        RECT 1049.360 34.350 1049.620 34.670 ;
        RECT 1055.340 34.350 1055.600 34.670 ;
        RECT 1049.420 2.400 1049.560 34.350 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
      LAYER via2 ;
        RECT 1540.170 1062.360 1540.450 1062.640 ;
        RECT 1541.090 1062.360 1541.370 1062.640 ;
        RECT 1540.170 965.800 1540.450 966.080 ;
        RECT 1541.550 965.800 1541.830 966.080 ;
        RECT 1539.710 434.720 1539.990 435.000 ;
        RECT 1540.630 434.720 1540.910 435.000 ;
        RECT 1539.710 220.520 1539.990 220.800 ;
        RECT 1541.090 220.520 1541.370 220.800 ;
      LAYER met3 ;
        RECT 1540.145 1062.650 1540.475 1062.665 ;
        RECT 1541.065 1062.650 1541.395 1062.665 ;
        RECT 1540.145 1062.350 1541.395 1062.650 ;
        RECT 1540.145 1062.335 1540.475 1062.350 ;
        RECT 1541.065 1062.335 1541.395 1062.350 ;
        RECT 1540.145 966.090 1540.475 966.105 ;
        RECT 1541.525 966.090 1541.855 966.105 ;
        RECT 1540.145 965.790 1541.855 966.090 ;
        RECT 1540.145 965.775 1540.475 965.790 ;
        RECT 1541.525 965.775 1541.855 965.790 ;
        RECT 1539.685 435.010 1540.015 435.025 ;
        RECT 1540.605 435.010 1540.935 435.025 ;
        RECT 1539.685 434.710 1540.935 435.010 ;
        RECT 1539.685 434.695 1540.015 434.710 ;
        RECT 1540.605 434.695 1540.935 434.710 ;
        RECT 1539.685 220.810 1540.015 220.825 ;
        RECT 1541.065 220.810 1541.395 220.825 ;
        RECT 1539.685 220.510 1541.395 220.810 ;
        RECT 1539.685 220.495 1540.015 220.510 ;
        RECT 1541.065 220.495 1541.395 220.510 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1547.125 1338.665 1547.295 1366.035 ;
        RECT 1547.585 697.085 1547.755 745.195 ;
        RECT 1546.665 512.125 1546.835 576.215 ;
        RECT 1547.125 427.805 1547.295 449.055 ;
      LAYER mcon ;
        RECT 1547.125 1365.865 1547.295 1366.035 ;
        RECT 1547.585 745.025 1547.755 745.195 ;
        RECT 1546.665 576.045 1546.835 576.215 ;
        RECT 1547.125 448.885 1547.295 449.055 ;
      LAYER met1 ;
        RECT 1547.050 1366.020 1547.370 1366.080 ;
        RECT 1546.855 1365.880 1547.370 1366.020 ;
        RECT 1547.050 1365.820 1547.370 1365.880 ;
        RECT 1547.050 1338.820 1547.370 1338.880 ;
        RECT 1546.855 1338.680 1547.370 1338.820 ;
        RECT 1547.050 1338.620 1547.370 1338.680 ;
        RECT 1546.590 1007.120 1546.910 1007.380 ;
        RECT 1546.680 1006.980 1546.820 1007.120 ;
        RECT 1547.050 1006.980 1547.370 1007.040 ;
        RECT 1546.680 1006.840 1547.370 1006.980 ;
        RECT 1547.050 1006.780 1547.370 1006.840 ;
        RECT 1547.510 745.180 1547.830 745.240 ;
        RECT 1547.315 745.040 1547.830 745.180 ;
        RECT 1547.510 744.980 1547.830 745.040 ;
        RECT 1547.510 697.240 1547.830 697.300 ;
        RECT 1547.315 697.100 1547.830 697.240 ;
        RECT 1547.510 697.040 1547.830 697.100 ;
        RECT 1547.510 672.760 1547.830 672.820 ;
        RECT 1548.430 672.760 1548.750 672.820 ;
        RECT 1547.510 672.620 1548.750 672.760 ;
        RECT 1547.510 672.560 1547.830 672.620 ;
        RECT 1548.430 672.560 1548.750 672.620 ;
        RECT 1547.050 600.680 1547.370 600.740 ;
        RECT 1548.430 600.680 1548.750 600.740 ;
        RECT 1547.050 600.540 1548.750 600.680 ;
        RECT 1547.050 600.480 1547.370 600.540 ;
        RECT 1548.430 600.480 1548.750 600.540 ;
        RECT 1546.590 576.200 1546.910 576.260 ;
        RECT 1546.395 576.060 1546.910 576.200 ;
        RECT 1546.590 576.000 1546.910 576.060 ;
        RECT 1546.590 512.280 1546.910 512.340 ;
        RECT 1546.395 512.140 1546.910 512.280 ;
        RECT 1546.590 512.080 1546.910 512.140 ;
        RECT 1547.050 449.040 1547.370 449.100 ;
        RECT 1546.855 448.900 1547.370 449.040 ;
        RECT 1547.050 448.840 1547.370 448.900 ;
        RECT 1547.050 427.960 1547.370 428.020 ;
        RECT 1546.855 427.820 1547.370 427.960 ;
        RECT 1547.050 427.760 1547.370 427.820 ;
        RECT 1546.590 331.060 1546.910 331.120 ;
        RECT 1547.050 331.060 1547.370 331.120 ;
        RECT 1546.590 330.920 1547.370 331.060 ;
        RECT 1546.590 330.860 1546.910 330.920 ;
        RECT 1547.050 330.860 1547.370 330.920 ;
        RECT 1547.050 282.920 1547.370 283.180 ;
        RECT 1547.140 282.440 1547.280 282.920 ;
        RECT 1547.510 282.440 1547.830 282.500 ;
        RECT 1547.140 282.300 1547.830 282.440 ;
        RECT 1547.510 282.240 1547.830 282.300 ;
        RECT 1069.110 64.500 1069.430 64.560 ;
        RECT 1546.590 64.500 1546.910 64.560 ;
        RECT 1069.110 64.360 1546.910 64.500 ;
        RECT 1069.110 64.300 1069.430 64.360 ;
        RECT 1546.590 64.300 1546.910 64.360 ;
      LAYER via ;
        RECT 1547.080 1365.820 1547.340 1366.080 ;
        RECT 1547.080 1338.620 1547.340 1338.880 ;
        RECT 1546.620 1007.120 1546.880 1007.380 ;
        RECT 1547.080 1006.780 1547.340 1007.040 ;
        RECT 1547.540 744.980 1547.800 745.240 ;
        RECT 1547.540 697.040 1547.800 697.300 ;
        RECT 1547.540 672.560 1547.800 672.820 ;
        RECT 1548.460 672.560 1548.720 672.820 ;
        RECT 1547.080 600.480 1547.340 600.740 ;
        RECT 1548.460 600.480 1548.720 600.740 ;
        RECT 1546.620 576.000 1546.880 576.260 ;
        RECT 1546.620 512.080 1546.880 512.340 ;
        RECT 1547.080 448.840 1547.340 449.100 ;
        RECT 1547.080 427.760 1547.340 428.020 ;
        RECT 1546.620 330.860 1546.880 331.120 ;
        RECT 1547.080 330.860 1547.340 331.120 ;
        RECT 1547.080 282.920 1547.340 283.180 ;
        RECT 1547.540 282.240 1547.800 282.500 ;
        RECT 1069.140 64.300 1069.400 64.560 ;
        RECT 1546.620 64.300 1546.880 64.560 ;
      LAYER met2 ;
        RECT 1551.605 1700.410 1551.885 1704.000 ;
        RECT 1550.820 1700.270 1551.885 1700.410 ;
        RECT 1550.820 1642.725 1550.960 1700.270 ;
        RECT 1551.605 1700.000 1551.885 1700.270 ;
        RECT 1550.750 1642.355 1551.030 1642.725 ;
        RECT 1547.070 1641.675 1547.350 1642.045 ;
        RECT 1547.140 1366.110 1547.280 1641.675 ;
        RECT 1547.080 1365.790 1547.340 1366.110 ;
        RECT 1547.080 1338.590 1547.340 1338.910 ;
        RECT 1547.140 1269.970 1547.280 1338.590 ;
        RECT 1546.680 1269.830 1547.280 1269.970 ;
        RECT 1546.680 1269.290 1546.820 1269.830 ;
        RECT 1546.680 1269.150 1547.280 1269.290 ;
        RECT 1547.140 1076.850 1547.280 1269.150 ;
        RECT 1546.680 1076.710 1547.280 1076.850 ;
        RECT 1546.680 1076.170 1546.820 1076.710 ;
        RECT 1546.680 1076.030 1547.280 1076.170 ;
        RECT 1547.140 1028.570 1547.280 1076.030 ;
        RECT 1547.140 1028.430 1547.740 1028.570 ;
        RECT 1547.600 1007.605 1547.740 1028.430 ;
        RECT 1546.610 1007.235 1546.890 1007.605 ;
        RECT 1547.530 1007.235 1547.810 1007.605 ;
        RECT 1546.620 1007.090 1546.880 1007.235 ;
        RECT 1547.080 1006.750 1547.340 1007.070 ;
        RECT 1547.140 883.730 1547.280 1006.750 ;
        RECT 1546.680 883.590 1547.280 883.730 ;
        RECT 1546.680 883.050 1546.820 883.590 ;
        RECT 1546.680 882.910 1547.280 883.050 ;
        RECT 1547.140 751.810 1547.280 882.910 ;
        RECT 1547.140 751.670 1547.740 751.810 ;
        RECT 1547.600 745.270 1547.740 751.670 ;
        RECT 1547.540 744.950 1547.800 745.270 ;
        RECT 1547.540 697.010 1547.800 697.330 ;
        RECT 1547.600 672.850 1547.740 697.010 ;
        RECT 1547.540 672.530 1547.800 672.850 ;
        RECT 1548.460 672.530 1548.720 672.850 ;
        RECT 1548.520 600.770 1548.660 672.530 ;
        RECT 1547.080 600.450 1547.340 600.770 ;
        RECT 1548.460 600.450 1548.720 600.770 ;
        RECT 1547.140 600.170 1547.280 600.450 ;
        RECT 1546.680 600.030 1547.280 600.170 ;
        RECT 1546.680 576.290 1546.820 600.030 ;
        RECT 1546.620 575.970 1546.880 576.290 ;
        RECT 1546.620 512.050 1546.880 512.370 ;
        RECT 1546.680 486.610 1546.820 512.050 ;
        RECT 1546.680 486.470 1547.280 486.610 ;
        RECT 1547.140 449.130 1547.280 486.470 ;
        RECT 1547.080 448.810 1547.340 449.130 ;
        RECT 1547.080 427.730 1547.340 428.050 ;
        RECT 1547.140 400.930 1547.280 427.730 ;
        RECT 1547.140 400.790 1547.740 400.930 ;
        RECT 1547.600 379.340 1547.740 400.790 ;
        RECT 1546.680 379.200 1547.740 379.340 ;
        RECT 1546.680 331.150 1546.820 379.200 ;
        RECT 1546.620 330.830 1546.880 331.150 ;
        RECT 1547.080 330.830 1547.340 331.150 ;
        RECT 1547.140 283.210 1547.280 330.830 ;
        RECT 1547.080 282.890 1547.340 283.210 ;
        RECT 1547.540 282.210 1547.800 282.530 ;
        RECT 1547.600 154.770 1547.740 282.210 ;
        RECT 1546.680 154.630 1547.740 154.770 ;
        RECT 1546.680 64.590 1546.820 154.630 ;
        RECT 1069.140 64.270 1069.400 64.590 ;
        RECT 1546.620 64.270 1546.880 64.590 ;
        RECT 1069.200 3.130 1069.340 64.270 ;
        RECT 1067.360 2.990 1069.340 3.130 ;
        RECT 1067.360 2.400 1067.500 2.990 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
      LAYER via2 ;
        RECT 1550.750 1642.400 1551.030 1642.680 ;
        RECT 1547.070 1641.720 1547.350 1642.000 ;
        RECT 1546.610 1007.280 1546.890 1007.560 ;
        RECT 1547.530 1007.280 1547.810 1007.560 ;
      LAYER met3 ;
        RECT 1550.725 1642.690 1551.055 1642.705 ;
        RECT 1546.830 1642.390 1551.055 1642.690 ;
        RECT 1546.830 1642.025 1547.130 1642.390 ;
        RECT 1550.725 1642.375 1551.055 1642.390 ;
        RECT 1546.830 1641.710 1547.375 1642.025 ;
        RECT 1547.045 1641.695 1547.375 1641.710 ;
        RECT 1546.585 1007.570 1546.915 1007.585 ;
        RECT 1547.505 1007.570 1547.835 1007.585 ;
        RECT 1546.585 1007.270 1547.835 1007.570 ;
        RECT 1546.585 1007.255 1546.915 1007.270 ;
        RECT 1547.505 1007.255 1547.835 1007.270 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1554.025 1483.505 1554.195 1490.815 ;
        RECT 1553.565 1339.005 1553.735 1367.055 ;
        RECT 1554.025 1199.945 1554.195 1283.415 ;
        RECT 1554.485 1072.785 1554.655 1097.095 ;
        RECT 1554.025 927.945 1554.195 1000.535 ;
        RECT 1554.025 848.725 1554.195 896.835 ;
        RECT 1554.025 620.925 1554.195 669.375 ;
      LAYER mcon ;
        RECT 1554.025 1490.645 1554.195 1490.815 ;
        RECT 1553.565 1366.885 1553.735 1367.055 ;
        RECT 1554.025 1283.245 1554.195 1283.415 ;
        RECT 1554.485 1096.925 1554.655 1097.095 ;
        RECT 1554.025 1000.365 1554.195 1000.535 ;
        RECT 1554.025 896.665 1554.195 896.835 ;
        RECT 1554.025 669.205 1554.195 669.375 ;
      LAYER met1 ;
        RECT 1554.410 1642.440 1554.730 1642.500 ;
        RECT 1557.170 1642.440 1557.490 1642.500 ;
        RECT 1554.410 1642.300 1557.490 1642.440 ;
        RECT 1554.410 1642.240 1554.730 1642.300 ;
        RECT 1557.170 1642.240 1557.490 1642.300 ;
        RECT 1553.965 1490.800 1554.255 1490.845 ;
        RECT 1554.410 1490.800 1554.730 1490.860 ;
        RECT 1553.965 1490.660 1554.730 1490.800 ;
        RECT 1553.965 1490.615 1554.255 1490.660 ;
        RECT 1554.410 1490.600 1554.730 1490.660 ;
        RECT 1553.950 1483.660 1554.270 1483.720 ;
        RECT 1553.755 1483.520 1554.270 1483.660 ;
        RECT 1553.950 1483.460 1554.270 1483.520 ;
        RECT 1553.950 1478.900 1554.270 1478.960 ;
        RECT 1554.870 1478.900 1555.190 1478.960 ;
        RECT 1553.950 1478.760 1555.190 1478.900 ;
        RECT 1553.950 1478.700 1554.270 1478.760 ;
        RECT 1554.870 1478.700 1555.190 1478.760 ;
        RECT 1553.490 1387.100 1553.810 1387.160 ;
        RECT 1553.950 1387.100 1554.270 1387.160 ;
        RECT 1553.490 1386.960 1554.270 1387.100 ;
        RECT 1553.490 1386.900 1553.810 1386.960 ;
        RECT 1553.950 1386.900 1554.270 1386.960 ;
        RECT 1553.490 1367.040 1553.810 1367.100 ;
        RECT 1553.295 1366.900 1553.810 1367.040 ;
        RECT 1553.490 1366.840 1553.810 1366.900 ;
        RECT 1553.505 1339.160 1553.795 1339.205 ;
        RECT 1553.950 1339.160 1554.270 1339.220 ;
        RECT 1553.505 1339.020 1554.270 1339.160 ;
        RECT 1553.505 1338.975 1553.795 1339.020 ;
        RECT 1553.950 1338.960 1554.270 1339.020 ;
        RECT 1553.950 1318.220 1554.270 1318.480 ;
        RECT 1554.040 1317.800 1554.180 1318.220 ;
        RECT 1553.950 1317.540 1554.270 1317.800 ;
        RECT 1553.965 1283.400 1554.255 1283.445 ;
        RECT 1554.410 1283.400 1554.730 1283.460 ;
        RECT 1553.965 1283.260 1554.730 1283.400 ;
        RECT 1553.965 1283.215 1554.255 1283.260 ;
        RECT 1554.410 1283.200 1554.730 1283.260 ;
        RECT 1553.950 1200.100 1554.270 1200.160 ;
        RECT 1553.755 1199.960 1554.270 1200.100 ;
        RECT 1553.950 1199.900 1554.270 1199.960 ;
        RECT 1553.490 1193.640 1553.810 1193.700 ;
        RECT 1553.950 1193.640 1554.270 1193.700 ;
        RECT 1553.490 1193.500 1554.270 1193.640 ;
        RECT 1553.490 1193.440 1553.810 1193.500 ;
        RECT 1553.950 1193.440 1554.270 1193.500 ;
        RECT 1554.410 1097.080 1554.730 1097.140 ;
        RECT 1554.215 1096.940 1554.730 1097.080 ;
        RECT 1554.410 1096.880 1554.730 1096.940 ;
        RECT 1554.410 1072.940 1554.730 1073.000 ;
        RECT 1554.215 1072.800 1554.730 1072.940 ;
        RECT 1554.410 1072.740 1554.730 1072.800 ;
        RECT 1553.950 1007.320 1554.270 1007.380 ;
        RECT 1554.410 1007.320 1554.730 1007.380 ;
        RECT 1553.950 1007.180 1554.730 1007.320 ;
        RECT 1553.950 1007.120 1554.270 1007.180 ;
        RECT 1554.410 1007.120 1554.730 1007.180 ;
        RECT 1553.950 1000.520 1554.270 1000.580 ;
        RECT 1553.755 1000.380 1554.270 1000.520 ;
        RECT 1553.950 1000.320 1554.270 1000.380 ;
        RECT 1552.110 928.100 1552.430 928.160 ;
        RECT 1553.965 928.100 1554.255 928.145 ;
        RECT 1552.110 927.960 1554.255 928.100 ;
        RECT 1552.110 927.900 1552.430 927.960 ;
        RECT 1553.965 927.915 1554.255 927.960 ;
        RECT 1553.950 896.820 1554.270 896.880 ;
        RECT 1553.755 896.680 1554.270 896.820 ;
        RECT 1553.950 896.620 1554.270 896.680 ;
        RECT 1553.965 848.880 1554.255 848.925 ;
        RECT 1554.410 848.880 1554.730 848.940 ;
        RECT 1553.965 848.740 1554.730 848.880 ;
        RECT 1553.965 848.695 1554.255 848.740 ;
        RECT 1554.410 848.680 1554.730 848.740 ;
        RECT 1554.410 807.060 1554.730 807.120 ;
        RECT 1554.870 807.060 1555.190 807.120 ;
        RECT 1554.410 806.920 1555.190 807.060 ;
        RECT 1554.410 806.860 1554.730 806.920 ;
        RECT 1554.870 806.860 1555.190 806.920 ;
        RECT 1553.950 669.360 1554.270 669.420 ;
        RECT 1553.755 669.220 1554.270 669.360 ;
        RECT 1553.950 669.160 1554.270 669.220 ;
        RECT 1553.950 621.080 1554.270 621.140 ;
        RECT 1553.755 620.940 1554.270 621.080 ;
        RECT 1553.950 620.880 1554.270 620.940 ;
        RECT 1553.950 572.940 1554.270 573.200 ;
        RECT 1554.040 572.460 1554.180 572.940 ;
        RECT 1554.410 572.460 1554.730 572.520 ;
        RECT 1554.040 572.320 1554.730 572.460 ;
        RECT 1554.410 572.260 1554.730 572.320 ;
        RECT 1554.410 517.380 1554.730 517.440 ;
        RECT 1555.330 517.380 1555.650 517.440 ;
        RECT 1554.410 517.240 1555.650 517.380 ;
        RECT 1554.410 517.180 1554.730 517.240 ;
        RECT 1555.330 517.180 1555.650 517.240 ;
        RECT 1554.410 324.600 1554.730 324.660 ;
        RECT 1554.870 324.600 1555.190 324.660 ;
        RECT 1554.410 324.460 1555.190 324.600 ;
        RECT 1554.410 324.400 1554.730 324.460 ;
        RECT 1554.870 324.400 1555.190 324.460 ;
        RECT 1553.950 294.000 1554.270 294.060 ;
        RECT 1554.870 294.000 1555.190 294.060 ;
        RECT 1553.950 293.860 1555.190 294.000 ;
        RECT 1553.950 293.800 1554.270 293.860 ;
        RECT 1554.870 293.800 1555.190 293.860 ;
        RECT 1553.950 90.340 1554.270 90.400 ;
        RECT 1553.580 90.200 1554.270 90.340 ;
        RECT 1553.580 90.060 1553.720 90.200 ;
        RECT 1553.950 90.140 1554.270 90.200 ;
        RECT 1553.490 89.800 1553.810 90.060 ;
        RECT 1089.810 64.160 1090.130 64.220 ;
        RECT 1553.490 64.160 1553.810 64.220 ;
        RECT 1089.810 64.020 1553.810 64.160 ;
        RECT 1089.810 63.960 1090.130 64.020 ;
        RECT 1553.490 63.960 1553.810 64.020 ;
        RECT 1085.210 2.960 1085.530 3.020 ;
        RECT 1089.810 2.960 1090.130 3.020 ;
        RECT 1085.210 2.820 1090.130 2.960 ;
        RECT 1085.210 2.760 1085.530 2.820 ;
        RECT 1089.810 2.760 1090.130 2.820 ;
      LAYER via ;
        RECT 1554.440 1642.240 1554.700 1642.500 ;
        RECT 1557.200 1642.240 1557.460 1642.500 ;
        RECT 1554.440 1490.600 1554.700 1490.860 ;
        RECT 1553.980 1483.460 1554.240 1483.720 ;
        RECT 1553.980 1478.700 1554.240 1478.960 ;
        RECT 1554.900 1478.700 1555.160 1478.960 ;
        RECT 1553.520 1386.900 1553.780 1387.160 ;
        RECT 1553.980 1386.900 1554.240 1387.160 ;
        RECT 1553.520 1366.840 1553.780 1367.100 ;
        RECT 1553.980 1338.960 1554.240 1339.220 ;
        RECT 1553.980 1318.220 1554.240 1318.480 ;
        RECT 1553.980 1317.540 1554.240 1317.800 ;
        RECT 1554.440 1283.200 1554.700 1283.460 ;
        RECT 1553.980 1199.900 1554.240 1200.160 ;
        RECT 1553.520 1193.440 1553.780 1193.700 ;
        RECT 1553.980 1193.440 1554.240 1193.700 ;
        RECT 1554.440 1096.880 1554.700 1097.140 ;
        RECT 1554.440 1072.740 1554.700 1073.000 ;
        RECT 1553.980 1007.120 1554.240 1007.380 ;
        RECT 1554.440 1007.120 1554.700 1007.380 ;
        RECT 1553.980 1000.320 1554.240 1000.580 ;
        RECT 1552.140 927.900 1552.400 928.160 ;
        RECT 1553.980 896.620 1554.240 896.880 ;
        RECT 1554.440 848.680 1554.700 848.940 ;
        RECT 1554.440 806.860 1554.700 807.120 ;
        RECT 1554.900 806.860 1555.160 807.120 ;
        RECT 1553.980 669.160 1554.240 669.420 ;
        RECT 1553.980 620.880 1554.240 621.140 ;
        RECT 1553.980 572.940 1554.240 573.200 ;
        RECT 1554.440 572.260 1554.700 572.520 ;
        RECT 1554.440 517.180 1554.700 517.440 ;
        RECT 1555.360 517.180 1555.620 517.440 ;
        RECT 1554.440 324.400 1554.700 324.660 ;
        RECT 1554.900 324.400 1555.160 324.660 ;
        RECT 1553.980 293.800 1554.240 294.060 ;
        RECT 1554.900 293.800 1555.160 294.060 ;
        RECT 1553.980 90.140 1554.240 90.400 ;
        RECT 1553.520 89.800 1553.780 90.060 ;
        RECT 1089.840 63.960 1090.100 64.220 ;
        RECT 1553.520 63.960 1553.780 64.220 ;
        RECT 1085.240 2.760 1085.500 3.020 ;
        RECT 1089.840 2.760 1090.100 3.020 ;
      LAYER met2 ;
        RECT 1558.505 1700.410 1558.785 1704.000 ;
        RECT 1557.260 1700.270 1558.785 1700.410 ;
        RECT 1557.260 1642.530 1557.400 1700.270 ;
        RECT 1558.505 1700.000 1558.785 1700.270 ;
        RECT 1554.440 1642.210 1554.700 1642.530 ;
        RECT 1557.200 1642.210 1557.460 1642.530 ;
        RECT 1554.500 1592.970 1554.640 1642.210 ;
        RECT 1554.040 1592.830 1554.640 1592.970 ;
        RECT 1554.040 1580.165 1554.180 1592.830 ;
        RECT 1553.970 1579.795 1554.250 1580.165 ;
        RECT 1554.430 1579.115 1554.710 1579.485 ;
        RECT 1554.500 1490.890 1554.640 1579.115 ;
        RECT 1554.440 1490.570 1554.700 1490.890 ;
        RECT 1553.980 1483.430 1554.240 1483.750 ;
        RECT 1554.040 1478.990 1554.180 1483.430 ;
        RECT 1553.980 1478.670 1554.240 1478.990 ;
        RECT 1554.900 1478.670 1555.160 1478.990 ;
        RECT 1554.960 1435.210 1555.100 1478.670 ;
        RECT 1554.040 1435.070 1555.100 1435.210 ;
        RECT 1554.040 1387.190 1554.180 1435.070 ;
        RECT 1553.520 1386.870 1553.780 1387.190 ;
        RECT 1553.980 1386.870 1554.240 1387.190 ;
        RECT 1553.580 1367.130 1553.720 1386.870 ;
        RECT 1553.520 1366.810 1553.780 1367.130 ;
        RECT 1553.980 1338.930 1554.240 1339.250 ;
        RECT 1554.040 1318.510 1554.180 1338.930 ;
        RECT 1553.980 1318.190 1554.240 1318.510 ;
        RECT 1553.980 1317.510 1554.240 1317.830 ;
        RECT 1554.040 1290.370 1554.180 1317.510 ;
        RECT 1554.040 1290.230 1554.640 1290.370 ;
        RECT 1554.500 1283.490 1554.640 1290.230 ;
        RECT 1554.440 1283.170 1554.700 1283.490 ;
        RECT 1553.980 1199.870 1554.240 1200.190 ;
        RECT 1554.040 1193.730 1554.180 1199.870 ;
        RECT 1553.520 1193.410 1553.780 1193.730 ;
        RECT 1553.980 1193.410 1554.240 1193.730 ;
        RECT 1553.580 1145.645 1553.720 1193.410 ;
        RECT 1553.510 1145.275 1553.790 1145.645 ;
        RECT 1554.890 1145.275 1555.170 1145.645 ;
        RECT 1554.960 1135.330 1555.100 1145.275 ;
        RECT 1554.500 1135.190 1555.100 1135.330 ;
        RECT 1554.500 1097.170 1554.640 1135.190 ;
        RECT 1554.440 1096.850 1554.700 1097.170 ;
        RECT 1554.440 1072.710 1554.700 1073.030 ;
        RECT 1554.500 1007.410 1554.640 1072.710 ;
        RECT 1553.980 1007.090 1554.240 1007.410 ;
        RECT 1554.440 1007.090 1554.700 1007.410 ;
        RECT 1554.040 1000.610 1554.180 1007.090 ;
        RECT 1553.980 1000.290 1554.240 1000.610 ;
        RECT 1552.140 927.870 1552.400 928.190 ;
        RECT 1552.200 904.245 1552.340 927.870 ;
        RECT 1552.130 903.875 1552.410 904.245 ;
        RECT 1553.970 903.875 1554.250 904.245 ;
        RECT 1554.040 896.910 1554.180 903.875 ;
        RECT 1553.980 896.590 1554.240 896.910 ;
        RECT 1554.440 848.650 1554.700 848.970 ;
        RECT 1554.500 807.150 1554.640 848.650 ;
        RECT 1554.440 806.830 1554.700 807.150 ;
        RECT 1554.900 806.830 1555.160 807.150 ;
        RECT 1554.960 747.730 1555.100 806.830 ;
        RECT 1554.500 747.590 1555.100 747.730 ;
        RECT 1554.500 669.530 1554.640 747.590 ;
        RECT 1554.040 669.450 1554.640 669.530 ;
        RECT 1553.980 669.390 1554.640 669.450 ;
        RECT 1553.980 669.130 1554.240 669.390 ;
        RECT 1554.040 668.975 1554.180 669.130 ;
        RECT 1553.980 620.850 1554.240 621.170 ;
        RECT 1554.040 573.230 1554.180 620.850 ;
        RECT 1553.980 572.910 1554.240 573.230 ;
        RECT 1554.440 572.230 1554.700 572.550 ;
        RECT 1554.500 517.470 1554.640 572.230 ;
        RECT 1554.440 517.150 1554.700 517.470 ;
        RECT 1555.360 517.150 1555.620 517.470 ;
        RECT 1555.420 469.725 1555.560 517.150 ;
        RECT 1555.350 469.355 1555.630 469.725 ;
        RECT 1554.890 468.675 1555.170 469.045 ;
        RECT 1554.960 372.370 1555.100 468.675 ;
        RECT 1554.500 372.230 1555.100 372.370 ;
        RECT 1554.500 324.690 1554.640 372.230 ;
        RECT 1554.440 324.370 1554.700 324.690 ;
        RECT 1554.900 324.370 1555.160 324.690 ;
        RECT 1554.960 294.090 1555.100 324.370 ;
        RECT 1553.980 293.770 1554.240 294.090 ;
        RECT 1554.900 293.770 1555.160 294.090 ;
        RECT 1554.040 258.810 1554.180 293.770 ;
        RECT 1554.040 258.670 1555.100 258.810 ;
        RECT 1554.960 186.730 1555.100 258.670 ;
        RECT 1554.040 186.590 1555.100 186.730 ;
        RECT 1554.040 90.430 1554.180 186.590 ;
        RECT 1553.980 90.110 1554.240 90.430 ;
        RECT 1553.520 89.770 1553.780 90.090 ;
        RECT 1553.580 64.250 1553.720 89.770 ;
        RECT 1089.840 63.930 1090.100 64.250 ;
        RECT 1553.520 63.930 1553.780 64.250 ;
        RECT 1089.900 3.050 1090.040 63.930 ;
        RECT 1085.240 2.730 1085.500 3.050 ;
        RECT 1089.840 2.730 1090.100 3.050 ;
        RECT 1085.300 2.400 1085.440 2.730 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
      LAYER via2 ;
        RECT 1553.970 1579.840 1554.250 1580.120 ;
        RECT 1554.430 1579.160 1554.710 1579.440 ;
        RECT 1553.510 1145.320 1553.790 1145.600 ;
        RECT 1554.890 1145.320 1555.170 1145.600 ;
        RECT 1552.130 903.920 1552.410 904.200 ;
        RECT 1553.970 903.920 1554.250 904.200 ;
        RECT 1555.350 469.400 1555.630 469.680 ;
        RECT 1554.890 468.720 1555.170 469.000 ;
      LAYER met3 ;
        RECT 1553.945 1580.130 1554.275 1580.145 ;
        RECT 1553.270 1579.830 1554.275 1580.130 ;
        RECT 1553.270 1579.450 1553.570 1579.830 ;
        RECT 1553.945 1579.815 1554.275 1579.830 ;
        RECT 1554.405 1579.450 1554.735 1579.465 ;
        RECT 1553.270 1579.150 1554.735 1579.450 ;
        RECT 1554.405 1579.135 1554.735 1579.150 ;
        RECT 1553.485 1145.610 1553.815 1145.625 ;
        RECT 1554.865 1145.610 1555.195 1145.625 ;
        RECT 1553.485 1145.310 1555.195 1145.610 ;
        RECT 1553.485 1145.295 1553.815 1145.310 ;
        RECT 1554.865 1145.295 1555.195 1145.310 ;
        RECT 1552.105 904.210 1552.435 904.225 ;
        RECT 1553.945 904.210 1554.275 904.225 ;
        RECT 1552.105 903.910 1554.275 904.210 ;
        RECT 1552.105 903.895 1552.435 903.910 ;
        RECT 1553.945 903.895 1554.275 903.910 ;
        RECT 1555.325 469.690 1555.655 469.705 ;
        RECT 1555.110 469.375 1555.655 469.690 ;
        RECT 1555.110 469.025 1555.410 469.375 ;
        RECT 1554.865 468.710 1555.410 469.025 ;
        RECT 1554.865 468.695 1555.195 468.710 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1560.850 1671.680 1561.170 1671.740 ;
        RECT 1563.150 1671.680 1563.470 1671.740 ;
        RECT 1560.850 1671.540 1563.470 1671.680 ;
        RECT 1560.850 1671.480 1561.170 1671.540 ;
        RECT 1563.150 1671.480 1563.470 1671.540 ;
        RECT 1103.610 63.820 1103.930 63.880 ;
        RECT 1560.850 63.820 1561.170 63.880 ;
        RECT 1103.610 63.680 1561.170 63.820 ;
        RECT 1103.610 63.620 1103.930 63.680 ;
        RECT 1560.850 63.620 1561.170 63.680 ;
        RECT 1102.690 2.960 1103.010 3.020 ;
        RECT 1103.610 2.960 1103.930 3.020 ;
        RECT 1102.690 2.820 1103.930 2.960 ;
        RECT 1102.690 2.760 1103.010 2.820 ;
        RECT 1103.610 2.760 1103.930 2.820 ;
      LAYER via ;
        RECT 1560.880 1671.480 1561.140 1671.740 ;
        RECT 1563.180 1671.480 1563.440 1671.740 ;
        RECT 1103.640 63.620 1103.900 63.880 ;
        RECT 1560.880 63.620 1561.140 63.880 ;
        RECT 1102.720 2.760 1102.980 3.020 ;
        RECT 1103.640 2.760 1103.900 3.020 ;
      LAYER met2 ;
        RECT 1564.945 1700.410 1565.225 1704.000 ;
        RECT 1563.240 1700.270 1565.225 1700.410 ;
        RECT 1563.240 1671.770 1563.380 1700.270 ;
        RECT 1564.945 1700.000 1565.225 1700.270 ;
        RECT 1560.880 1671.450 1561.140 1671.770 ;
        RECT 1563.180 1671.450 1563.440 1671.770 ;
        RECT 1560.940 63.910 1561.080 1671.450 ;
        RECT 1103.640 63.590 1103.900 63.910 ;
        RECT 1560.880 63.590 1561.140 63.910 ;
        RECT 1103.700 3.050 1103.840 63.590 ;
        RECT 1102.720 2.730 1102.980 3.050 ;
        RECT 1103.640 2.730 1103.900 3.050 ;
        RECT 1102.780 2.400 1102.920 2.730 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1567.825 807.245 1567.995 855.355 ;
        RECT 1568.285 752.165 1568.455 753.015 ;
        RECT 1568.285 512.125 1568.455 565.675 ;
        RECT 1568.285 372.725 1568.455 420.835 ;
      LAYER mcon ;
        RECT 1567.825 855.185 1567.995 855.355 ;
        RECT 1568.285 752.845 1568.455 753.015 ;
        RECT 1568.285 565.505 1568.455 565.675 ;
        RECT 1568.285 420.665 1568.455 420.835 ;
      LAYER met1 ;
        RECT 1567.290 1531.940 1567.610 1532.000 ;
        RECT 1567.750 1531.940 1568.070 1532.000 ;
        RECT 1567.290 1531.800 1568.070 1531.940 ;
        RECT 1567.290 1531.740 1567.610 1531.800 ;
        RECT 1567.750 1531.740 1568.070 1531.800 ;
        RECT 1567.750 1007.320 1568.070 1007.380 ;
        RECT 1568.210 1007.320 1568.530 1007.380 ;
        RECT 1567.750 1007.180 1568.530 1007.320 ;
        RECT 1567.750 1007.120 1568.070 1007.180 ;
        RECT 1568.210 1007.120 1568.530 1007.180 ;
        RECT 1568.210 903.960 1568.530 904.020 ;
        RECT 1568.670 903.960 1568.990 904.020 ;
        RECT 1568.210 903.820 1568.990 903.960 ;
        RECT 1568.210 903.760 1568.530 903.820 ;
        RECT 1568.670 903.760 1568.990 903.820 ;
        RECT 1567.750 855.340 1568.070 855.400 ;
        RECT 1567.555 855.200 1568.070 855.340 ;
        RECT 1567.750 855.140 1568.070 855.200 ;
        RECT 1567.765 807.400 1568.055 807.445 ;
        RECT 1569.130 807.400 1569.450 807.460 ;
        RECT 1567.765 807.260 1569.450 807.400 ;
        RECT 1567.765 807.215 1568.055 807.260 ;
        RECT 1569.130 807.200 1569.450 807.260 ;
        RECT 1568.225 753.000 1568.515 753.045 ;
        RECT 1569.130 753.000 1569.450 753.060 ;
        RECT 1568.225 752.860 1569.450 753.000 ;
        RECT 1568.225 752.815 1568.515 752.860 ;
        RECT 1569.130 752.800 1569.450 752.860 ;
        RECT 1568.210 752.320 1568.530 752.380 ;
        RECT 1568.015 752.180 1568.530 752.320 ;
        RECT 1568.210 752.120 1568.530 752.180 ;
        RECT 1568.210 565.660 1568.530 565.720 ;
        RECT 1568.015 565.520 1568.530 565.660 ;
        RECT 1568.210 565.460 1568.530 565.520 ;
        RECT 1567.290 512.280 1567.610 512.340 ;
        RECT 1568.225 512.280 1568.515 512.325 ;
        RECT 1567.290 512.140 1568.515 512.280 ;
        RECT 1567.290 512.080 1567.610 512.140 ;
        RECT 1568.225 512.095 1568.515 512.140 ;
        RECT 1567.290 427.960 1567.610 428.020 ;
        RECT 1568.210 427.960 1568.530 428.020 ;
        RECT 1567.290 427.820 1568.530 427.960 ;
        RECT 1567.290 427.760 1567.610 427.820 ;
        RECT 1568.210 427.760 1568.530 427.820 ;
        RECT 1568.210 420.820 1568.530 420.880 ;
        RECT 1568.015 420.680 1568.530 420.820 ;
        RECT 1568.210 420.620 1568.530 420.680 ;
        RECT 1568.225 372.880 1568.515 372.925 ;
        RECT 1568.670 372.880 1568.990 372.940 ;
        RECT 1568.225 372.740 1568.990 372.880 ;
        RECT 1568.225 372.695 1568.515 372.740 ;
        RECT 1568.670 372.680 1568.990 372.740 ;
        RECT 1568.670 283.260 1568.990 283.520 ;
        RECT 1568.760 282.840 1568.900 283.260 ;
        RECT 1568.670 282.580 1568.990 282.840 ;
        RECT 1567.750 207.300 1568.070 207.360 ;
        RECT 1568.670 207.300 1568.990 207.360 ;
        RECT 1567.750 207.160 1568.990 207.300 ;
        RECT 1567.750 207.100 1568.070 207.160 ;
        RECT 1568.670 207.100 1568.990 207.160 ;
        RECT 1124.310 63.480 1124.630 63.540 ;
        RECT 1567.750 63.480 1568.070 63.540 ;
        RECT 1124.310 63.340 1568.070 63.480 ;
        RECT 1124.310 63.280 1124.630 63.340 ;
        RECT 1567.750 63.280 1568.070 63.340 ;
        RECT 1120.630 2.960 1120.950 3.020 ;
        RECT 1124.310 2.960 1124.630 3.020 ;
        RECT 1120.630 2.820 1124.630 2.960 ;
        RECT 1120.630 2.760 1120.950 2.820 ;
        RECT 1124.310 2.760 1124.630 2.820 ;
      LAYER via ;
        RECT 1567.320 1531.740 1567.580 1532.000 ;
        RECT 1567.780 1531.740 1568.040 1532.000 ;
        RECT 1567.780 1007.120 1568.040 1007.380 ;
        RECT 1568.240 1007.120 1568.500 1007.380 ;
        RECT 1568.240 903.760 1568.500 904.020 ;
        RECT 1568.700 903.760 1568.960 904.020 ;
        RECT 1567.780 855.140 1568.040 855.400 ;
        RECT 1569.160 807.200 1569.420 807.460 ;
        RECT 1569.160 752.800 1569.420 753.060 ;
        RECT 1568.240 752.120 1568.500 752.380 ;
        RECT 1568.240 565.460 1568.500 565.720 ;
        RECT 1567.320 512.080 1567.580 512.340 ;
        RECT 1567.320 427.760 1567.580 428.020 ;
        RECT 1568.240 427.760 1568.500 428.020 ;
        RECT 1568.240 420.620 1568.500 420.880 ;
        RECT 1568.700 372.680 1568.960 372.940 ;
        RECT 1568.700 283.260 1568.960 283.520 ;
        RECT 1568.700 282.580 1568.960 282.840 ;
        RECT 1567.780 207.100 1568.040 207.360 ;
        RECT 1568.700 207.100 1568.960 207.360 ;
        RECT 1124.340 63.280 1124.600 63.540 ;
        RECT 1567.780 63.280 1568.040 63.540 ;
        RECT 1120.660 2.760 1120.920 3.020 ;
        RECT 1124.340 2.760 1124.600 3.020 ;
      LAYER met2 ;
        RECT 1571.845 1700.410 1572.125 1704.000 ;
        RECT 1570.140 1700.270 1572.125 1700.410 ;
        RECT 1570.140 1642.725 1570.280 1700.270 ;
        RECT 1571.845 1700.000 1572.125 1700.270 ;
        RECT 1570.070 1642.355 1570.350 1642.725 ;
        RECT 1568.690 1641.675 1568.970 1642.045 ;
        RECT 1568.760 1611.330 1568.900 1641.675 ;
        RECT 1568.300 1611.190 1568.900 1611.330 ;
        RECT 1568.300 1580.165 1568.440 1611.190 ;
        RECT 1567.310 1579.795 1567.590 1580.165 ;
        RECT 1568.230 1579.795 1568.510 1580.165 ;
        RECT 1567.380 1532.030 1567.520 1579.795 ;
        RECT 1567.320 1531.710 1567.580 1532.030 ;
        RECT 1567.780 1531.710 1568.040 1532.030 ;
        RECT 1567.840 1442.690 1567.980 1531.710 ;
        RECT 1567.840 1442.550 1568.440 1442.690 ;
        RECT 1568.300 1007.410 1568.440 1442.550 ;
        RECT 1567.780 1007.090 1568.040 1007.410 ;
        RECT 1568.240 1007.090 1568.500 1007.410 ;
        RECT 1567.840 952.410 1567.980 1007.090 ;
        RECT 1567.840 952.270 1568.440 952.410 ;
        RECT 1568.300 904.050 1568.440 952.270 ;
        RECT 1568.240 903.730 1568.500 904.050 ;
        RECT 1568.700 903.730 1568.960 904.050 ;
        RECT 1568.760 855.850 1568.900 903.730 ;
        RECT 1567.840 855.710 1568.900 855.850 ;
        RECT 1567.840 855.430 1567.980 855.710 ;
        RECT 1567.780 855.110 1568.040 855.430 ;
        RECT 1569.160 807.170 1569.420 807.490 ;
        RECT 1569.220 753.090 1569.360 807.170 ;
        RECT 1569.160 752.770 1569.420 753.090 ;
        RECT 1568.240 752.090 1568.500 752.410 ;
        RECT 1568.300 565.750 1568.440 752.090 ;
        RECT 1568.240 565.430 1568.500 565.750 ;
        RECT 1567.320 512.050 1567.580 512.370 ;
        RECT 1567.380 428.050 1567.520 512.050 ;
        RECT 1567.320 427.730 1567.580 428.050 ;
        RECT 1568.240 427.730 1568.500 428.050 ;
        RECT 1568.300 420.910 1568.440 427.730 ;
        RECT 1568.240 420.590 1568.500 420.910 ;
        RECT 1568.700 372.650 1568.960 372.970 ;
        RECT 1568.760 283.550 1568.900 372.650 ;
        RECT 1568.700 283.230 1568.960 283.550 ;
        RECT 1568.700 282.550 1568.960 282.870 ;
        RECT 1568.760 207.390 1568.900 282.550 ;
        RECT 1567.780 207.070 1568.040 207.390 ;
        RECT 1568.700 207.070 1568.960 207.390 ;
        RECT 1567.840 63.570 1567.980 207.070 ;
        RECT 1124.340 63.250 1124.600 63.570 ;
        RECT 1567.780 63.250 1568.040 63.570 ;
        RECT 1124.400 3.050 1124.540 63.250 ;
        RECT 1120.660 2.730 1120.920 3.050 ;
        RECT 1124.340 2.730 1124.600 3.050 ;
        RECT 1120.720 2.400 1120.860 2.730 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
      LAYER via2 ;
        RECT 1570.070 1642.400 1570.350 1642.680 ;
        RECT 1568.690 1641.720 1568.970 1642.000 ;
        RECT 1567.310 1579.840 1567.590 1580.120 ;
        RECT 1568.230 1579.840 1568.510 1580.120 ;
      LAYER met3 ;
        RECT 1570.045 1642.690 1570.375 1642.705 ;
        RECT 1567.990 1642.390 1570.375 1642.690 ;
        RECT 1567.990 1642.010 1568.290 1642.390 ;
        RECT 1570.045 1642.375 1570.375 1642.390 ;
        RECT 1568.665 1642.010 1568.995 1642.025 ;
        RECT 1567.990 1641.710 1568.995 1642.010 ;
        RECT 1568.665 1641.695 1568.995 1641.710 ;
        RECT 1567.285 1580.130 1567.615 1580.145 ;
        RECT 1568.205 1580.130 1568.535 1580.145 ;
        RECT 1567.285 1579.830 1568.535 1580.130 ;
        RECT 1567.285 1579.815 1567.615 1579.830 ;
        RECT 1568.205 1579.815 1568.535 1579.830 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1574.650 1651.280 1574.970 1651.340 ;
        RECT 1576.950 1651.280 1577.270 1651.340 ;
        RECT 1574.650 1651.140 1577.270 1651.280 ;
        RECT 1574.650 1651.080 1574.970 1651.140 ;
        RECT 1576.950 1651.080 1577.270 1651.140 ;
        RECT 1145.010 63.140 1145.330 63.200 ;
        RECT 1574.650 63.140 1574.970 63.200 ;
        RECT 1145.010 63.000 1574.970 63.140 ;
        RECT 1145.010 62.940 1145.330 63.000 ;
        RECT 1574.650 62.940 1574.970 63.000 ;
        RECT 1138.570 37.980 1138.890 38.040 ;
        RECT 1145.010 37.980 1145.330 38.040 ;
        RECT 1138.570 37.840 1145.330 37.980 ;
        RECT 1138.570 37.780 1138.890 37.840 ;
        RECT 1145.010 37.780 1145.330 37.840 ;
      LAYER via ;
        RECT 1574.680 1651.080 1574.940 1651.340 ;
        RECT 1576.980 1651.080 1577.240 1651.340 ;
        RECT 1145.040 62.940 1145.300 63.200 ;
        RECT 1574.680 62.940 1574.940 63.200 ;
        RECT 1138.600 37.780 1138.860 38.040 ;
        RECT 1145.040 37.780 1145.300 38.040 ;
      LAYER met2 ;
        RECT 1578.745 1700.410 1579.025 1704.000 ;
        RECT 1577.040 1700.270 1579.025 1700.410 ;
        RECT 1577.040 1651.370 1577.180 1700.270 ;
        RECT 1578.745 1700.000 1579.025 1700.270 ;
        RECT 1574.680 1651.050 1574.940 1651.370 ;
        RECT 1576.980 1651.050 1577.240 1651.370 ;
        RECT 1574.740 63.230 1574.880 1651.050 ;
        RECT 1145.040 62.910 1145.300 63.230 ;
        RECT 1574.680 62.910 1574.940 63.230 ;
        RECT 1145.100 38.070 1145.240 62.910 ;
        RECT 1138.600 37.750 1138.860 38.070 ;
        RECT 1145.040 37.750 1145.300 38.070 ;
        RECT 1138.660 2.400 1138.800 37.750 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1581.625 1490.645 1581.795 1538.755 ;
        RECT 1581.165 1435.225 1581.335 1442.535 ;
        RECT 1581.165 952.425 1581.335 959.395 ;
        RECT 1581.625 662.405 1581.795 710.515 ;
        RECT 1156.585 48.365 1156.755 62.815 ;
      LAYER mcon ;
        RECT 1581.625 1538.585 1581.795 1538.755 ;
        RECT 1581.165 1442.365 1581.335 1442.535 ;
        RECT 1581.165 959.225 1581.335 959.395 ;
        RECT 1581.625 710.345 1581.795 710.515 ;
        RECT 1156.585 62.645 1156.755 62.815 ;
      LAYER met1 ;
        RECT 1582.010 1642.440 1582.330 1642.500 ;
        RECT 1582.930 1642.440 1583.250 1642.500 ;
        RECT 1582.010 1642.300 1583.250 1642.440 ;
        RECT 1582.010 1642.240 1582.330 1642.300 ;
        RECT 1582.930 1642.240 1583.250 1642.300 ;
        RECT 1582.010 1594.500 1582.330 1594.560 ;
        RECT 1581.640 1594.360 1582.330 1594.500 ;
        RECT 1581.640 1593.880 1581.780 1594.360 ;
        RECT 1582.010 1594.300 1582.330 1594.360 ;
        RECT 1581.550 1593.620 1581.870 1593.880 ;
        RECT 1581.550 1538.740 1581.870 1538.800 ;
        RECT 1581.355 1538.600 1581.870 1538.740 ;
        RECT 1581.550 1538.540 1581.870 1538.600 ;
        RECT 1581.550 1490.800 1581.870 1490.860 ;
        RECT 1581.355 1490.660 1581.870 1490.800 ;
        RECT 1581.550 1490.600 1581.870 1490.660 ;
        RECT 1581.105 1442.520 1581.395 1442.565 ;
        RECT 1581.550 1442.520 1581.870 1442.580 ;
        RECT 1581.105 1442.380 1581.870 1442.520 ;
        RECT 1581.105 1442.335 1581.395 1442.380 ;
        RECT 1581.550 1442.320 1581.870 1442.380 ;
        RECT 1581.090 1435.380 1581.410 1435.440 ;
        RECT 1580.895 1435.240 1581.410 1435.380 ;
        RECT 1581.090 1435.180 1581.410 1435.240 ;
        RECT 1581.090 1393.900 1581.410 1393.960 ;
        RECT 1581.550 1393.900 1581.870 1393.960 ;
        RECT 1581.090 1393.760 1581.870 1393.900 ;
        RECT 1581.090 1393.700 1581.410 1393.760 ;
        RECT 1581.550 1393.700 1581.870 1393.760 ;
        RECT 1581.090 1104.220 1581.410 1104.280 ;
        RECT 1581.550 1104.220 1581.870 1104.280 ;
        RECT 1581.090 1104.080 1581.870 1104.220 ;
        RECT 1581.090 1104.020 1581.410 1104.080 ;
        RECT 1581.550 1104.020 1581.870 1104.080 ;
        RECT 1581.550 1055.600 1581.870 1055.660 ;
        RECT 1582.470 1055.600 1582.790 1055.660 ;
        RECT 1581.550 1055.460 1582.790 1055.600 ;
        RECT 1581.550 1055.400 1581.870 1055.460 ;
        RECT 1582.470 1055.400 1582.790 1055.460 ;
        RECT 1581.105 959.380 1581.395 959.425 ;
        RECT 1581.550 959.380 1581.870 959.440 ;
        RECT 1581.105 959.240 1581.870 959.380 ;
        RECT 1581.105 959.195 1581.395 959.240 ;
        RECT 1581.550 959.180 1581.870 959.240 ;
        RECT 1581.090 952.580 1581.410 952.640 ;
        RECT 1580.895 952.440 1581.410 952.580 ;
        RECT 1581.090 952.380 1581.410 952.440 ;
        RECT 1581.090 911.100 1581.410 911.160 ;
        RECT 1581.550 911.100 1581.870 911.160 ;
        RECT 1581.090 910.960 1581.870 911.100 ;
        RECT 1581.090 910.900 1581.410 910.960 ;
        RECT 1581.550 910.900 1581.870 910.960 ;
        RECT 1581.550 772.720 1581.870 772.780 ;
        RECT 1582.010 772.720 1582.330 772.780 ;
        RECT 1581.550 772.580 1582.330 772.720 ;
        RECT 1581.550 772.520 1581.870 772.580 ;
        RECT 1582.010 772.520 1582.330 772.580 ;
        RECT 1581.550 710.500 1581.870 710.560 ;
        RECT 1581.355 710.360 1581.870 710.500 ;
        RECT 1581.550 710.300 1581.870 710.360 ;
        RECT 1581.550 662.560 1581.870 662.620 ;
        RECT 1581.355 662.420 1581.870 662.560 ;
        RECT 1581.550 662.360 1581.870 662.420 ;
        RECT 1581.550 621.420 1581.870 621.480 ;
        RECT 1581.180 621.280 1581.870 621.420 ;
        RECT 1581.180 621.140 1581.320 621.280 ;
        RECT 1581.550 621.220 1581.870 621.280 ;
        RECT 1581.090 620.880 1581.410 621.140 ;
        RECT 1581.090 572.800 1581.410 572.860 ;
        RECT 1581.550 572.800 1581.870 572.860 ;
        RECT 1581.090 572.660 1581.870 572.800 ;
        RECT 1581.090 572.600 1581.410 572.660 ;
        RECT 1581.550 572.600 1581.870 572.660 ;
        RECT 1156.525 62.800 1156.815 62.845 ;
        RECT 1581.090 62.800 1581.410 62.860 ;
        RECT 1156.525 62.660 1581.410 62.800 ;
        RECT 1156.525 62.615 1156.815 62.660 ;
        RECT 1581.090 62.600 1581.410 62.660 ;
        RECT 1156.510 48.520 1156.830 48.580 ;
        RECT 1156.315 48.380 1156.830 48.520 ;
        RECT 1156.510 48.320 1156.830 48.380 ;
      LAYER via ;
        RECT 1582.040 1642.240 1582.300 1642.500 ;
        RECT 1582.960 1642.240 1583.220 1642.500 ;
        RECT 1582.040 1594.300 1582.300 1594.560 ;
        RECT 1581.580 1593.620 1581.840 1593.880 ;
        RECT 1581.580 1538.540 1581.840 1538.800 ;
        RECT 1581.580 1490.600 1581.840 1490.860 ;
        RECT 1581.580 1442.320 1581.840 1442.580 ;
        RECT 1581.120 1435.180 1581.380 1435.440 ;
        RECT 1581.120 1393.700 1581.380 1393.960 ;
        RECT 1581.580 1393.700 1581.840 1393.960 ;
        RECT 1581.120 1104.020 1581.380 1104.280 ;
        RECT 1581.580 1104.020 1581.840 1104.280 ;
        RECT 1581.580 1055.400 1581.840 1055.660 ;
        RECT 1582.500 1055.400 1582.760 1055.660 ;
        RECT 1581.580 959.180 1581.840 959.440 ;
        RECT 1581.120 952.380 1581.380 952.640 ;
        RECT 1581.120 910.900 1581.380 911.160 ;
        RECT 1581.580 910.900 1581.840 911.160 ;
        RECT 1581.580 772.520 1581.840 772.780 ;
        RECT 1582.040 772.520 1582.300 772.780 ;
        RECT 1581.580 710.300 1581.840 710.560 ;
        RECT 1581.580 662.360 1581.840 662.620 ;
        RECT 1581.580 621.220 1581.840 621.480 ;
        RECT 1581.120 620.880 1581.380 621.140 ;
        RECT 1581.120 572.600 1581.380 572.860 ;
        RECT 1581.580 572.600 1581.840 572.860 ;
        RECT 1581.120 62.600 1581.380 62.860 ;
        RECT 1156.540 48.320 1156.800 48.580 ;
      LAYER met2 ;
        RECT 1585.185 1700.410 1585.465 1704.000 ;
        RECT 1583.480 1700.270 1585.465 1700.410 ;
        RECT 1583.480 1667.090 1583.620 1700.270 ;
        RECT 1585.185 1700.000 1585.465 1700.270 ;
        RECT 1583.020 1666.950 1583.620 1667.090 ;
        RECT 1583.020 1642.530 1583.160 1666.950 ;
        RECT 1582.040 1642.210 1582.300 1642.530 ;
        RECT 1582.960 1642.210 1583.220 1642.530 ;
        RECT 1582.100 1594.590 1582.240 1642.210 ;
        RECT 1582.040 1594.270 1582.300 1594.590 ;
        RECT 1581.580 1593.590 1581.840 1593.910 ;
        RECT 1581.640 1538.830 1581.780 1593.590 ;
        RECT 1581.580 1538.510 1581.840 1538.830 ;
        RECT 1581.580 1490.570 1581.840 1490.890 ;
        RECT 1581.640 1442.610 1581.780 1490.570 ;
        RECT 1581.580 1442.290 1581.840 1442.610 ;
        RECT 1581.120 1435.150 1581.380 1435.470 ;
        RECT 1581.180 1393.990 1581.320 1435.150 ;
        RECT 1581.120 1393.670 1581.380 1393.990 ;
        RECT 1581.580 1393.670 1581.840 1393.990 ;
        RECT 1581.640 1152.330 1581.780 1393.670 ;
        RECT 1581.180 1152.190 1581.780 1152.330 ;
        RECT 1581.180 1104.310 1581.320 1152.190 ;
        RECT 1581.120 1103.990 1581.380 1104.310 ;
        RECT 1581.580 1103.990 1581.840 1104.310 ;
        RECT 1581.640 1055.690 1581.780 1103.990 ;
        RECT 1581.580 1055.370 1581.840 1055.690 ;
        RECT 1582.500 1055.370 1582.760 1055.690 ;
        RECT 1582.560 1007.605 1582.700 1055.370 ;
        RECT 1581.570 1007.235 1581.850 1007.605 ;
        RECT 1582.490 1007.235 1582.770 1007.605 ;
        RECT 1581.640 959.470 1581.780 1007.235 ;
        RECT 1581.580 959.150 1581.840 959.470 ;
        RECT 1581.120 952.350 1581.380 952.670 ;
        RECT 1581.180 911.190 1581.320 952.350 ;
        RECT 1581.120 910.870 1581.380 911.190 ;
        RECT 1581.580 910.870 1581.840 911.190 ;
        RECT 1581.640 772.810 1581.780 910.870 ;
        RECT 1581.580 772.490 1581.840 772.810 ;
        RECT 1582.040 772.490 1582.300 772.810 ;
        RECT 1582.100 717.810 1582.240 772.490 ;
        RECT 1581.640 717.670 1582.240 717.810 ;
        RECT 1581.640 710.590 1581.780 717.670 ;
        RECT 1581.580 710.270 1581.840 710.590 ;
        RECT 1581.580 662.330 1581.840 662.650 ;
        RECT 1581.640 621.510 1581.780 662.330 ;
        RECT 1581.580 621.190 1581.840 621.510 ;
        RECT 1581.120 620.850 1581.380 621.170 ;
        RECT 1581.180 572.890 1581.320 620.850 ;
        RECT 1581.120 572.570 1581.380 572.890 ;
        RECT 1581.580 572.570 1581.840 572.890 ;
        RECT 1581.640 103.090 1581.780 572.570 ;
        RECT 1581.180 102.950 1581.780 103.090 ;
        RECT 1581.180 62.890 1581.320 102.950 ;
        RECT 1581.120 62.570 1581.380 62.890 ;
        RECT 1156.540 48.290 1156.800 48.610 ;
        RECT 1156.600 2.400 1156.740 48.290 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
      LAYER via2 ;
        RECT 1581.570 1007.280 1581.850 1007.560 ;
        RECT 1582.490 1007.280 1582.770 1007.560 ;
      LAYER met3 ;
        RECT 1581.545 1007.570 1581.875 1007.585 ;
        RECT 1582.465 1007.570 1582.795 1007.585 ;
        RECT 1581.545 1007.270 1582.795 1007.570 ;
        RECT 1581.545 1007.255 1581.875 1007.270 ;
        RECT 1582.465 1007.255 1582.795 1007.270 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 675.810 66.200 676.130 66.260 ;
        RECT 1401.690 66.200 1402.010 66.260 ;
        RECT 675.810 66.060 1402.010 66.200 ;
        RECT 675.810 66.000 676.130 66.060 ;
        RECT 1401.690 66.000 1402.010 66.060 ;
      LAYER via ;
        RECT 675.840 66.000 676.100 66.260 ;
        RECT 1401.720 66.000 1401.980 66.260 ;
      LAYER met2 ;
        RECT 1403.485 1700.410 1403.765 1704.000 ;
        RECT 1401.780 1700.270 1403.765 1700.410 ;
        RECT 1401.780 66.290 1401.920 1700.270 ;
        RECT 1403.485 1700.000 1403.765 1700.270 ;
        RECT 675.840 65.970 676.100 66.290 ;
        RECT 1401.720 65.970 1401.980 66.290 ;
        RECT 675.900 3.130 676.040 65.970 ;
        RECT 674.520 2.990 676.040 3.130 ;
        RECT 674.520 2.400 674.660 2.990 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1589.370 1594.500 1589.690 1594.560 ;
        RECT 1589.000 1594.360 1589.690 1594.500 ;
        RECT 1589.000 1594.220 1589.140 1594.360 ;
        RECT 1589.370 1594.300 1589.690 1594.360 ;
        RECT 1588.910 1593.960 1589.230 1594.220 ;
        RECT 1173.990 37.980 1174.310 38.040 ;
        RECT 1588.910 37.980 1589.230 38.040 ;
        RECT 1173.990 37.840 1589.230 37.980 ;
        RECT 1173.990 37.780 1174.310 37.840 ;
        RECT 1588.910 37.780 1589.230 37.840 ;
      LAYER via ;
        RECT 1589.400 1594.300 1589.660 1594.560 ;
        RECT 1588.940 1593.960 1589.200 1594.220 ;
        RECT 1174.020 37.780 1174.280 38.040 ;
        RECT 1588.940 37.780 1589.200 38.040 ;
      LAYER met2 ;
        RECT 1592.085 1700.410 1592.365 1704.000 ;
        RECT 1590.380 1700.270 1592.365 1700.410 ;
        RECT 1590.380 1642.610 1590.520 1700.270 ;
        RECT 1592.085 1700.000 1592.365 1700.270 ;
        RECT 1589.460 1642.470 1590.520 1642.610 ;
        RECT 1589.460 1594.590 1589.600 1642.470 ;
        RECT 1589.400 1594.270 1589.660 1594.590 ;
        RECT 1588.940 1593.930 1589.200 1594.250 ;
        RECT 1589.000 38.070 1589.140 1593.930 ;
        RECT 1174.020 37.750 1174.280 38.070 ;
        RECT 1588.940 37.750 1589.200 38.070 ;
        RECT 1174.080 2.400 1174.220 37.750 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1595.885 1642.285 1596.055 1671.015 ;
      LAYER mcon ;
        RECT 1595.885 1670.845 1596.055 1671.015 ;
      LAYER met1 ;
        RECT 1595.825 1671.000 1596.115 1671.045 ;
        RECT 1597.190 1671.000 1597.510 1671.060 ;
        RECT 1595.825 1670.860 1597.510 1671.000 ;
        RECT 1595.825 1670.815 1596.115 1670.860 ;
        RECT 1597.190 1670.800 1597.510 1670.860 ;
        RECT 1595.810 1642.440 1596.130 1642.500 ;
        RECT 1595.615 1642.300 1596.130 1642.440 ;
        RECT 1595.810 1642.240 1596.130 1642.300 ;
        RECT 1191.930 38.320 1192.250 38.380 ;
        RECT 1595.810 38.320 1596.130 38.380 ;
        RECT 1191.930 38.180 1596.130 38.320 ;
        RECT 1191.930 38.120 1192.250 38.180 ;
        RECT 1595.810 38.120 1596.130 38.180 ;
      LAYER via ;
        RECT 1597.220 1670.800 1597.480 1671.060 ;
        RECT 1595.840 1642.240 1596.100 1642.500 ;
        RECT 1191.960 38.120 1192.220 38.380 ;
        RECT 1595.840 38.120 1596.100 38.380 ;
      LAYER met2 ;
        RECT 1598.525 1700.410 1598.805 1704.000 ;
        RECT 1597.280 1700.270 1598.805 1700.410 ;
        RECT 1597.280 1671.090 1597.420 1700.270 ;
        RECT 1598.525 1700.000 1598.805 1700.270 ;
        RECT 1597.220 1670.770 1597.480 1671.090 ;
        RECT 1595.840 1642.210 1596.100 1642.530 ;
        RECT 1595.900 38.410 1596.040 1642.210 ;
        RECT 1191.960 38.090 1192.220 38.410 ;
        RECT 1595.840 38.090 1596.100 38.410 ;
        RECT 1192.020 2.400 1192.160 38.090 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1601.330 1678.140 1601.650 1678.200 ;
        RECT 1603.630 1678.140 1603.950 1678.200 ;
        RECT 1601.330 1678.000 1603.950 1678.140 ;
        RECT 1601.330 1677.940 1601.650 1678.000 ;
        RECT 1603.630 1677.940 1603.950 1678.000 ;
        RECT 1209.870 38.660 1210.190 38.720 ;
        RECT 1601.330 38.660 1601.650 38.720 ;
        RECT 1209.870 38.520 1601.650 38.660 ;
        RECT 1209.870 38.460 1210.190 38.520 ;
        RECT 1601.330 38.460 1601.650 38.520 ;
      LAYER via ;
        RECT 1601.360 1677.940 1601.620 1678.200 ;
        RECT 1603.660 1677.940 1603.920 1678.200 ;
        RECT 1209.900 38.460 1210.160 38.720 ;
        RECT 1601.360 38.460 1601.620 38.720 ;
      LAYER met2 ;
        RECT 1605.425 1700.410 1605.705 1704.000 ;
        RECT 1603.720 1700.270 1605.705 1700.410 ;
        RECT 1603.720 1678.230 1603.860 1700.270 ;
        RECT 1605.425 1700.000 1605.705 1700.270 ;
        RECT 1601.360 1677.910 1601.620 1678.230 ;
        RECT 1603.660 1677.910 1603.920 1678.230 ;
        RECT 1601.420 38.750 1601.560 1677.910 ;
        RECT 1209.900 38.430 1210.160 38.750 ;
        RECT 1601.360 38.430 1601.620 38.750 ;
        RECT 1209.960 2.400 1210.100 38.430 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1608.230 1678.140 1608.550 1678.200 ;
        RECT 1610.990 1678.140 1611.310 1678.200 ;
        RECT 1608.230 1678.000 1611.310 1678.140 ;
        RECT 1608.230 1677.940 1608.550 1678.000 ;
        RECT 1610.990 1677.940 1611.310 1678.000 ;
        RECT 1227.810 39.000 1228.130 39.060 ;
        RECT 1608.230 39.000 1608.550 39.060 ;
        RECT 1227.810 38.860 1608.550 39.000 ;
        RECT 1227.810 38.800 1228.130 38.860 ;
        RECT 1608.230 38.800 1608.550 38.860 ;
      LAYER via ;
        RECT 1608.260 1677.940 1608.520 1678.200 ;
        RECT 1611.020 1677.940 1611.280 1678.200 ;
        RECT 1227.840 38.800 1228.100 39.060 ;
        RECT 1608.260 38.800 1608.520 39.060 ;
      LAYER met2 ;
        RECT 1612.325 1700.410 1612.605 1704.000 ;
        RECT 1611.080 1700.270 1612.605 1700.410 ;
        RECT 1611.080 1678.230 1611.220 1700.270 ;
        RECT 1612.325 1700.000 1612.605 1700.270 ;
        RECT 1608.260 1677.910 1608.520 1678.230 ;
        RECT 1611.020 1677.910 1611.280 1678.230 ;
        RECT 1608.320 39.090 1608.460 1677.910 ;
        RECT 1227.840 38.770 1228.100 39.090 ;
        RECT 1608.260 38.770 1608.520 39.090 ;
        RECT 1227.900 2.400 1228.040 38.770 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1615.130 1678.480 1615.450 1678.540 ;
        RECT 1617.430 1678.480 1617.750 1678.540 ;
        RECT 1615.130 1678.340 1617.750 1678.480 ;
        RECT 1615.130 1678.280 1615.450 1678.340 ;
        RECT 1617.430 1678.280 1617.750 1678.340 ;
        RECT 1245.750 39.340 1246.070 39.400 ;
        RECT 1615.130 39.340 1615.450 39.400 ;
        RECT 1245.750 39.200 1615.450 39.340 ;
        RECT 1245.750 39.140 1246.070 39.200 ;
        RECT 1615.130 39.140 1615.450 39.200 ;
      LAYER via ;
        RECT 1615.160 1678.280 1615.420 1678.540 ;
        RECT 1617.460 1678.280 1617.720 1678.540 ;
        RECT 1245.780 39.140 1246.040 39.400 ;
        RECT 1615.160 39.140 1615.420 39.400 ;
      LAYER met2 ;
        RECT 1618.765 1700.410 1619.045 1704.000 ;
        RECT 1617.520 1700.270 1619.045 1700.410 ;
        RECT 1617.520 1678.570 1617.660 1700.270 ;
        RECT 1618.765 1700.000 1619.045 1700.270 ;
        RECT 1615.160 1678.250 1615.420 1678.570 ;
        RECT 1617.460 1678.250 1617.720 1678.570 ;
        RECT 1615.220 39.430 1615.360 1678.250 ;
        RECT 1245.780 39.110 1246.040 39.430 ;
        RECT 1615.160 39.110 1615.420 39.430 ;
        RECT 1245.840 2.400 1245.980 39.110 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1623.485 1641.605 1623.655 1683.595 ;
        RECT 1623.025 1449.505 1623.195 1497.275 ;
        RECT 1622.565 1317.245 1622.735 1393.575 ;
        RECT 1623.025 1256.045 1623.195 1304.155 ;
        RECT 1623.025 772.905 1623.195 821.015 ;
        RECT 1623.485 524.365 1623.655 531.675 ;
        RECT 1623.025 265.285 1623.195 331.075 ;
        RECT 1623.025 96.645 1623.195 144.755 ;
      LAYER mcon ;
        RECT 1623.485 1683.425 1623.655 1683.595 ;
        RECT 1623.025 1497.105 1623.195 1497.275 ;
        RECT 1622.565 1393.405 1622.735 1393.575 ;
        RECT 1623.025 1303.985 1623.195 1304.155 ;
        RECT 1623.025 820.845 1623.195 821.015 ;
        RECT 1623.485 531.505 1623.655 531.675 ;
        RECT 1623.025 330.905 1623.195 331.075 ;
        RECT 1623.025 144.585 1623.195 144.755 ;
      LAYER met1 ;
        RECT 1623.410 1683.580 1623.730 1683.640 ;
        RECT 1623.215 1683.440 1623.730 1683.580 ;
        RECT 1623.410 1683.380 1623.730 1683.440 ;
        RECT 1623.425 1641.760 1623.715 1641.805 ;
        RECT 1623.870 1641.760 1624.190 1641.820 ;
        RECT 1623.425 1641.620 1624.190 1641.760 ;
        RECT 1623.425 1641.575 1623.715 1641.620 ;
        RECT 1623.870 1641.560 1624.190 1641.620 ;
        RECT 1622.950 1593.480 1623.270 1593.540 ;
        RECT 1623.870 1593.480 1624.190 1593.540 ;
        RECT 1622.950 1593.340 1624.190 1593.480 ;
        RECT 1622.950 1593.280 1623.270 1593.340 ;
        RECT 1623.870 1593.280 1624.190 1593.340 ;
        RECT 1622.965 1497.260 1623.255 1497.305 ;
        RECT 1623.410 1497.260 1623.730 1497.320 ;
        RECT 1622.965 1497.120 1623.730 1497.260 ;
        RECT 1622.965 1497.075 1623.255 1497.120 ;
        RECT 1623.410 1497.060 1623.730 1497.120 ;
        RECT 1622.950 1449.660 1623.270 1449.720 ;
        RECT 1622.755 1449.520 1623.270 1449.660 ;
        RECT 1622.950 1449.460 1623.270 1449.520 ;
        RECT 1622.950 1448.780 1623.270 1449.040 ;
        RECT 1623.040 1448.640 1623.180 1448.780 ;
        RECT 1623.870 1448.640 1624.190 1448.700 ;
        RECT 1623.040 1448.500 1624.190 1448.640 ;
        RECT 1623.870 1448.440 1624.190 1448.500 ;
        RECT 1622.490 1400.700 1622.810 1400.760 ;
        RECT 1623.870 1400.700 1624.190 1400.760 ;
        RECT 1622.490 1400.560 1624.190 1400.700 ;
        RECT 1622.490 1400.500 1622.810 1400.560 ;
        RECT 1623.870 1400.500 1624.190 1400.560 ;
        RECT 1622.490 1393.560 1622.810 1393.620 ;
        RECT 1622.295 1393.420 1622.810 1393.560 ;
        RECT 1622.490 1393.360 1622.810 1393.420 ;
        RECT 1622.505 1317.400 1622.795 1317.445 ;
        RECT 1623.410 1317.400 1623.730 1317.460 ;
        RECT 1622.505 1317.260 1623.730 1317.400 ;
        RECT 1622.505 1317.215 1622.795 1317.260 ;
        RECT 1623.410 1317.200 1623.730 1317.260 ;
        RECT 1622.965 1304.140 1623.255 1304.185 ;
        RECT 1623.410 1304.140 1623.730 1304.200 ;
        RECT 1622.965 1304.000 1623.730 1304.140 ;
        RECT 1622.965 1303.955 1623.255 1304.000 ;
        RECT 1623.410 1303.940 1623.730 1304.000 ;
        RECT 1622.950 1256.200 1623.270 1256.260 ;
        RECT 1622.755 1256.060 1623.270 1256.200 ;
        RECT 1622.950 1256.000 1623.270 1256.060 ;
        RECT 1623.870 1207.580 1624.190 1207.640 ;
        RECT 1624.330 1207.580 1624.650 1207.640 ;
        RECT 1623.870 1207.440 1624.650 1207.580 ;
        RECT 1623.870 1207.380 1624.190 1207.440 ;
        RECT 1624.330 1207.380 1624.650 1207.440 ;
        RECT 1622.950 1159.300 1623.270 1159.360 ;
        RECT 1624.330 1159.300 1624.650 1159.360 ;
        RECT 1622.950 1159.160 1624.650 1159.300 ;
        RECT 1622.950 1159.100 1623.270 1159.160 ;
        RECT 1624.330 1159.100 1624.650 1159.160 ;
        RECT 1622.950 1062.740 1623.270 1062.800 ;
        RECT 1624.330 1062.740 1624.650 1062.800 ;
        RECT 1622.950 1062.600 1624.650 1062.740 ;
        RECT 1622.950 1062.540 1623.270 1062.600 ;
        RECT 1624.330 1062.540 1624.650 1062.600 ;
        RECT 1622.950 966.180 1623.270 966.240 ;
        RECT 1623.410 966.180 1623.730 966.240 ;
        RECT 1622.950 966.040 1623.730 966.180 ;
        RECT 1622.950 965.980 1623.270 966.040 ;
        RECT 1623.410 965.980 1623.730 966.040 ;
        RECT 1622.490 910.760 1622.810 910.820 ;
        RECT 1623.410 910.760 1623.730 910.820 ;
        RECT 1622.490 910.620 1623.730 910.760 ;
        RECT 1622.490 910.560 1622.810 910.620 ;
        RECT 1623.410 910.560 1623.730 910.620 ;
        RECT 1622.965 821.000 1623.255 821.045 ;
        RECT 1623.410 821.000 1623.730 821.060 ;
        RECT 1622.965 820.860 1623.730 821.000 ;
        RECT 1622.965 820.815 1623.255 820.860 ;
        RECT 1623.410 820.800 1623.730 820.860 ;
        RECT 1622.950 773.060 1623.270 773.120 ;
        RECT 1622.755 772.920 1623.270 773.060 ;
        RECT 1622.950 772.860 1623.270 772.920 ;
        RECT 1622.950 738.520 1623.270 738.780 ;
        RECT 1623.040 738.100 1623.180 738.520 ;
        RECT 1622.950 737.840 1623.270 738.100 ;
        RECT 1622.950 655.420 1623.270 655.480 ;
        RECT 1624.330 655.420 1624.650 655.480 ;
        RECT 1622.950 655.280 1624.650 655.420 ;
        RECT 1622.950 655.220 1623.270 655.280 ;
        RECT 1624.330 655.220 1624.650 655.280 ;
        RECT 1623.410 531.660 1623.730 531.720 ;
        RECT 1623.215 531.520 1623.730 531.660 ;
        RECT 1623.410 531.460 1623.730 531.520 ;
        RECT 1623.410 524.520 1623.730 524.580 ;
        RECT 1623.215 524.380 1623.730 524.520 ;
        RECT 1623.410 524.320 1623.730 524.380 ;
        RECT 1623.410 497.320 1623.730 497.380 ;
        RECT 1623.040 497.180 1623.730 497.320 ;
        RECT 1623.040 496.700 1623.180 497.180 ;
        RECT 1623.410 497.120 1623.730 497.180 ;
        RECT 1622.950 496.440 1623.270 496.700 ;
        RECT 1622.950 411.780 1623.270 412.040 ;
        RECT 1623.040 411.360 1623.180 411.780 ;
        RECT 1622.950 411.100 1623.270 411.360 ;
        RECT 1622.950 338.680 1623.270 338.940 ;
        RECT 1623.040 338.260 1623.180 338.680 ;
        RECT 1622.950 338.000 1623.270 338.260 ;
        RECT 1622.950 331.060 1623.270 331.120 ;
        RECT 1622.755 330.920 1623.270 331.060 ;
        RECT 1622.950 330.860 1623.270 330.920 ;
        RECT 1622.965 265.440 1623.255 265.485 ;
        RECT 1623.870 265.440 1624.190 265.500 ;
        RECT 1622.965 265.300 1624.190 265.440 ;
        RECT 1622.965 265.255 1623.255 265.300 ;
        RECT 1623.870 265.240 1624.190 265.300 ;
        RECT 1623.870 192.820 1624.190 193.080 ;
        RECT 1623.960 192.400 1624.100 192.820 ;
        RECT 1623.870 192.140 1624.190 192.400 ;
        RECT 1622.950 144.740 1623.270 144.800 ;
        RECT 1622.755 144.600 1623.270 144.740 ;
        RECT 1622.950 144.540 1623.270 144.600 ;
        RECT 1622.950 96.800 1623.270 96.860 ;
        RECT 1622.755 96.660 1623.270 96.800 ;
        RECT 1622.950 96.600 1623.270 96.660 ;
        RECT 1263.230 39.680 1263.550 39.740 ;
        RECT 1622.950 39.680 1623.270 39.740 ;
        RECT 1263.230 39.540 1623.270 39.680 ;
        RECT 1263.230 39.480 1263.550 39.540 ;
        RECT 1622.950 39.480 1623.270 39.540 ;
      LAYER via ;
        RECT 1623.440 1683.380 1623.700 1683.640 ;
        RECT 1623.900 1641.560 1624.160 1641.820 ;
        RECT 1622.980 1593.280 1623.240 1593.540 ;
        RECT 1623.900 1593.280 1624.160 1593.540 ;
        RECT 1623.440 1497.060 1623.700 1497.320 ;
        RECT 1622.980 1449.460 1623.240 1449.720 ;
        RECT 1622.980 1448.780 1623.240 1449.040 ;
        RECT 1623.900 1448.440 1624.160 1448.700 ;
        RECT 1622.520 1400.500 1622.780 1400.760 ;
        RECT 1623.900 1400.500 1624.160 1400.760 ;
        RECT 1622.520 1393.360 1622.780 1393.620 ;
        RECT 1623.440 1317.200 1623.700 1317.460 ;
        RECT 1623.440 1303.940 1623.700 1304.200 ;
        RECT 1622.980 1256.000 1623.240 1256.260 ;
        RECT 1623.900 1207.380 1624.160 1207.640 ;
        RECT 1624.360 1207.380 1624.620 1207.640 ;
        RECT 1622.980 1159.100 1623.240 1159.360 ;
        RECT 1624.360 1159.100 1624.620 1159.360 ;
        RECT 1622.980 1062.540 1623.240 1062.800 ;
        RECT 1624.360 1062.540 1624.620 1062.800 ;
        RECT 1622.980 965.980 1623.240 966.240 ;
        RECT 1623.440 965.980 1623.700 966.240 ;
        RECT 1622.520 910.560 1622.780 910.820 ;
        RECT 1623.440 910.560 1623.700 910.820 ;
        RECT 1623.440 820.800 1623.700 821.060 ;
        RECT 1622.980 772.860 1623.240 773.120 ;
        RECT 1622.980 738.520 1623.240 738.780 ;
        RECT 1622.980 737.840 1623.240 738.100 ;
        RECT 1622.980 655.220 1623.240 655.480 ;
        RECT 1624.360 655.220 1624.620 655.480 ;
        RECT 1623.440 531.460 1623.700 531.720 ;
        RECT 1623.440 524.320 1623.700 524.580 ;
        RECT 1623.440 497.120 1623.700 497.380 ;
        RECT 1622.980 496.440 1623.240 496.700 ;
        RECT 1622.980 411.780 1623.240 412.040 ;
        RECT 1622.980 411.100 1623.240 411.360 ;
        RECT 1622.980 338.680 1623.240 338.940 ;
        RECT 1622.980 338.000 1623.240 338.260 ;
        RECT 1622.980 330.860 1623.240 331.120 ;
        RECT 1623.900 265.240 1624.160 265.500 ;
        RECT 1623.900 192.820 1624.160 193.080 ;
        RECT 1623.900 192.140 1624.160 192.400 ;
        RECT 1622.980 144.540 1623.240 144.800 ;
        RECT 1622.980 96.600 1623.240 96.860 ;
        RECT 1263.260 39.480 1263.520 39.740 ;
        RECT 1622.980 39.480 1623.240 39.740 ;
      LAYER met2 ;
        RECT 1625.665 1700.000 1625.945 1704.000 ;
        RECT 1625.800 1691.685 1625.940 1700.000 ;
        RECT 1625.730 1691.315 1626.010 1691.685 ;
        RECT 1622.970 1690.890 1623.250 1691.005 ;
        RECT 1622.970 1690.750 1623.640 1690.890 ;
        RECT 1622.970 1690.635 1623.250 1690.750 ;
        RECT 1623.500 1683.670 1623.640 1690.750 ;
        RECT 1623.440 1683.350 1623.700 1683.670 ;
        RECT 1623.900 1641.530 1624.160 1641.850 ;
        RECT 1623.960 1607.250 1624.100 1641.530 ;
        RECT 1623.040 1607.110 1624.100 1607.250 ;
        RECT 1623.040 1593.570 1623.180 1607.110 ;
        RECT 1622.980 1593.250 1623.240 1593.570 ;
        RECT 1623.900 1593.250 1624.160 1593.570 ;
        RECT 1623.960 1558.970 1624.100 1593.250 ;
        RECT 1623.500 1558.830 1624.100 1558.970 ;
        RECT 1623.500 1497.350 1623.640 1558.830 ;
        RECT 1623.440 1497.030 1623.700 1497.350 ;
        RECT 1622.980 1449.430 1623.240 1449.750 ;
        RECT 1623.040 1449.070 1623.180 1449.430 ;
        RECT 1622.980 1448.750 1623.240 1449.070 ;
        RECT 1623.900 1448.410 1624.160 1448.730 ;
        RECT 1623.960 1400.790 1624.100 1448.410 ;
        RECT 1622.520 1400.470 1622.780 1400.790 ;
        RECT 1623.900 1400.470 1624.160 1400.790 ;
        RECT 1622.580 1393.650 1622.720 1400.470 ;
        RECT 1622.520 1393.330 1622.780 1393.650 ;
        RECT 1623.440 1317.170 1623.700 1317.490 ;
        RECT 1623.500 1304.230 1623.640 1317.170 ;
        RECT 1623.440 1303.910 1623.700 1304.230 ;
        RECT 1622.980 1255.970 1623.240 1256.290 ;
        RECT 1623.040 1255.805 1623.180 1255.970 ;
        RECT 1622.970 1255.435 1623.250 1255.805 ;
        RECT 1623.890 1255.435 1624.170 1255.805 ;
        RECT 1623.960 1207.670 1624.100 1255.435 ;
        RECT 1623.900 1207.350 1624.160 1207.670 ;
        RECT 1624.360 1207.350 1624.620 1207.670 ;
        RECT 1624.420 1159.390 1624.560 1207.350 ;
        RECT 1622.980 1159.245 1623.240 1159.390 ;
        RECT 1624.360 1159.245 1624.620 1159.390 ;
        RECT 1622.970 1158.875 1623.250 1159.245 ;
        RECT 1624.350 1158.875 1624.630 1159.245 ;
        RECT 1624.420 1062.830 1624.560 1158.875 ;
        RECT 1622.980 1062.510 1623.240 1062.830 ;
        RECT 1624.360 1062.510 1624.620 1062.830 ;
        RECT 1623.040 1038.770 1623.180 1062.510 ;
        RECT 1623.040 1038.630 1623.640 1038.770 ;
        RECT 1623.500 966.270 1623.640 1038.630 ;
        RECT 1622.980 965.950 1623.240 966.270 ;
        RECT 1623.440 965.950 1623.700 966.270 ;
        RECT 1623.040 931.330 1623.180 965.950 ;
        RECT 1623.040 931.190 1623.640 931.330 ;
        RECT 1623.500 910.850 1623.640 931.190 ;
        RECT 1622.520 910.530 1622.780 910.850 ;
        RECT 1623.440 910.530 1623.700 910.850 ;
        RECT 1622.580 862.765 1622.720 910.530 ;
        RECT 1622.510 862.395 1622.790 862.765 ;
        RECT 1623.430 862.395 1623.710 862.765 ;
        RECT 1623.500 821.090 1623.640 862.395 ;
        RECT 1623.440 820.770 1623.700 821.090 ;
        RECT 1622.980 772.830 1623.240 773.150 ;
        RECT 1623.040 738.810 1623.180 772.830 ;
        RECT 1622.980 738.490 1623.240 738.810 ;
        RECT 1622.980 737.810 1623.240 738.130 ;
        RECT 1623.040 724.725 1623.180 737.810 ;
        RECT 1622.970 724.355 1623.250 724.725 ;
        RECT 1623.890 724.355 1624.170 724.725 ;
        RECT 1623.960 677.125 1624.100 724.355 ;
        RECT 1623.890 676.755 1624.170 677.125 ;
        RECT 1622.970 676.075 1623.250 676.445 ;
        RECT 1623.040 655.510 1623.180 676.075 ;
        RECT 1622.980 655.190 1623.240 655.510 ;
        RECT 1624.360 655.190 1624.620 655.510 ;
        RECT 1624.420 579.885 1624.560 655.190 ;
        RECT 1623.430 579.515 1623.710 579.885 ;
        RECT 1624.350 579.515 1624.630 579.885 ;
        RECT 1623.500 531.750 1623.640 579.515 ;
        RECT 1623.440 531.430 1623.700 531.750 ;
        RECT 1623.440 524.290 1623.700 524.610 ;
        RECT 1623.500 497.410 1623.640 524.290 ;
        RECT 1623.440 497.090 1623.700 497.410 ;
        RECT 1622.980 496.410 1623.240 496.730 ;
        RECT 1623.040 412.070 1623.180 496.410 ;
        RECT 1622.980 411.750 1623.240 412.070 ;
        RECT 1622.980 411.070 1623.240 411.390 ;
        RECT 1623.040 338.970 1623.180 411.070 ;
        RECT 1622.980 338.650 1623.240 338.970 ;
        RECT 1622.980 337.970 1623.240 338.290 ;
        RECT 1623.040 331.150 1623.180 337.970 ;
        RECT 1622.980 330.830 1623.240 331.150 ;
        RECT 1623.900 265.210 1624.160 265.530 ;
        RECT 1623.960 193.110 1624.100 265.210 ;
        RECT 1623.900 192.790 1624.160 193.110 ;
        RECT 1623.900 192.110 1624.160 192.430 ;
        RECT 1623.960 168.370 1624.100 192.110 ;
        RECT 1623.040 168.230 1624.100 168.370 ;
        RECT 1623.040 144.830 1623.180 168.230 ;
        RECT 1622.980 144.510 1623.240 144.830 ;
        RECT 1622.980 96.570 1623.240 96.890 ;
        RECT 1623.040 39.770 1623.180 96.570 ;
        RECT 1263.260 39.450 1263.520 39.770 ;
        RECT 1622.980 39.450 1623.240 39.770 ;
        RECT 1263.320 2.400 1263.460 39.450 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
      LAYER via2 ;
        RECT 1625.730 1691.360 1626.010 1691.640 ;
        RECT 1622.970 1690.680 1623.250 1690.960 ;
        RECT 1622.970 1255.480 1623.250 1255.760 ;
        RECT 1623.890 1255.480 1624.170 1255.760 ;
        RECT 1622.970 1158.920 1623.250 1159.200 ;
        RECT 1624.350 1158.920 1624.630 1159.200 ;
        RECT 1622.510 862.440 1622.790 862.720 ;
        RECT 1623.430 862.440 1623.710 862.720 ;
        RECT 1622.970 724.400 1623.250 724.680 ;
        RECT 1623.890 724.400 1624.170 724.680 ;
        RECT 1623.890 676.800 1624.170 677.080 ;
        RECT 1622.970 676.120 1623.250 676.400 ;
        RECT 1623.430 579.560 1623.710 579.840 ;
        RECT 1624.350 579.560 1624.630 579.840 ;
      LAYER met3 ;
        RECT 1625.705 1691.650 1626.035 1691.665 ;
        RECT 1622.270 1691.350 1626.035 1691.650 ;
        RECT 1622.270 1690.970 1622.570 1691.350 ;
        RECT 1625.705 1691.335 1626.035 1691.350 ;
        RECT 1622.945 1690.970 1623.275 1690.985 ;
        RECT 1622.270 1690.670 1623.275 1690.970 ;
        RECT 1622.945 1690.655 1623.275 1690.670 ;
        RECT 1622.945 1255.770 1623.275 1255.785 ;
        RECT 1623.865 1255.770 1624.195 1255.785 ;
        RECT 1622.945 1255.470 1624.195 1255.770 ;
        RECT 1622.945 1255.455 1623.275 1255.470 ;
        RECT 1623.865 1255.455 1624.195 1255.470 ;
        RECT 1622.945 1159.210 1623.275 1159.225 ;
        RECT 1624.325 1159.210 1624.655 1159.225 ;
        RECT 1622.945 1158.910 1624.655 1159.210 ;
        RECT 1622.945 1158.895 1623.275 1158.910 ;
        RECT 1624.325 1158.895 1624.655 1158.910 ;
        RECT 1622.485 862.730 1622.815 862.745 ;
        RECT 1623.405 862.730 1623.735 862.745 ;
        RECT 1622.485 862.430 1623.735 862.730 ;
        RECT 1622.485 862.415 1622.815 862.430 ;
        RECT 1623.405 862.415 1623.735 862.430 ;
        RECT 1622.945 724.690 1623.275 724.705 ;
        RECT 1623.865 724.690 1624.195 724.705 ;
        RECT 1622.945 724.390 1624.195 724.690 ;
        RECT 1622.945 724.375 1623.275 724.390 ;
        RECT 1623.865 724.375 1624.195 724.390 ;
        RECT 1623.865 677.090 1624.195 677.105 ;
        RECT 1622.270 676.790 1624.195 677.090 ;
        RECT 1622.270 676.410 1622.570 676.790 ;
        RECT 1623.865 676.775 1624.195 676.790 ;
        RECT 1622.945 676.410 1623.275 676.425 ;
        RECT 1622.270 676.110 1623.275 676.410 ;
        RECT 1622.945 676.095 1623.275 676.110 ;
        RECT 1623.405 579.850 1623.735 579.865 ;
        RECT 1624.325 579.850 1624.655 579.865 ;
        RECT 1623.405 579.550 1624.655 579.850 ;
        RECT 1623.405 579.535 1623.735 579.550 ;
        RECT 1624.325 579.535 1624.655 579.550 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1629.925 1449.165 1630.095 1473.475 ;
      LAYER mcon ;
        RECT 1629.925 1473.305 1630.095 1473.475 ;
      LAYER met1 ;
        RECT 1629.850 1607.900 1630.170 1608.160 ;
        RECT 1629.940 1607.080 1630.080 1607.900 ;
        RECT 1630.310 1607.080 1630.630 1607.140 ;
        RECT 1629.940 1606.940 1630.630 1607.080 ;
        RECT 1630.310 1606.880 1630.630 1606.940 ;
        RECT 1629.865 1473.460 1630.155 1473.505 ;
        RECT 1630.310 1473.460 1630.630 1473.520 ;
        RECT 1629.865 1473.320 1630.630 1473.460 ;
        RECT 1629.865 1473.275 1630.155 1473.320 ;
        RECT 1630.310 1473.260 1630.630 1473.320 ;
        RECT 1629.850 1449.320 1630.170 1449.380 ;
        RECT 1629.655 1449.180 1630.170 1449.320 ;
        RECT 1629.850 1449.120 1630.170 1449.180 ;
        RECT 1629.850 1365.820 1630.170 1366.080 ;
        RECT 1629.940 1365.400 1630.080 1365.820 ;
        RECT 1629.850 1365.140 1630.170 1365.400 ;
        RECT 1629.850 1269.260 1630.170 1269.520 ;
        RECT 1629.940 1268.840 1630.080 1269.260 ;
        RECT 1629.850 1268.580 1630.170 1268.840 ;
        RECT 1629.850 1172.700 1630.170 1172.960 ;
        RECT 1629.940 1172.280 1630.080 1172.700 ;
        RECT 1629.850 1172.020 1630.170 1172.280 ;
        RECT 1629.850 1076.140 1630.170 1076.400 ;
        RECT 1629.940 1075.720 1630.080 1076.140 ;
        RECT 1629.850 1075.460 1630.170 1075.720 ;
        RECT 1629.850 979.580 1630.170 979.840 ;
        RECT 1629.940 979.160 1630.080 979.580 ;
        RECT 1629.850 978.900 1630.170 979.160 ;
        RECT 1629.850 786.460 1630.170 786.720 ;
        RECT 1629.940 786.040 1630.080 786.460 ;
        RECT 1629.850 785.780 1630.170 786.040 ;
        RECT 1629.850 400.220 1630.170 400.480 ;
        RECT 1629.940 399.800 1630.080 400.220 ;
        RECT 1629.850 399.540 1630.170 399.800 ;
        RECT 1629.850 338.540 1630.170 338.600 ;
        RECT 1629.480 338.400 1630.170 338.540 ;
        RECT 1629.480 338.260 1629.620 338.400 ;
        RECT 1629.850 338.340 1630.170 338.400 ;
        RECT 1629.390 338.000 1629.710 338.260 ;
        RECT 1629.390 290.060 1629.710 290.320 ;
        RECT 1629.480 289.640 1629.620 290.060 ;
        RECT 1629.390 289.380 1629.710 289.640 ;
        RECT 1629.390 234.160 1629.710 234.220 ;
        RECT 1630.770 234.160 1631.090 234.220 ;
        RECT 1629.390 234.020 1631.090 234.160 ;
        RECT 1629.390 233.960 1629.710 234.020 ;
        RECT 1630.770 233.960 1631.090 234.020 ;
        RECT 1629.850 62.460 1630.170 62.520 ;
        RECT 1629.480 62.320 1630.170 62.460 ;
        RECT 1629.480 62.180 1629.620 62.320 ;
        RECT 1629.850 62.260 1630.170 62.320 ;
        RECT 1629.390 61.920 1629.710 62.180 ;
        RECT 1281.170 40.020 1281.490 40.080 ;
        RECT 1629.390 40.020 1629.710 40.080 ;
        RECT 1281.170 39.880 1629.710 40.020 ;
        RECT 1281.170 39.820 1281.490 39.880 ;
        RECT 1629.390 39.820 1629.710 39.880 ;
      LAYER via ;
        RECT 1629.880 1607.900 1630.140 1608.160 ;
        RECT 1630.340 1606.880 1630.600 1607.140 ;
        RECT 1630.340 1473.260 1630.600 1473.520 ;
        RECT 1629.880 1449.120 1630.140 1449.380 ;
        RECT 1629.880 1365.820 1630.140 1366.080 ;
        RECT 1629.880 1365.140 1630.140 1365.400 ;
        RECT 1629.880 1269.260 1630.140 1269.520 ;
        RECT 1629.880 1268.580 1630.140 1268.840 ;
        RECT 1629.880 1172.700 1630.140 1172.960 ;
        RECT 1629.880 1172.020 1630.140 1172.280 ;
        RECT 1629.880 1076.140 1630.140 1076.400 ;
        RECT 1629.880 1075.460 1630.140 1075.720 ;
        RECT 1629.880 979.580 1630.140 979.840 ;
        RECT 1629.880 978.900 1630.140 979.160 ;
        RECT 1629.880 786.460 1630.140 786.720 ;
        RECT 1629.880 785.780 1630.140 786.040 ;
        RECT 1629.880 400.220 1630.140 400.480 ;
        RECT 1629.880 399.540 1630.140 399.800 ;
        RECT 1629.880 338.340 1630.140 338.600 ;
        RECT 1629.420 338.000 1629.680 338.260 ;
        RECT 1629.420 290.060 1629.680 290.320 ;
        RECT 1629.420 289.380 1629.680 289.640 ;
        RECT 1629.420 233.960 1629.680 234.220 ;
        RECT 1630.800 233.960 1631.060 234.220 ;
        RECT 1629.880 62.260 1630.140 62.520 ;
        RECT 1629.420 61.920 1629.680 62.180 ;
        RECT 1281.200 39.820 1281.460 40.080 ;
        RECT 1629.420 39.820 1629.680 40.080 ;
      LAYER met2 ;
        RECT 1632.565 1700.410 1632.845 1704.000 ;
        RECT 1631.320 1700.270 1632.845 1700.410 ;
        RECT 1631.320 1677.970 1631.460 1700.270 ;
        RECT 1632.565 1700.000 1632.845 1700.270 ;
        RECT 1629.940 1677.830 1631.460 1677.970 ;
        RECT 1629.940 1608.190 1630.080 1677.830 ;
        RECT 1629.880 1607.870 1630.140 1608.190 ;
        RECT 1630.340 1606.850 1630.600 1607.170 ;
        RECT 1630.400 1473.550 1630.540 1606.850 ;
        RECT 1630.340 1473.230 1630.600 1473.550 ;
        RECT 1629.880 1449.090 1630.140 1449.410 ;
        RECT 1629.940 1366.110 1630.080 1449.090 ;
        RECT 1629.880 1365.790 1630.140 1366.110 ;
        RECT 1629.880 1365.110 1630.140 1365.430 ;
        RECT 1629.940 1269.550 1630.080 1365.110 ;
        RECT 1629.880 1269.230 1630.140 1269.550 ;
        RECT 1629.880 1268.550 1630.140 1268.870 ;
        RECT 1629.940 1172.990 1630.080 1268.550 ;
        RECT 1629.880 1172.670 1630.140 1172.990 ;
        RECT 1629.880 1171.990 1630.140 1172.310 ;
        RECT 1629.940 1076.430 1630.080 1171.990 ;
        RECT 1629.880 1076.110 1630.140 1076.430 ;
        RECT 1629.880 1075.430 1630.140 1075.750 ;
        RECT 1629.940 979.870 1630.080 1075.430 ;
        RECT 1629.880 979.550 1630.140 979.870 ;
        RECT 1629.880 978.870 1630.140 979.190 ;
        RECT 1629.940 883.730 1630.080 978.870 ;
        RECT 1629.480 883.590 1630.080 883.730 ;
        RECT 1629.480 883.050 1629.620 883.590 ;
        RECT 1629.480 882.910 1630.080 883.050 ;
        RECT 1629.940 786.750 1630.080 882.910 ;
        RECT 1629.880 786.430 1630.140 786.750 ;
        RECT 1629.880 785.750 1630.140 786.070 ;
        RECT 1629.940 497.490 1630.080 785.750 ;
        RECT 1629.480 497.350 1630.080 497.490 ;
        RECT 1629.480 496.810 1629.620 497.350 ;
        RECT 1629.480 496.670 1630.080 496.810 ;
        RECT 1629.940 400.510 1630.080 496.670 ;
        RECT 1629.880 400.190 1630.140 400.510 ;
        RECT 1629.880 399.510 1630.140 399.830 ;
        RECT 1629.940 338.630 1630.080 399.510 ;
        RECT 1629.880 338.310 1630.140 338.630 ;
        RECT 1629.420 337.970 1629.680 338.290 ;
        RECT 1629.480 290.350 1629.620 337.970 ;
        RECT 1629.420 290.030 1629.680 290.350 ;
        RECT 1629.420 289.350 1629.680 289.670 ;
        RECT 1629.480 234.250 1629.620 289.350 ;
        RECT 1629.420 233.930 1629.680 234.250 ;
        RECT 1630.800 233.930 1631.060 234.250 ;
        RECT 1630.860 192.850 1631.000 233.930 ;
        RECT 1630.400 192.710 1631.000 192.850 ;
        RECT 1630.400 122.130 1630.540 192.710 ;
        RECT 1629.940 121.990 1630.540 122.130 ;
        RECT 1629.940 62.550 1630.080 121.990 ;
        RECT 1629.880 62.230 1630.140 62.550 ;
        RECT 1629.420 61.890 1629.680 62.210 ;
        RECT 1629.480 40.110 1629.620 61.890 ;
        RECT 1281.200 39.790 1281.460 40.110 ;
        RECT 1629.420 39.790 1629.680 40.110 ;
        RECT 1281.260 2.400 1281.400 39.790 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1637.285 1642.285 1637.455 1656.055 ;
        RECT 1637.285 1545.725 1637.455 1593.835 ;
        RECT 1636.365 1442.025 1636.535 1490.475 ;
        RECT 1636.365 1213.205 1636.535 1255.875 ;
        RECT 1636.825 855.525 1636.995 903.975 ;
        RECT 1636.825 737.885 1636.995 767.635 ;
        RECT 1636.825 641.325 1636.995 676.175 ;
        RECT 1636.825 476.085 1636.995 524.195 ;
        RECT 1636.825 386.325 1636.995 434.435 ;
        RECT 1636.825 331.245 1636.995 338.215 ;
        RECT 1636.365 48.365 1636.535 96.475 ;
      LAYER mcon ;
        RECT 1637.285 1655.885 1637.455 1656.055 ;
        RECT 1637.285 1593.665 1637.455 1593.835 ;
        RECT 1636.365 1490.305 1636.535 1490.475 ;
        RECT 1636.365 1255.705 1636.535 1255.875 ;
        RECT 1636.825 903.805 1636.995 903.975 ;
        RECT 1636.825 767.465 1636.995 767.635 ;
        RECT 1636.825 676.005 1636.995 676.175 ;
        RECT 1636.825 524.025 1636.995 524.195 ;
        RECT 1636.825 434.265 1636.995 434.435 ;
        RECT 1636.825 338.045 1636.995 338.215 ;
        RECT 1636.365 96.305 1636.535 96.475 ;
      LAYER met1 ;
        RECT 1637.210 1656.040 1637.530 1656.100 ;
        RECT 1637.015 1655.900 1637.530 1656.040 ;
        RECT 1637.210 1655.840 1637.530 1655.900 ;
        RECT 1637.210 1642.440 1637.530 1642.500 ;
        RECT 1637.015 1642.300 1637.530 1642.440 ;
        RECT 1637.210 1642.240 1637.530 1642.300 ;
        RECT 1637.210 1593.820 1637.530 1593.880 ;
        RECT 1637.015 1593.680 1637.530 1593.820 ;
        RECT 1637.210 1593.620 1637.530 1593.680 ;
        RECT 1637.210 1545.880 1637.530 1545.940 ;
        RECT 1637.015 1545.740 1637.530 1545.880 ;
        RECT 1637.210 1545.680 1637.530 1545.740 ;
        RECT 1636.290 1497.260 1636.610 1497.320 ;
        RECT 1637.210 1497.260 1637.530 1497.320 ;
        RECT 1636.290 1497.120 1637.530 1497.260 ;
        RECT 1636.290 1497.060 1636.610 1497.120 ;
        RECT 1637.210 1497.060 1637.530 1497.120 ;
        RECT 1636.290 1490.460 1636.610 1490.520 ;
        RECT 1636.095 1490.320 1636.610 1490.460 ;
        RECT 1636.290 1490.260 1636.610 1490.320 ;
        RECT 1636.305 1442.180 1636.595 1442.225 ;
        RECT 1637.670 1442.180 1637.990 1442.240 ;
        RECT 1636.305 1442.040 1637.990 1442.180 ;
        RECT 1636.305 1441.995 1636.595 1442.040 ;
        RECT 1637.670 1441.980 1637.990 1442.040 ;
        RECT 1637.670 1400.700 1637.990 1400.760 ;
        RECT 1636.840 1400.560 1637.990 1400.700 ;
        RECT 1636.840 1400.420 1636.980 1400.560 ;
        RECT 1637.670 1400.500 1637.990 1400.560 ;
        RECT 1636.750 1400.160 1637.070 1400.420 ;
        RECT 1636.305 1255.860 1636.595 1255.905 ;
        RECT 1636.750 1255.860 1637.070 1255.920 ;
        RECT 1636.305 1255.720 1637.070 1255.860 ;
        RECT 1636.305 1255.675 1636.595 1255.720 ;
        RECT 1636.750 1255.660 1637.070 1255.720 ;
        RECT 1636.290 1213.360 1636.610 1213.420 ;
        RECT 1636.095 1213.220 1636.610 1213.360 ;
        RECT 1636.290 1213.160 1636.610 1213.220 ;
        RECT 1636.290 1200.440 1636.610 1200.500 ;
        RECT 1636.750 1200.440 1637.070 1200.500 ;
        RECT 1636.290 1200.300 1637.070 1200.440 ;
        RECT 1636.290 1200.240 1636.610 1200.300 ;
        RECT 1636.750 1200.240 1637.070 1200.300 ;
        RECT 1636.750 1104.220 1637.070 1104.280 ;
        RECT 1637.670 1104.220 1637.990 1104.280 ;
        RECT 1636.750 1104.080 1637.990 1104.220 ;
        RECT 1636.750 1104.020 1637.070 1104.080 ;
        RECT 1637.670 1104.020 1637.990 1104.080 ;
        RECT 1636.750 1076.820 1637.070 1077.080 ;
        RECT 1636.840 1076.400 1636.980 1076.820 ;
        RECT 1636.750 1076.140 1637.070 1076.400 ;
        RECT 1636.750 1055.600 1637.070 1055.660 ;
        RECT 1637.670 1055.600 1637.990 1055.660 ;
        RECT 1636.750 1055.460 1637.990 1055.600 ;
        RECT 1636.750 1055.400 1637.070 1055.460 ;
        RECT 1637.670 1055.400 1637.990 1055.460 ;
        RECT 1636.750 980.260 1637.070 980.520 ;
        RECT 1636.840 979.840 1636.980 980.260 ;
        RECT 1636.750 979.580 1637.070 979.840 ;
        RECT 1636.750 931.640 1637.070 931.900 ;
        RECT 1636.840 931.160 1636.980 931.640 ;
        RECT 1637.210 931.160 1637.530 931.220 ;
        RECT 1636.840 931.020 1637.530 931.160 ;
        RECT 1637.210 930.960 1637.530 931.020 ;
        RECT 1636.765 903.960 1637.055 904.005 ;
        RECT 1637.210 903.960 1637.530 904.020 ;
        RECT 1636.765 903.820 1637.530 903.960 ;
        RECT 1636.765 903.775 1637.055 903.820 ;
        RECT 1637.210 903.760 1637.530 903.820 ;
        RECT 1636.750 855.680 1637.070 855.740 ;
        RECT 1636.555 855.540 1637.070 855.680 ;
        RECT 1636.750 855.480 1637.070 855.540 ;
        RECT 1636.750 767.620 1637.070 767.680 ;
        RECT 1636.555 767.480 1637.070 767.620 ;
        RECT 1636.750 767.420 1637.070 767.480 ;
        RECT 1636.750 738.040 1637.070 738.100 ;
        RECT 1636.555 737.900 1637.070 738.040 ;
        RECT 1636.750 737.840 1637.070 737.900 ;
        RECT 1636.750 676.160 1637.070 676.220 ;
        RECT 1636.555 676.020 1637.070 676.160 ;
        RECT 1636.750 675.960 1637.070 676.020 ;
        RECT 1636.750 641.480 1637.070 641.540 ;
        RECT 1636.555 641.340 1637.070 641.480 ;
        RECT 1636.750 641.280 1637.070 641.340 ;
        RECT 1636.765 524.180 1637.055 524.225 ;
        RECT 1637.210 524.180 1637.530 524.240 ;
        RECT 1636.765 524.040 1637.530 524.180 ;
        RECT 1636.765 523.995 1637.055 524.040 ;
        RECT 1637.210 523.980 1637.530 524.040 ;
        RECT 1636.750 476.240 1637.070 476.300 ;
        RECT 1636.555 476.100 1637.070 476.240 ;
        RECT 1636.750 476.040 1637.070 476.100 ;
        RECT 1636.750 434.420 1637.070 434.480 ;
        RECT 1636.555 434.280 1637.070 434.420 ;
        RECT 1636.750 434.220 1637.070 434.280 ;
        RECT 1636.750 386.480 1637.070 386.540 ;
        RECT 1636.555 386.340 1637.070 386.480 ;
        RECT 1636.750 386.280 1637.070 386.340 ;
        RECT 1636.750 338.200 1637.070 338.260 ;
        RECT 1636.555 338.060 1637.070 338.200 ;
        RECT 1636.750 338.000 1637.070 338.060 ;
        RECT 1636.750 331.400 1637.070 331.460 ;
        RECT 1636.555 331.260 1637.070 331.400 ;
        RECT 1636.750 331.200 1637.070 331.260 ;
        RECT 1636.750 265.780 1637.070 265.840 ;
        RECT 1636.380 265.640 1637.070 265.780 ;
        RECT 1636.380 265.500 1636.520 265.640 ;
        RECT 1636.750 265.580 1637.070 265.640 ;
        RECT 1636.290 265.240 1636.610 265.500 ;
        RECT 1636.290 144.740 1636.610 144.800 ;
        RECT 1637.210 144.740 1637.530 144.800 ;
        RECT 1636.290 144.600 1637.530 144.740 ;
        RECT 1636.290 144.540 1636.610 144.600 ;
        RECT 1637.210 144.540 1637.530 144.600 ;
        RECT 1636.305 96.460 1636.595 96.505 ;
        RECT 1636.750 96.460 1637.070 96.520 ;
        RECT 1636.305 96.320 1637.070 96.460 ;
        RECT 1636.305 96.275 1636.595 96.320 ;
        RECT 1636.750 96.260 1637.070 96.320 ;
        RECT 1636.290 48.520 1636.610 48.580 ;
        RECT 1636.095 48.380 1636.610 48.520 ;
        RECT 1636.290 48.320 1636.610 48.380 ;
        RECT 1299.110 40.360 1299.430 40.420 ;
        RECT 1636.290 40.360 1636.610 40.420 ;
        RECT 1299.110 40.220 1636.610 40.360 ;
        RECT 1299.110 40.160 1299.430 40.220 ;
        RECT 1636.290 40.160 1636.610 40.220 ;
      LAYER via ;
        RECT 1637.240 1655.840 1637.500 1656.100 ;
        RECT 1637.240 1642.240 1637.500 1642.500 ;
        RECT 1637.240 1593.620 1637.500 1593.880 ;
        RECT 1637.240 1545.680 1637.500 1545.940 ;
        RECT 1636.320 1497.060 1636.580 1497.320 ;
        RECT 1637.240 1497.060 1637.500 1497.320 ;
        RECT 1636.320 1490.260 1636.580 1490.520 ;
        RECT 1637.700 1441.980 1637.960 1442.240 ;
        RECT 1637.700 1400.500 1637.960 1400.760 ;
        RECT 1636.780 1400.160 1637.040 1400.420 ;
        RECT 1636.780 1255.660 1637.040 1255.920 ;
        RECT 1636.320 1213.160 1636.580 1213.420 ;
        RECT 1636.320 1200.240 1636.580 1200.500 ;
        RECT 1636.780 1200.240 1637.040 1200.500 ;
        RECT 1636.780 1104.020 1637.040 1104.280 ;
        RECT 1637.700 1104.020 1637.960 1104.280 ;
        RECT 1636.780 1076.820 1637.040 1077.080 ;
        RECT 1636.780 1076.140 1637.040 1076.400 ;
        RECT 1636.780 1055.400 1637.040 1055.660 ;
        RECT 1637.700 1055.400 1637.960 1055.660 ;
        RECT 1636.780 980.260 1637.040 980.520 ;
        RECT 1636.780 979.580 1637.040 979.840 ;
        RECT 1636.780 931.640 1637.040 931.900 ;
        RECT 1637.240 930.960 1637.500 931.220 ;
        RECT 1637.240 903.760 1637.500 904.020 ;
        RECT 1636.780 855.480 1637.040 855.740 ;
        RECT 1636.780 767.420 1637.040 767.680 ;
        RECT 1636.780 737.840 1637.040 738.100 ;
        RECT 1636.780 675.960 1637.040 676.220 ;
        RECT 1636.780 641.280 1637.040 641.540 ;
        RECT 1637.240 523.980 1637.500 524.240 ;
        RECT 1636.780 476.040 1637.040 476.300 ;
        RECT 1636.780 434.220 1637.040 434.480 ;
        RECT 1636.780 386.280 1637.040 386.540 ;
        RECT 1636.780 338.000 1637.040 338.260 ;
        RECT 1636.780 331.200 1637.040 331.460 ;
        RECT 1636.780 265.580 1637.040 265.840 ;
        RECT 1636.320 265.240 1636.580 265.500 ;
        RECT 1636.320 144.540 1636.580 144.800 ;
        RECT 1637.240 144.540 1637.500 144.800 ;
        RECT 1636.780 96.260 1637.040 96.520 ;
        RECT 1636.320 48.320 1636.580 48.580 ;
        RECT 1299.140 40.160 1299.400 40.420 ;
        RECT 1636.320 40.160 1636.580 40.420 ;
      LAYER met2 ;
        RECT 1639.005 1701.090 1639.285 1704.000 ;
        RECT 1637.300 1700.950 1639.285 1701.090 ;
        RECT 1637.300 1656.130 1637.440 1700.950 ;
        RECT 1639.005 1700.000 1639.285 1700.950 ;
        RECT 1637.240 1655.810 1637.500 1656.130 ;
        RECT 1637.240 1642.210 1637.500 1642.530 ;
        RECT 1637.300 1593.910 1637.440 1642.210 ;
        RECT 1637.240 1593.590 1637.500 1593.910 ;
        RECT 1637.240 1545.650 1637.500 1545.970 ;
        RECT 1637.300 1497.350 1637.440 1545.650 ;
        RECT 1636.320 1497.030 1636.580 1497.350 ;
        RECT 1637.240 1497.030 1637.500 1497.350 ;
        RECT 1636.380 1490.550 1636.520 1497.030 ;
        RECT 1636.320 1490.230 1636.580 1490.550 ;
        RECT 1637.700 1441.950 1637.960 1442.270 ;
        RECT 1637.760 1400.790 1637.900 1441.950 ;
        RECT 1637.700 1400.470 1637.960 1400.790 ;
        RECT 1636.780 1400.130 1637.040 1400.450 ;
        RECT 1636.840 1393.845 1636.980 1400.130 ;
        RECT 1636.770 1393.475 1637.050 1393.845 ;
        RECT 1638.150 1393.475 1638.430 1393.845 ;
        RECT 1638.220 1268.610 1638.360 1393.475 ;
        RECT 1636.840 1268.470 1638.360 1268.610 ;
        RECT 1636.840 1255.950 1636.980 1268.470 ;
        RECT 1636.780 1255.630 1637.040 1255.950 ;
        RECT 1636.320 1213.130 1636.580 1213.450 ;
        RECT 1636.380 1200.530 1636.520 1213.130 ;
        RECT 1636.320 1200.210 1636.580 1200.530 ;
        RECT 1636.780 1200.210 1637.040 1200.530 ;
        RECT 1636.840 1152.445 1636.980 1200.210 ;
        RECT 1636.770 1152.075 1637.050 1152.445 ;
        RECT 1637.690 1152.075 1637.970 1152.445 ;
        RECT 1637.760 1104.310 1637.900 1152.075 ;
        RECT 1636.780 1103.990 1637.040 1104.310 ;
        RECT 1637.700 1103.990 1637.960 1104.310 ;
        RECT 1636.840 1077.110 1636.980 1103.990 ;
        RECT 1636.780 1076.790 1637.040 1077.110 ;
        RECT 1636.780 1076.110 1637.040 1076.430 ;
        RECT 1636.840 1055.690 1636.980 1076.110 ;
        RECT 1636.780 1055.370 1637.040 1055.690 ;
        RECT 1637.700 1055.370 1637.960 1055.690 ;
        RECT 1637.760 1007.605 1637.900 1055.370 ;
        RECT 1636.770 1007.235 1637.050 1007.605 ;
        RECT 1637.690 1007.235 1637.970 1007.605 ;
        RECT 1636.840 980.550 1636.980 1007.235 ;
        RECT 1636.780 980.230 1637.040 980.550 ;
        RECT 1636.780 979.550 1637.040 979.870 ;
        RECT 1636.840 931.930 1636.980 979.550 ;
        RECT 1636.780 931.610 1637.040 931.930 ;
        RECT 1637.240 930.930 1637.500 931.250 ;
        RECT 1637.300 904.050 1637.440 930.930 ;
        RECT 1637.240 903.730 1637.500 904.050 ;
        RECT 1636.780 855.450 1637.040 855.770 ;
        RECT 1636.840 767.710 1636.980 855.450 ;
        RECT 1636.780 767.390 1637.040 767.710 ;
        RECT 1636.780 737.810 1637.040 738.130 ;
        RECT 1636.840 724.610 1636.980 737.810 ;
        RECT 1636.840 724.470 1637.440 724.610 ;
        RECT 1637.300 691.405 1637.440 724.470 ;
        RECT 1637.230 691.035 1637.510 691.405 ;
        RECT 1636.770 676.075 1637.050 676.445 ;
        RECT 1636.780 675.930 1637.040 676.075 ;
        RECT 1636.780 641.250 1637.040 641.570 ;
        RECT 1636.840 628.050 1636.980 641.250 ;
        RECT 1636.840 627.910 1637.440 628.050 ;
        RECT 1637.300 604.250 1637.440 627.910 ;
        RECT 1637.300 604.110 1637.900 604.250 ;
        RECT 1637.760 532.285 1637.900 604.110 ;
        RECT 1637.690 531.915 1637.970 532.285 ;
        RECT 1637.230 531.235 1637.510 531.605 ;
        RECT 1637.300 524.270 1637.440 531.235 ;
        RECT 1637.240 523.950 1637.500 524.270 ;
        RECT 1636.780 476.010 1637.040 476.330 ;
        RECT 1636.840 434.510 1636.980 476.010 ;
        RECT 1636.780 434.190 1637.040 434.510 ;
        RECT 1636.780 386.250 1637.040 386.570 ;
        RECT 1636.840 338.290 1636.980 386.250 ;
        RECT 1636.780 337.970 1637.040 338.290 ;
        RECT 1636.780 331.170 1637.040 331.490 ;
        RECT 1636.840 265.870 1636.980 331.170 ;
        RECT 1636.780 265.550 1637.040 265.870 ;
        RECT 1636.320 265.210 1636.580 265.530 ;
        RECT 1636.380 193.530 1636.520 265.210 ;
        RECT 1636.380 193.390 1636.980 193.530 ;
        RECT 1636.840 169.050 1636.980 193.390 ;
        RECT 1636.380 168.910 1636.980 169.050 ;
        RECT 1636.380 158.170 1636.520 168.910 ;
        RECT 1636.380 158.030 1637.440 158.170 ;
        RECT 1637.300 144.830 1637.440 158.030 ;
        RECT 1636.320 144.510 1636.580 144.830 ;
        RECT 1637.240 144.510 1637.500 144.830 ;
        RECT 1636.380 96.970 1636.520 144.510 ;
        RECT 1636.380 96.830 1636.980 96.970 ;
        RECT 1636.840 96.550 1636.980 96.830 ;
        RECT 1636.780 96.230 1637.040 96.550 ;
        RECT 1636.320 48.290 1636.580 48.610 ;
        RECT 1636.380 40.450 1636.520 48.290 ;
        RECT 1299.140 40.130 1299.400 40.450 ;
        RECT 1636.320 40.130 1636.580 40.450 ;
        RECT 1299.200 2.400 1299.340 40.130 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
      LAYER via2 ;
        RECT 1636.770 1393.520 1637.050 1393.800 ;
        RECT 1638.150 1393.520 1638.430 1393.800 ;
        RECT 1636.770 1152.120 1637.050 1152.400 ;
        RECT 1637.690 1152.120 1637.970 1152.400 ;
        RECT 1636.770 1007.280 1637.050 1007.560 ;
        RECT 1637.690 1007.280 1637.970 1007.560 ;
        RECT 1637.230 691.080 1637.510 691.360 ;
        RECT 1636.770 676.120 1637.050 676.400 ;
        RECT 1637.690 531.960 1637.970 532.240 ;
        RECT 1637.230 531.280 1637.510 531.560 ;
      LAYER met3 ;
        RECT 1636.745 1393.810 1637.075 1393.825 ;
        RECT 1638.125 1393.810 1638.455 1393.825 ;
        RECT 1636.745 1393.510 1638.455 1393.810 ;
        RECT 1636.745 1393.495 1637.075 1393.510 ;
        RECT 1638.125 1393.495 1638.455 1393.510 ;
        RECT 1636.745 1152.410 1637.075 1152.425 ;
        RECT 1637.665 1152.410 1637.995 1152.425 ;
        RECT 1636.745 1152.110 1637.995 1152.410 ;
        RECT 1636.745 1152.095 1637.075 1152.110 ;
        RECT 1637.665 1152.095 1637.995 1152.110 ;
        RECT 1636.745 1007.570 1637.075 1007.585 ;
        RECT 1637.665 1007.570 1637.995 1007.585 ;
        RECT 1636.745 1007.270 1637.995 1007.570 ;
        RECT 1636.745 1007.255 1637.075 1007.270 ;
        RECT 1637.665 1007.255 1637.995 1007.270 ;
        RECT 1637.205 691.380 1637.535 691.385 ;
        RECT 1636.950 691.370 1637.535 691.380 ;
        RECT 1636.750 691.070 1637.535 691.370 ;
        RECT 1636.950 691.060 1637.535 691.070 ;
        RECT 1637.205 691.055 1637.535 691.060 ;
        RECT 1636.745 676.420 1637.075 676.425 ;
        RECT 1636.745 676.410 1637.330 676.420 ;
        RECT 1636.520 676.110 1637.330 676.410 ;
        RECT 1636.745 676.100 1637.330 676.110 ;
        RECT 1636.745 676.095 1637.075 676.100 ;
        RECT 1637.665 532.250 1637.995 532.265 ;
        RECT 1636.990 531.950 1637.995 532.250 ;
        RECT 1636.990 531.585 1637.290 531.950 ;
        RECT 1637.665 531.935 1637.995 531.950 ;
        RECT 1636.990 531.270 1637.535 531.585 ;
        RECT 1637.205 531.255 1637.535 531.270 ;
      LAYER via3 ;
        RECT 1636.980 691.060 1637.300 691.380 ;
        RECT 1636.980 676.100 1637.300 676.420 ;
      LAYER met4 ;
        RECT 1636.975 691.055 1637.305 691.385 ;
        RECT 1636.990 676.425 1637.290 691.055 ;
        RECT 1636.975 676.095 1637.305 676.425 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1642.345 593.045 1642.515 627.895 ;
        RECT 1642.805 138.125 1642.975 159.375 ;
        RECT 1642.345 61.625 1642.515 113.815 ;
      LAYER mcon ;
        RECT 1642.345 627.725 1642.515 627.895 ;
        RECT 1642.805 159.205 1642.975 159.375 ;
        RECT 1642.345 113.645 1642.515 113.815 ;
      LAYER met1 ;
        RECT 1642.730 1642.440 1643.050 1642.500 ;
        RECT 1644.110 1642.440 1644.430 1642.500 ;
        RECT 1642.730 1642.300 1644.430 1642.440 ;
        RECT 1642.730 1642.240 1643.050 1642.300 ;
        RECT 1644.110 1642.240 1644.430 1642.300 ;
        RECT 1642.730 1593.820 1643.050 1593.880 ;
        RECT 1643.650 1593.820 1643.970 1593.880 ;
        RECT 1642.730 1593.680 1643.970 1593.820 ;
        RECT 1642.730 1593.620 1643.050 1593.680 ;
        RECT 1643.650 1593.620 1643.970 1593.680 ;
        RECT 1642.730 1462.920 1643.050 1462.980 ;
        RECT 1643.650 1462.920 1643.970 1462.980 ;
        RECT 1642.730 1462.780 1643.970 1462.920 ;
        RECT 1642.730 1462.720 1643.050 1462.780 ;
        RECT 1643.650 1462.720 1643.970 1462.780 ;
        RECT 1642.730 676.160 1643.050 676.220 ;
        RECT 1643.650 676.160 1643.970 676.220 ;
        RECT 1642.730 676.020 1643.970 676.160 ;
        RECT 1642.730 675.960 1643.050 676.020 ;
        RECT 1643.650 675.960 1643.970 676.020 ;
        RECT 1642.270 627.880 1642.590 627.940 ;
        RECT 1642.270 627.740 1642.785 627.880 ;
        RECT 1642.270 627.680 1642.590 627.740 ;
        RECT 1642.285 593.200 1642.575 593.245 ;
        RECT 1642.730 593.200 1643.050 593.260 ;
        RECT 1642.285 593.060 1643.050 593.200 ;
        RECT 1642.285 593.015 1642.575 593.060 ;
        RECT 1642.730 593.000 1643.050 593.060 ;
        RECT 1642.730 352.280 1643.050 352.540 ;
        RECT 1642.820 351.860 1642.960 352.280 ;
        RECT 1642.730 351.600 1643.050 351.860 ;
        RECT 1642.730 159.360 1643.050 159.420 ;
        RECT 1642.535 159.220 1643.050 159.360 ;
        RECT 1642.730 159.160 1643.050 159.220 ;
        RECT 1642.730 138.280 1643.050 138.340 ;
        RECT 1642.535 138.140 1643.050 138.280 ;
        RECT 1642.730 138.080 1643.050 138.140 ;
        RECT 1642.285 113.800 1642.575 113.845 ;
        RECT 1642.730 113.800 1643.050 113.860 ;
        RECT 1642.285 113.660 1643.050 113.800 ;
        RECT 1642.285 113.615 1642.575 113.660 ;
        RECT 1642.730 113.600 1643.050 113.660 ;
        RECT 1642.285 61.780 1642.575 61.825 ;
        RECT 1642.730 61.780 1643.050 61.840 ;
        RECT 1642.285 61.640 1643.050 61.780 ;
        RECT 1642.285 61.595 1642.575 61.640 ;
        RECT 1642.730 61.580 1643.050 61.640 ;
        RECT 1317.050 40.700 1317.370 40.760 ;
        RECT 1642.270 40.700 1642.590 40.760 ;
        RECT 1317.050 40.560 1642.590 40.700 ;
        RECT 1317.050 40.500 1317.370 40.560 ;
        RECT 1642.270 40.500 1642.590 40.560 ;
      LAYER via ;
        RECT 1642.760 1642.240 1643.020 1642.500 ;
        RECT 1644.140 1642.240 1644.400 1642.500 ;
        RECT 1642.760 1593.620 1643.020 1593.880 ;
        RECT 1643.680 1593.620 1643.940 1593.880 ;
        RECT 1642.760 1462.720 1643.020 1462.980 ;
        RECT 1643.680 1462.720 1643.940 1462.980 ;
        RECT 1642.760 675.960 1643.020 676.220 ;
        RECT 1643.680 675.960 1643.940 676.220 ;
        RECT 1642.300 627.680 1642.560 627.940 ;
        RECT 1642.760 593.000 1643.020 593.260 ;
        RECT 1642.760 352.280 1643.020 352.540 ;
        RECT 1642.760 351.600 1643.020 351.860 ;
        RECT 1642.760 159.160 1643.020 159.420 ;
        RECT 1642.760 138.080 1643.020 138.340 ;
        RECT 1642.760 113.600 1643.020 113.860 ;
        RECT 1642.760 61.580 1643.020 61.840 ;
        RECT 1317.080 40.500 1317.340 40.760 ;
        RECT 1642.300 40.500 1642.560 40.760 ;
      LAYER met2 ;
        RECT 1645.905 1700.410 1646.185 1704.000 ;
        RECT 1644.200 1700.270 1646.185 1700.410 ;
        RECT 1644.200 1642.530 1644.340 1700.270 ;
        RECT 1645.905 1700.000 1646.185 1700.270 ;
        RECT 1642.760 1642.210 1643.020 1642.530 ;
        RECT 1644.140 1642.210 1644.400 1642.530 ;
        RECT 1642.820 1593.910 1642.960 1642.210 ;
        RECT 1642.760 1593.590 1643.020 1593.910 ;
        RECT 1643.680 1593.590 1643.940 1593.910 ;
        RECT 1643.740 1463.010 1643.880 1593.590 ;
        RECT 1642.760 1462.690 1643.020 1463.010 ;
        RECT 1643.680 1462.690 1643.940 1463.010 ;
        RECT 1642.820 1414.810 1642.960 1462.690 ;
        RECT 1642.360 1414.670 1642.960 1414.810 ;
        RECT 1642.360 1414.130 1642.500 1414.670 ;
        RECT 1642.360 1413.990 1642.960 1414.130 ;
        RECT 1642.820 1318.250 1642.960 1413.990 ;
        RECT 1642.360 1318.110 1642.960 1318.250 ;
        RECT 1642.360 1317.570 1642.500 1318.110 ;
        RECT 1642.360 1317.430 1642.960 1317.570 ;
        RECT 1642.820 1221.690 1642.960 1317.430 ;
        RECT 1642.360 1221.550 1642.960 1221.690 ;
        RECT 1642.360 1221.010 1642.500 1221.550 ;
        RECT 1642.360 1220.870 1642.960 1221.010 ;
        RECT 1642.820 1125.130 1642.960 1220.870 ;
        RECT 1642.360 1124.990 1642.960 1125.130 ;
        RECT 1642.360 1124.450 1642.500 1124.990 ;
        RECT 1642.360 1124.310 1642.960 1124.450 ;
        RECT 1642.820 1028.570 1642.960 1124.310 ;
        RECT 1642.360 1028.430 1642.960 1028.570 ;
        RECT 1642.360 1027.890 1642.500 1028.430 ;
        RECT 1642.360 1027.750 1642.960 1027.890 ;
        RECT 1642.820 932.010 1642.960 1027.750 ;
        RECT 1642.360 931.870 1642.960 932.010 ;
        RECT 1642.360 931.330 1642.500 931.870 ;
        RECT 1642.360 931.190 1642.960 931.330 ;
        RECT 1642.820 835.450 1642.960 931.190 ;
        RECT 1642.360 835.310 1642.960 835.450 ;
        RECT 1642.360 834.770 1642.500 835.310 ;
        RECT 1642.360 834.630 1642.960 834.770 ;
        RECT 1642.820 738.890 1642.960 834.630 ;
        RECT 1642.360 738.750 1642.960 738.890 ;
        RECT 1642.360 738.210 1642.500 738.750 ;
        RECT 1642.360 738.070 1642.960 738.210 ;
        RECT 1642.820 676.250 1642.960 738.070 ;
        RECT 1642.760 675.930 1643.020 676.250 ;
        RECT 1643.680 675.930 1643.940 676.250 ;
        RECT 1643.740 628.165 1643.880 675.930 ;
        RECT 1642.290 627.795 1642.570 628.165 ;
        RECT 1643.670 627.795 1643.950 628.165 ;
        RECT 1642.300 627.650 1642.560 627.795 ;
        RECT 1642.760 592.970 1643.020 593.290 ;
        RECT 1642.820 545.770 1642.960 592.970 ;
        RECT 1642.360 545.630 1642.960 545.770 ;
        RECT 1642.360 545.090 1642.500 545.630 ;
        RECT 1642.360 544.950 1642.960 545.090 ;
        RECT 1642.820 449.210 1642.960 544.950 ;
        RECT 1642.360 449.070 1642.960 449.210 ;
        RECT 1642.360 448.530 1642.500 449.070 ;
        RECT 1642.360 448.390 1642.960 448.530 ;
        RECT 1642.820 352.570 1642.960 448.390 ;
        RECT 1642.760 352.250 1643.020 352.570 ;
        RECT 1642.760 351.570 1643.020 351.890 ;
        RECT 1642.820 255.410 1642.960 351.570 ;
        RECT 1642.360 255.270 1642.960 255.410 ;
        RECT 1642.360 254.730 1642.500 255.270 ;
        RECT 1642.360 254.590 1642.960 254.730 ;
        RECT 1642.820 159.450 1642.960 254.590 ;
        RECT 1642.760 159.130 1643.020 159.450 ;
        RECT 1642.760 138.050 1643.020 138.370 ;
        RECT 1642.820 113.890 1642.960 138.050 ;
        RECT 1642.760 113.570 1643.020 113.890 ;
        RECT 1642.760 61.550 1643.020 61.870 ;
        RECT 1642.820 48.010 1642.960 61.550 ;
        RECT 1642.360 47.870 1642.960 48.010 ;
        RECT 1642.360 40.790 1642.500 47.870 ;
        RECT 1317.080 40.470 1317.340 40.790 ;
        RECT 1642.300 40.470 1642.560 40.790 ;
        RECT 1317.140 2.400 1317.280 40.470 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 1642.290 627.840 1642.570 628.120 ;
        RECT 1643.670 627.840 1643.950 628.120 ;
      LAYER met3 ;
        RECT 1642.265 628.130 1642.595 628.145 ;
        RECT 1643.645 628.130 1643.975 628.145 ;
        RECT 1642.265 627.830 1643.975 628.130 ;
        RECT 1642.265 627.815 1642.595 627.830 ;
        RECT 1643.645 627.815 1643.975 627.830 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1649.630 1678.140 1649.950 1678.200 ;
        RECT 1651.470 1678.140 1651.790 1678.200 ;
        RECT 1649.630 1678.000 1651.790 1678.140 ;
        RECT 1649.630 1677.940 1649.950 1678.000 ;
        RECT 1651.470 1677.940 1651.790 1678.000 ;
        RECT 1334.990 41.040 1335.310 41.100 ;
        RECT 1649.630 41.040 1649.950 41.100 ;
        RECT 1334.990 40.900 1649.950 41.040 ;
        RECT 1334.990 40.840 1335.310 40.900 ;
        RECT 1649.630 40.840 1649.950 40.900 ;
      LAYER via ;
        RECT 1649.660 1677.940 1649.920 1678.200 ;
        RECT 1651.500 1677.940 1651.760 1678.200 ;
        RECT 1335.020 40.840 1335.280 41.100 ;
        RECT 1649.660 40.840 1649.920 41.100 ;
      LAYER met2 ;
        RECT 1652.805 1700.410 1653.085 1704.000 ;
        RECT 1651.560 1700.270 1653.085 1700.410 ;
        RECT 1651.560 1678.230 1651.700 1700.270 ;
        RECT 1652.805 1700.000 1653.085 1700.270 ;
        RECT 1649.660 1677.910 1649.920 1678.230 ;
        RECT 1651.500 1677.910 1651.760 1678.230 ;
        RECT 1649.720 41.130 1649.860 1677.910 ;
        RECT 1335.020 40.810 1335.280 41.130 ;
        RECT 1649.660 40.810 1649.920 41.130 ;
        RECT 1335.080 2.400 1335.220 40.810 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 37.640 692.690 37.700 ;
        RECT 1409.050 37.640 1409.370 37.700 ;
        RECT 692.370 37.500 1409.370 37.640 ;
        RECT 692.370 37.440 692.690 37.500 ;
        RECT 1409.050 37.440 1409.370 37.500 ;
      LAYER via ;
        RECT 692.400 37.440 692.660 37.700 ;
        RECT 1409.080 37.440 1409.340 37.700 ;
      LAYER met2 ;
        RECT 1410.385 1700.410 1410.665 1704.000 ;
        RECT 1409.140 1700.270 1410.665 1700.410 ;
        RECT 1409.140 37.730 1409.280 1700.270 ;
        RECT 1410.385 1700.000 1410.665 1700.270 ;
        RECT 692.400 37.410 692.660 37.730 ;
        RECT 1409.080 37.410 1409.340 37.730 ;
        RECT 692.460 2.400 692.600 37.410 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.910 1687.320 1359.230 1687.380 ;
        RECT 1659.290 1687.320 1659.610 1687.380 ;
        RECT 1358.910 1687.180 1659.610 1687.320 ;
        RECT 1358.910 1687.120 1359.230 1687.180 ;
        RECT 1659.290 1687.120 1659.610 1687.180 ;
        RECT 1352.470 19.280 1352.790 19.340 ;
        RECT 1358.910 19.280 1359.230 19.340 ;
        RECT 1352.470 19.140 1359.230 19.280 ;
        RECT 1352.470 19.080 1352.790 19.140 ;
        RECT 1358.910 19.080 1359.230 19.140 ;
      LAYER via ;
        RECT 1358.940 1687.120 1359.200 1687.380 ;
        RECT 1659.320 1687.120 1659.580 1687.380 ;
        RECT 1352.500 19.080 1352.760 19.340 ;
        RECT 1358.940 19.080 1359.200 19.340 ;
      LAYER met2 ;
        RECT 1659.245 1700.000 1659.525 1704.000 ;
        RECT 1659.380 1687.410 1659.520 1700.000 ;
        RECT 1358.940 1687.090 1359.200 1687.410 ;
        RECT 1659.320 1687.090 1659.580 1687.410 ;
        RECT 1359.000 19.370 1359.140 1687.090 ;
        RECT 1352.500 19.050 1352.760 19.370 ;
        RECT 1358.940 19.050 1359.200 19.370 ;
        RECT 1352.560 2.400 1352.700 19.050 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1372.710 1687.660 1373.030 1687.720 ;
        RECT 1666.190 1687.660 1666.510 1687.720 ;
        RECT 1372.710 1687.520 1666.510 1687.660 ;
        RECT 1372.710 1687.460 1373.030 1687.520 ;
        RECT 1666.190 1687.460 1666.510 1687.520 ;
        RECT 1370.410 20.640 1370.730 20.700 ;
        RECT 1372.710 20.640 1373.030 20.700 ;
        RECT 1370.410 20.500 1373.030 20.640 ;
        RECT 1370.410 20.440 1370.730 20.500 ;
        RECT 1372.710 20.440 1373.030 20.500 ;
      LAYER via ;
        RECT 1372.740 1687.460 1373.000 1687.720 ;
        RECT 1666.220 1687.460 1666.480 1687.720 ;
        RECT 1370.440 20.440 1370.700 20.700 ;
        RECT 1372.740 20.440 1373.000 20.700 ;
      LAYER met2 ;
        RECT 1666.145 1700.000 1666.425 1704.000 ;
        RECT 1666.280 1687.750 1666.420 1700.000 ;
        RECT 1372.740 1687.430 1373.000 1687.750 ;
        RECT 1666.220 1687.430 1666.480 1687.750 ;
        RECT 1372.800 20.730 1372.940 1687.430 ;
        RECT 1370.440 20.410 1370.700 20.730 ;
        RECT 1372.740 20.410 1373.000 20.730 ;
        RECT 1370.500 2.400 1370.640 20.410 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1486.865 1686.485 1487.035 1689.715 ;
      LAYER mcon ;
        RECT 1486.865 1689.545 1487.035 1689.715 ;
      LAYER met1 ;
        RECT 1486.805 1689.700 1487.095 1689.745 ;
        RECT 1672.630 1689.700 1672.950 1689.760 ;
        RECT 1486.805 1689.560 1672.950 1689.700 ;
        RECT 1486.805 1689.515 1487.095 1689.560 ;
        RECT 1672.630 1689.500 1672.950 1689.560 ;
        RECT 1440.330 1686.640 1440.650 1686.700 ;
        RECT 1486.805 1686.640 1487.095 1686.685 ;
        RECT 1440.330 1686.500 1487.095 1686.640 ;
        RECT 1440.330 1686.440 1440.650 1686.500 ;
        RECT 1486.805 1686.455 1487.095 1686.500 ;
        RECT 1388.350 18.260 1388.670 18.320 ;
        RECT 1438.490 18.260 1438.810 18.320 ;
        RECT 1388.350 18.120 1438.810 18.260 ;
        RECT 1388.350 18.060 1388.670 18.120 ;
        RECT 1438.490 18.060 1438.810 18.120 ;
      LAYER via ;
        RECT 1672.660 1689.500 1672.920 1689.760 ;
        RECT 1440.360 1686.440 1440.620 1686.700 ;
        RECT 1388.380 18.060 1388.640 18.320 ;
        RECT 1438.520 18.060 1438.780 18.320 ;
      LAYER met2 ;
        RECT 1672.585 1700.000 1672.865 1704.000 ;
        RECT 1672.720 1689.790 1672.860 1700.000 ;
        RECT 1672.660 1689.470 1672.920 1689.790 ;
        RECT 1440.360 1686.410 1440.620 1686.730 ;
        RECT 1440.420 1671.170 1440.560 1686.410 ;
        RECT 1438.580 1671.030 1440.560 1671.170 ;
        RECT 1438.580 18.350 1438.720 1671.030 ;
        RECT 1388.380 18.030 1388.640 18.350 ;
        RECT 1438.520 18.030 1438.780 18.350 ;
        RECT 1388.440 2.400 1388.580 18.030 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1470.305 1647.045 1470.475 1690.055 ;
        RECT 1423.385 19.465 1423.555 20.655 ;
      LAYER mcon ;
        RECT 1470.305 1689.885 1470.475 1690.055 ;
        RECT 1423.385 20.485 1423.555 20.655 ;
      LAYER met1 ;
        RECT 1470.245 1690.040 1470.535 1690.085 ;
        RECT 1679.530 1690.040 1679.850 1690.100 ;
        RECT 1470.245 1689.900 1679.850 1690.040 ;
        RECT 1470.245 1689.855 1470.535 1689.900 ;
        RECT 1679.530 1689.840 1679.850 1689.900 ;
        RECT 1452.290 1647.200 1452.610 1647.260 ;
        RECT 1470.245 1647.200 1470.535 1647.245 ;
        RECT 1452.290 1647.060 1470.535 1647.200 ;
        RECT 1452.290 1647.000 1452.610 1647.060 ;
        RECT 1470.245 1647.015 1470.535 1647.060 ;
        RECT 1406.290 20.640 1406.610 20.700 ;
        RECT 1423.325 20.640 1423.615 20.685 ;
        RECT 1406.290 20.500 1423.615 20.640 ;
        RECT 1406.290 20.440 1406.610 20.500 ;
        RECT 1423.325 20.455 1423.615 20.500 ;
        RECT 1423.325 19.620 1423.615 19.665 ;
        RECT 1452.290 19.620 1452.610 19.680 ;
        RECT 1423.325 19.480 1452.610 19.620 ;
        RECT 1423.325 19.435 1423.615 19.480 ;
        RECT 1452.290 19.420 1452.610 19.480 ;
      LAYER via ;
        RECT 1679.560 1689.840 1679.820 1690.100 ;
        RECT 1452.320 1647.000 1452.580 1647.260 ;
        RECT 1406.320 20.440 1406.580 20.700 ;
        RECT 1452.320 19.420 1452.580 19.680 ;
      LAYER met2 ;
        RECT 1679.485 1700.000 1679.765 1704.000 ;
        RECT 1679.620 1690.130 1679.760 1700.000 ;
        RECT 1679.560 1689.810 1679.820 1690.130 ;
        RECT 1452.320 1646.970 1452.580 1647.290 ;
        RECT 1406.320 20.410 1406.580 20.730 ;
        RECT 1406.380 2.400 1406.520 20.410 ;
        RECT 1452.380 19.710 1452.520 1646.970 ;
        RECT 1452.320 19.390 1452.580 19.710 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1427.910 1689.020 1428.230 1689.080 ;
        RECT 1686.430 1689.020 1686.750 1689.080 ;
        RECT 1427.910 1688.880 1686.750 1689.020 ;
        RECT 1427.910 1688.820 1428.230 1688.880 ;
        RECT 1686.430 1688.820 1686.750 1688.880 ;
        RECT 1423.770 20.640 1424.090 20.700 ;
        RECT 1427.910 20.640 1428.230 20.700 ;
        RECT 1423.770 20.500 1428.230 20.640 ;
        RECT 1423.770 20.440 1424.090 20.500 ;
        RECT 1427.910 20.440 1428.230 20.500 ;
      LAYER via ;
        RECT 1427.940 1688.820 1428.200 1689.080 ;
        RECT 1686.460 1688.820 1686.720 1689.080 ;
        RECT 1423.800 20.440 1424.060 20.700 ;
        RECT 1427.940 20.440 1428.200 20.700 ;
      LAYER met2 ;
        RECT 1686.385 1700.000 1686.665 1704.000 ;
        RECT 1686.520 1689.110 1686.660 1700.000 ;
        RECT 1427.940 1688.790 1428.200 1689.110 ;
        RECT 1686.460 1688.790 1686.720 1689.110 ;
        RECT 1428.000 20.730 1428.140 1688.790 ;
        RECT 1423.800 20.410 1424.060 20.730 ;
        RECT 1427.940 20.410 1428.200 20.730 ;
        RECT 1423.860 2.400 1424.000 20.410 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 18.260 1442.030 18.320 ;
        RECT 1691.490 18.260 1691.810 18.320 ;
        RECT 1441.710 18.120 1691.810 18.260 ;
        RECT 1441.710 18.060 1442.030 18.120 ;
        RECT 1691.490 18.060 1691.810 18.120 ;
      LAYER via ;
        RECT 1441.740 18.060 1442.000 18.320 ;
        RECT 1691.520 18.060 1691.780 18.320 ;
      LAYER met2 ;
        RECT 1692.825 1700.410 1693.105 1704.000 ;
        RECT 1691.580 1700.270 1693.105 1700.410 ;
        RECT 1691.580 18.350 1691.720 1700.270 ;
        RECT 1692.825 1700.000 1693.105 1700.270 ;
        RECT 1441.740 18.030 1442.000 18.350 ;
        RECT 1691.520 18.030 1691.780 18.350 ;
        RECT 1441.800 2.400 1441.940 18.030 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1510.785 1689.205 1510.955 1690.395 ;
      LAYER mcon ;
        RECT 1510.785 1690.225 1510.955 1690.395 ;
      LAYER met1 ;
        RECT 1462.410 1690.380 1462.730 1690.440 ;
        RECT 1510.725 1690.380 1511.015 1690.425 ;
        RECT 1462.410 1690.240 1511.015 1690.380 ;
        RECT 1462.410 1690.180 1462.730 1690.240 ;
        RECT 1510.725 1690.195 1511.015 1690.240 ;
        RECT 1510.725 1689.360 1511.015 1689.405 ;
        RECT 1699.770 1689.360 1700.090 1689.420 ;
        RECT 1510.725 1689.220 1700.090 1689.360 ;
        RECT 1510.725 1689.175 1511.015 1689.220 ;
        RECT 1699.770 1689.160 1700.090 1689.220 ;
        RECT 1459.650 20.640 1459.970 20.700 ;
        RECT 1462.410 20.640 1462.730 20.700 ;
        RECT 1459.650 20.500 1462.730 20.640 ;
        RECT 1459.650 20.440 1459.970 20.500 ;
        RECT 1462.410 20.440 1462.730 20.500 ;
      LAYER via ;
        RECT 1462.440 1690.180 1462.700 1690.440 ;
        RECT 1699.800 1689.160 1700.060 1689.420 ;
        RECT 1459.680 20.440 1459.940 20.700 ;
        RECT 1462.440 20.440 1462.700 20.700 ;
      LAYER met2 ;
        RECT 1699.725 1700.000 1700.005 1704.000 ;
        RECT 1462.440 1690.150 1462.700 1690.470 ;
        RECT 1462.500 20.730 1462.640 1690.150 ;
        RECT 1699.860 1689.450 1700.000 1700.000 ;
        RECT 1699.800 1689.130 1700.060 1689.450 ;
        RECT 1459.680 20.410 1459.940 20.730 ;
        RECT 1462.440 20.410 1462.700 20.730 ;
        RECT 1459.740 2.400 1459.880 20.410 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1630.845 1685.805 1631.935 1685.975 ;
      LAYER mcon ;
        RECT 1631.765 1685.805 1631.935 1685.975 ;
      LAYER met1 ;
        RECT 1563.610 1685.960 1563.930 1686.020 ;
        RECT 1630.785 1685.960 1631.075 1686.005 ;
        RECT 1563.610 1685.820 1631.075 1685.960 ;
        RECT 1563.610 1685.760 1563.930 1685.820 ;
        RECT 1630.785 1685.775 1631.075 1685.820 ;
        RECT 1631.705 1685.960 1631.995 1686.005 ;
        RECT 1706.670 1685.960 1706.990 1686.020 ;
        RECT 1631.705 1685.820 1706.990 1685.960 ;
        RECT 1631.705 1685.775 1631.995 1685.820 ;
        RECT 1706.670 1685.760 1706.990 1685.820 ;
        RECT 1477.590 15.540 1477.910 15.600 ;
        RECT 1562.690 15.540 1563.010 15.600 ;
        RECT 1477.590 15.400 1563.010 15.540 ;
        RECT 1477.590 15.340 1477.910 15.400 ;
        RECT 1562.690 15.340 1563.010 15.400 ;
      LAYER via ;
        RECT 1563.640 1685.760 1563.900 1686.020 ;
        RECT 1706.700 1685.760 1706.960 1686.020 ;
        RECT 1477.620 15.340 1477.880 15.600 ;
        RECT 1562.720 15.340 1562.980 15.600 ;
      LAYER met2 ;
        RECT 1706.625 1700.000 1706.905 1704.000 ;
        RECT 1706.760 1686.050 1706.900 1700.000 ;
        RECT 1563.640 1685.730 1563.900 1686.050 ;
        RECT 1706.700 1685.730 1706.960 1686.050 ;
        RECT 1563.700 1671.170 1563.840 1685.730 ;
        RECT 1562.780 1671.030 1563.840 1671.170 ;
        RECT 1562.780 15.630 1562.920 1671.030 ;
        RECT 1477.620 15.310 1477.880 15.630 ;
        RECT 1562.720 15.310 1562.980 15.630 ;
        RECT 1477.680 2.400 1477.820 15.310 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1607.845 16.745 1608.015 19.975 ;
      LAYER mcon ;
        RECT 1607.845 19.805 1608.015 19.975 ;
      LAYER met1 ;
        RECT 1639.050 1683.920 1639.370 1683.980 ;
        RECT 1713.110 1683.920 1713.430 1683.980 ;
        RECT 1639.050 1683.780 1713.430 1683.920 ;
        RECT 1639.050 1683.720 1639.370 1683.780 ;
        RECT 1713.110 1683.720 1713.430 1683.780 ;
        RECT 1607.785 19.960 1608.075 20.005 ;
        RECT 1639.050 19.960 1639.370 20.020 ;
        RECT 1607.785 19.820 1639.370 19.960 ;
        RECT 1607.785 19.775 1608.075 19.820 ;
        RECT 1639.050 19.760 1639.370 19.820 ;
        RECT 1546.220 17.100 1559.700 17.240 ;
        RECT 1495.530 16.560 1495.850 16.620 ;
        RECT 1546.220 16.560 1546.360 17.100 ;
        RECT 1559.560 16.900 1559.700 17.100 ;
        RECT 1607.785 16.900 1608.075 16.945 ;
        RECT 1559.560 16.760 1608.075 16.900 ;
        RECT 1607.785 16.715 1608.075 16.760 ;
        RECT 1495.530 16.420 1546.360 16.560 ;
        RECT 1495.530 16.360 1495.850 16.420 ;
      LAYER via ;
        RECT 1639.080 1683.720 1639.340 1683.980 ;
        RECT 1713.140 1683.720 1713.400 1683.980 ;
        RECT 1639.080 19.760 1639.340 20.020 ;
        RECT 1495.560 16.360 1495.820 16.620 ;
      LAYER met2 ;
        RECT 1713.065 1700.000 1713.345 1704.000 ;
        RECT 1713.200 1684.010 1713.340 1700.000 ;
        RECT 1639.080 1683.690 1639.340 1684.010 ;
        RECT 1713.140 1683.690 1713.400 1684.010 ;
        RECT 1639.140 20.050 1639.280 1683.690 ;
        RECT 1639.080 19.730 1639.340 20.050 ;
        RECT 1495.560 16.330 1495.820 16.650 ;
        RECT 1495.620 2.400 1495.760 16.330 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1689.725 1686.485 1689.895 1689.035 ;
      LAYER mcon ;
        RECT 1689.725 1688.865 1689.895 1689.035 ;
      LAYER met1 ;
        RECT 1689.665 1689.020 1689.955 1689.065 ;
        RECT 1720.010 1689.020 1720.330 1689.080 ;
        RECT 1689.665 1688.880 1720.330 1689.020 ;
        RECT 1689.665 1688.835 1689.955 1688.880 ;
        RECT 1720.010 1688.820 1720.330 1688.880 ;
        RECT 1517.610 1686.640 1517.930 1686.700 ;
        RECT 1689.665 1686.640 1689.955 1686.685 ;
        RECT 1517.610 1686.500 1689.955 1686.640 ;
        RECT 1517.610 1686.440 1517.930 1686.500 ;
        RECT 1689.665 1686.455 1689.955 1686.500 ;
        RECT 1513.010 14.520 1513.330 14.580 ;
        RECT 1517.610 14.520 1517.930 14.580 ;
        RECT 1513.010 14.380 1517.930 14.520 ;
        RECT 1513.010 14.320 1513.330 14.380 ;
        RECT 1517.610 14.320 1517.930 14.380 ;
      LAYER via ;
        RECT 1720.040 1688.820 1720.300 1689.080 ;
        RECT 1517.640 1686.440 1517.900 1686.700 ;
        RECT 1513.040 14.320 1513.300 14.580 ;
        RECT 1517.640 14.320 1517.900 14.580 ;
      LAYER met2 ;
        RECT 1719.965 1700.000 1720.245 1704.000 ;
        RECT 1720.100 1689.110 1720.240 1700.000 ;
        RECT 1720.040 1688.790 1720.300 1689.110 ;
        RECT 1517.640 1686.410 1517.900 1686.730 ;
        RECT 1517.700 14.610 1517.840 1686.410 ;
        RECT 1513.040 14.290 1513.300 14.610 ;
        RECT 1517.640 14.290 1517.900 14.610 ;
        RECT 1513.100 2.400 1513.240 14.290 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 710.310 37.300 710.630 37.360 ;
        RECT 1415.950 37.300 1416.270 37.360 ;
        RECT 710.310 37.160 1416.270 37.300 ;
        RECT 710.310 37.100 710.630 37.160 ;
        RECT 1415.950 37.100 1416.270 37.160 ;
      LAYER via ;
        RECT 710.340 37.100 710.600 37.360 ;
        RECT 1415.980 37.100 1416.240 37.360 ;
      LAYER met2 ;
        RECT 1416.825 1700.410 1417.105 1704.000 ;
        RECT 1416.040 1700.270 1417.105 1700.410 ;
        RECT 1416.040 37.390 1416.180 1700.270 ;
        RECT 1416.825 1700.000 1417.105 1700.270 ;
        RECT 710.340 37.070 710.600 37.390 ;
        RECT 1415.980 37.070 1416.240 37.390 ;
        RECT 710.400 2.400 710.540 37.070 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1631.765 14.705 1631.935 16.235 ;
      LAYER mcon ;
        RECT 1631.765 16.065 1631.935 16.235 ;
      LAYER met1 ;
        RECT 1673.550 1689.700 1673.870 1689.760 ;
        RECT 1726.910 1689.700 1727.230 1689.760 ;
        RECT 1673.550 1689.560 1727.230 1689.700 ;
        RECT 1673.550 1689.500 1673.870 1689.560 ;
        RECT 1726.910 1689.500 1727.230 1689.560 ;
        RECT 1530.950 16.220 1531.270 16.280 ;
        RECT 1631.705 16.220 1631.995 16.265 ;
        RECT 1530.950 16.080 1631.995 16.220 ;
        RECT 1530.950 16.020 1531.270 16.080 ;
        RECT 1631.705 16.035 1631.995 16.080 ;
        RECT 1631.705 14.860 1631.995 14.905 ;
        RECT 1673.090 14.860 1673.410 14.920 ;
        RECT 1631.705 14.720 1673.410 14.860 ;
        RECT 1631.705 14.675 1631.995 14.720 ;
        RECT 1673.090 14.660 1673.410 14.720 ;
      LAYER via ;
        RECT 1673.580 1689.500 1673.840 1689.760 ;
        RECT 1726.940 1689.500 1727.200 1689.760 ;
        RECT 1530.980 16.020 1531.240 16.280 ;
        RECT 1673.120 14.660 1673.380 14.920 ;
      LAYER met2 ;
        RECT 1726.865 1700.000 1727.145 1704.000 ;
        RECT 1727.000 1689.790 1727.140 1700.000 ;
        RECT 1673.580 1689.470 1673.840 1689.790 ;
        RECT 1726.940 1689.470 1727.200 1689.790 ;
        RECT 1530.980 15.990 1531.240 16.310 ;
        RECT 1531.040 2.400 1531.180 15.990 ;
        RECT 1673.640 15.370 1673.780 1689.470 ;
        RECT 1673.180 15.230 1673.780 15.370 ;
        RECT 1673.180 14.950 1673.320 15.230 ;
        RECT 1673.120 14.630 1673.380 14.950 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1733.350 1685.620 1733.670 1685.680 ;
        RECT 1715.960 1685.480 1733.670 1685.620 ;
        RECT 1715.960 1685.280 1716.100 1685.480 ;
        RECT 1733.350 1685.420 1733.670 1685.480 ;
        RECT 1709.520 1685.140 1716.100 1685.280 ;
        RECT 1693.790 1684.260 1694.110 1684.320 ;
        RECT 1709.520 1684.260 1709.660 1685.140 ;
        RECT 1693.790 1684.120 1709.660 1684.260 ;
        RECT 1693.790 1684.060 1694.110 1684.120 ;
        RECT 1548.890 16.560 1549.210 16.620 ;
        RECT 1693.790 16.560 1694.110 16.620 ;
        RECT 1548.890 16.420 1694.110 16.560 ;
        RECT 1548.890 16.360 1549.210 16.420 ;
        RECT 1693.790 16.360 1694.110 16.420 ;
      LAYER via ;
        RECT 1733.380 1685.420 1733.640 1685.680 ;
        RECT 1693.820 1684.060 1694.080 1684.320 ;
        RECT 1548.920 16.360 1549.180 16.620 ;
        RECT 1693.820 16.360 1694.080 16.620 ;
      LAYER met2 ;
        RECT 1733.305 1700.000 1733.585 1704.000 ;
        RECT 1733.440 1685.710 1733.580 1700.000 ;
        RECT 1733.380 1685.390 1733.640 1685.710 ;
        RECT 1693.820 1684.030 1694.080 1684.350 ;
        RECT 1693.880 16.650 1694.020 1684.030 ;
        RECT 1548.920 16.330 1549.180 16.650 ;
        RECT 1693.820 16.330 1694.080 16.650 ;
        RECT 1548.980 2.400 1549.120 16.330 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1709.890 1684.940 1710.210 1685.000 ;
        RECT 1740.250 1684.940 1740.570 1685.000 ;
        RECT 1709.890 1684.800 1740.570 1684.940 ;
        RECT 1709.890 1684.740 1710.210 1684.800 ;
        RECT 1740.250 1684.740 1740.570 1684.800 ;
        RECT 1707.590 15.540 1707.910 15.600 ;
        RECT 1632.240 15.400 1707.910 15.540 ;
        RECT 1566.830 15.200 1567.150 15.260 ;
        RECT 1632.240 15.200 1632.380 15.400 ;
        RECT 1707.590 15.340 1707.910 15.400 ;
        RECT 1566.830 15.060 1632.380 15.200 ;
        RECT 1566.830 15.000 1567.150 15.060 ;
      LAYER via ;
        RECT 1709.920 1684.740 1710.180 1685.000 ;
        RECT 1740.280 1684.740 1740.540 1685.000 ;
        RECT 1566.860 15.000 1567.120 15.260 ;
        RECT 1707.620 15.340 1707.880 15.600 ;
      LAYER met2 ;
        RECT 1740.205 1700.000 1740.485 1704.000 ;
        RECT 1740.340 1685.030 1740.480 1700.000 ;
        RECT 1709.920 1684.710 1710.180 1685.030 ;
        RECT 1740.280 1684.710 1740.540 1685.030 ;
        RECT 1709.980 1677.290 1710.120 1684.710 ;
        RECT 1707.680 1677.150 1710.120 1677.290 ;
        RECT 1707.680 15.630 1707.820 1677.150 ;
        RECT 1707.620 15.310 1707.880 15.630 ;
        RECT 1566.860 14.970 1567.120 15.290 ;
        RECT 1566.920 2.400 1567.060 14.970 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1723.230 1684.260 1723.550 1684.320 ;
        RECT 1746.690 1684.260 1747.010 1684.320 ;
        RECT 1723.230 1684.120 1747.010 1684.260 ;
        RECT 1723.230 1684.060 1723.550 1684.120 ;
        RECT 1746.690 1684.060 1747.010 1684.120 ;
        RECT 1584.770 19.280 1585.090 19.340 ;
        RECT 1720.930 19.280 1721.250 19.340 ;
        RECT 1584.770 19.140 1721.250 19.280 ;
        RECT 1584.770 19.080 1585.090 19.140 ;
        RECT 1720.930 19.080 1721.250 19.140 ;
      LAYER via ;
        RECT 1723.260 1684.060 1723.520 1684.320 ;
        RECT 1746.720 1684.060 1746.980 1684.320 ;
        RECT 1584.800 19.080 1585.060 19.340 ;
        RECT 1720.960 19.080 1721.220 19.340 ;
      LAYER met2 ;
        RECT 1746.645 1700.000 1746.925 1704.000 ;
        RECT 1746.780 1684.350 1746.920 1700.000 ;
        RECT 1723.260 1684.030 1723.520 1684.350 ;
        RECT 1746.720 1684.030 1746.980 1684.350 ;
        RECT 1723.320 1677.290 1723.460 1684.030 ;
        RECT 1721.480 1677.150 1723.460 1677.290 ;
        RECT 1721.480 21.490 1721.620 1677.150 ;
        RECT 1721.020 21.350 1721.620 21.490 ;
        RECT 1721.020 19.370 1721.160 21.350 ;
        RECT 1584.800 19.050 1585.060 19.370 ;
        RECT 1720.960 19.050 1721.220 19.370 ;
        RECT 1584.860 2.400 1585.000 19.050 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1753.590 1686.300 1753.910 1686.360 ;
        RECT 1631.320 1686.160 1753.910 1686.300 ;
        RECT 1607.310 1685.620 1607.630 1685.680 ;
        RECT 1631.320 1685.620 1631.460 1686.160 ;
        RECT 1753.590 1686.100 1753.910 1686.160 ;
        RECT 1607.310 1685.480 1631.460 1685.620 ;
        RECT 1607.310 1685.420 1607.630 1685.480 ;
        RECT 1602.250 19.960 1602.570 20.020 ;
        RECT 1607.310 19.960 1607.630 20.020 ;
        RECT 1602.250 19.820 1607.630 19.960 ;
        RECT 1602.250 19.760 1602.570 19.820 ;
        RECT 1607.310 19.760 1607.630 19.820 ;
      LAYER via ;
        RECT 1607.340 1685.420 1607.600 1685.680 ;
        RECT 1753.620 1686.100 1753.880 1686.360 ;
        RECT 1602.280 19.760 1602.540 20.020 ;
        RECT 1607.340 19.760 1607.600 20.020 ;
      LAYER met2 ;
        RECT 1753.545 1700.000 1753.825 1704.000 ;
        RECT 1753.680 1686.390 1753.820 1700.000 ;
        RECT 1753.620 1686.070 1753.880 1686.390 ;
        RECT 1607.340 1685.390 1607.600 1685.710 ;
        RECT 1607.400 20.050 1607.540 1685.390 ;
        RECT 1602.280 19.730 1602.540 20.050 ;
        RECT 1607.340 19.730 1607.600 20.050 ;
        RECT 1602.340 2.400 1602.480 19.730 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1722.845 17.765 1723.015 19.635 ;
      LAYER mcon ;
        RECT 1722.845 19.465 1723.015 19.635 ;
      LAYER met1 ;
        RECT 1722.785 19.620 1723.075 19.665 ;
        RECT 1760.490 19.620 1760.810 19.680 ;
        RECT 1722.785 19.480 1760.810 19.620 ;
        RECT 1722.785 19.435 1723.075 19.480 ;
        RECT 1760.490 19.420 1760.810 19.480 ;
        RECT 1620.190 17.920 1620.510 17.980 ;
        RECT 1722.785 17.920 1723.075 17.965 ;
        RECT 1620.190 17.780 1723.075 17.920 ;
        RECT 1620.190 17.720 1620.510 17.780 ;
        RECT 1722.785 17.735 1723.075 17.780 ;
      LAYER via ;
        RECT 1760.520 19.420 1760.780 19.680 ;
        RECT 1620.220 17.720 1620.480 17.980 ;
      LAYER met2 ;
        RECT 1760.445 1700.000 1760.725 1704.000 ;
        RECT 1760.580 19.710 1760.720 1700.000 ;
        RECT 1760.520 19.390 1760.780 19.710 ;
        RECT 1620.220 17.690 1620.480 18.010 ;
        RECT 1620.280 2.400 1620.420 17.690 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1762.790 1688.680 1763.110 1688.740 ;
        RECT 1766.930 1688.680 1767.250 1688.740 ;
        RECT 1762.790 1688.540 1767.250 1688.680 ;
        RECT 1762.790 1688.480 1763.110 1688.540 ;
        RECT 1766.930 1688.480 1767.250 1688.540 ;
        RECT 1638.130 15.880 1638.450 15.940 ;
        RECT 1762.330 15.880 1762.650 15.940 ;
        RECT 1638.130 15.740 1762.650 15.880 ;
        RECT 1638.130 15.680 1638.450 15.740 ;
        RECT 1762.330 15.680 1762.650 15.740 ;
      LAYER via ;
        RECT 1762.820 1688.480 1763.080 1688.740 ;
        RECT 1766.960 1688.480 1767.220 1688.740 ;
        RECT 1638.160 15.680 1638.420 15.940 ;
        RECT 1762.360 15.680 1762.620 15.940 ;
      LAYER met2 ;
        RECT 1766.885 1700.000 1767.165 1704.000 ;
        RECT 1767.020 1688.770 1767.160 1700.000 ;
        RECT 1762.820 1688.450 1763.080 1688.770 ;
        RECT 1766.960 1688.450 1767.220 1688.770 ;
        RECT 1762.880 18.090 1763.020 1688.450 ;
        RECT 1762.420 17.950 1763.020 18.090 ;
        RECT 1762.420 15.970 1762.560 17.950 ;
        RECT 1638.160 15.650 1638.420 15.970 ;
        RECT 1762.360 15.650 1762.620 15.970 ;
        RECT 1638.220 2.400 1638.360 15.650 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1728.290 1685.960 1728.610 1686.020 ;
        RECT 1773.830 1685.960 1774.150 1686.020 ;
        RECT 1728.290 1685.820 1774.150 1685.960 ;
        RECT 1728.290 1685.760 1728.610 1685.820 ;
        RECT 1773.830 1685.760 1774.150 1685.820 ;
        RECT 1656.070 14.520 1656.390 14.580 ;
        RECT 1728.290 14.520 1728.610 14.580 ;
        RECT 1656.070 14.380 1728.610 14.520 ;
        RECT 1656.070 14.320 1656.390 14.380 ;
        RECT 1728.290 14.320 1728.610 14.380 ;
      LAYER via ;
        RECT 1728.320 1685.760 1728.580 1686.020 ;
        RECT 1773.860 1685.760 1774.120 1686.020 ;
        RECT 1656.100 14.320 1656.360 14.580 ;
        RECT 1728.320 14.320 1728.580 14.580 ;
      LAYER met2 ;
        RECT 1773.785 1700.000 1774.065 1704.000 ;
        RECT 1773.920 1686.050 1774.060 1700.000 ;
        RECT 1728.320 1685.730 1728.580 1686.050 ;
        RECT 1773.860 1685.730 1774.120 1686.050 ;
        RECT 1728.380 14.610 1728.520 1685.730 ;
        RECT 1656.100 14.290 1656.360 14.610 ;
        RECT 1728.320 14.290 1728.580 14.610 ;
        RECT 1656.160 2.400 1656.300 14.290 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1673.550 14.860 1673.870 14.920 ;
        RECT 1782.110 14.860 1782.430 14.920 ;
        RECT 1673.550 14.720 1782.430 14.860 ;
        RECT 1673.550 14.660 1673.870 14.720 ;
        RECT 1782.110 14.660 1782.430 14.720 ;
      LAYER via ;
        RECT 1673.580 14.660 1673.840 14.920 ;
        RECT 1782.140 14.660 1782.400 14.920 ;
      LAYER met2 ;
        RECT 1780.685 1700.410 1780.965 1704.000 ;
        RECT 1780.685 1700.270 1782.340 1700.410 ;
        RECT 1780.685 1700.000 1780.965 1700.270 ;
        RECT 1782.200 14.950 1782.340 1700.270 ;
        RECT 1673.580 14.630 1673.840 14.950 ;
        RECT 1782.140 14.630 1782.400 14.950 ;
        RECT 1673.640 2.400 1673.780 14.630 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1765.165 1687.505 1765.335 1690.395 ;
      LAYER mcon ;
        RECT 1765.165 1690.225 1765.335 1690.395 ;
      LAYER met1 ;
        RECT 1765.105 1690.380 1765.395 1690.425 ;
        RECT 1787.170 1690.380 1787.490 1690.440 ;
        RECT 1765.105 1690.240 1787.490 1690.380 ;
        RECT 1765.105 1690.195 1765.395 1690.240 ;
        RECT 1787.170 1690.180 1787.490 1690.240 ;
        RECT 1742.090 1687.660 1742.410 1687.720 ;
        RECT 1765.105 1687.660 1765.395 1687.705 ;
        RECT 1742.090 1687.520 1765.395 1687.660 ;
        RECT 1742.090 1687.460 1742.410 1687.520 ;
        RECT 1765.105 1687.475 1765.395 1687.520 ;
        RECT 1691.490 16.220 1691.810 16.280 ;
        RECT 1742.090 16.220 1742.410 16.280 ;
        RECT 1691.490 16.080 1742.410 16.220 ;
        RECT 1691.490 16.020 1691.810 16.080 ;
        RECT 1742.090 16.020 1742.410 16.080 ;
      LAYER via ;
        RECT 1787.200 1690.180 1787.460 1690.440 ;
        RECT 1742.120 1687.460 1742.380 1687.720 ;
        RECT 1691.520 16.020 1691.780 16.280 ;
        RECT 1742.120 16.020 1742.380 16.280 ;
      LAYER met2 ;
        RECT 1787.125 1700.000 1787.405 1704.000 ;
        RECT 1787.260 1690.470 1787.400 1700.000 ;
        RECT 1787.200 1690.150 1787.460 1690.470 ;
        RECT 1742.120 1687.430 1742.380 1687.750 ;
        RECT 1742.180 16.310 1742.320 1687.430 ;
        RECT 1691.520 15.990 1691.780 16.310 ;
        RECT 1742.120 15.990 1742.380 16.310 ;
        RECT 1691.580 2.400 1691.720 15.990 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 728.250 36.960 728.570 37.020 ;
        RECT 1422.850 36.960 1423.170 37.020 ;
        RECT 728.250 36.820 1423.170 36.960 ;
        RECT 728.250 36.760 728.570 36.820 ;
        RECT 1422.850 36.760 1423.170 36.820 ;
      LAYER via ;
        RECT 728.280 36.760 728.540 37.020 ;
        RECT 1422.880 36.760 1423.140 37.020 ;
      LAYER met2 ;
        RECT 1423.725 1700.410 1424.005 1704.000 ;
        RECT 1422.940 1700.270 1424.005 1700.410 ;
        RECT 1422.940 37.050 1423.080 1700.270 ;
        RECT 1423.725 1700.000 1424.005 1700.270 ;
        RECT 728.280 36.730 728.540 37.050 ;
        RECT 1422.880 36.730 1423.140 37.050 ;
        RECT 728.340 2.400 728.480 36.730 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1709.430 18.260 1709.750 18.320 ;
        RECT 1794.070 18.260 1794.390 18.320 ;
        RECT 1709.430 18.120 1794.390 18.260 ;
        RECT 1709.430 18.060 1709.750 18.120 ;
        RECT 1794.070 18.060 1794.390 18.120 ;
      LAYER via ;
        RECT 1709.460 18.060 1709.720 18.320 ;
        RECT 1794.100 18.060 1794.360 18.320 ;
      LAYER met2 ;
        RECT 1794.025 1700.000 1794.305 1704.000 ;
        RECT 1794.160 18.350 1794.300 1700.000 ;
        RECT 1709.460 18.030 1709.720 18.350 ;
        RECT 1794.100 18.030 1794.360 18.350 ;
        RECT 1709.520 2.400 1709.660 18.030 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1748.990 1690.380 1749.310 1690.440 ;
        RECT 1748.990 1690.240 1764.860 1690.380 ;
        RECT 1748.990 1690.180 1749.310 1690.240 ;
        RECT 1764.720 1690.040 1764.860 1690.240 ;
        RECT 1800.970 1690.040 1801.290 1690.100 ;
        RECT 1764.720 1689.900 1801.290 1690.040 ;
        RECT 1800.970 1689.840 1801.290 1689.900 ;
        RECT 1727.370 20.640 1727.690 20.700 ;
        RECT 1748.990 20.640 1749.310 20.700 ;
        RECT 1727.370 20.500 1749.310 20.640 ;
        RECT 1727.370 20.440 1727.690 20.500 ;
        RECT 1748.990 20.440 1749.310 20.500 ;
      LAYER via ;
        RECT 1749.020 1690.180 1749.280 1690.440 ;
        RECT 1801.000 1689.840 1801.260 1690.100 ;
        RECT 1727.400 20.440 1727.660 20.700 ;
        RECT 1749.020 20.440 1749.280 20.700 ;
      LAYER met2 ;
        RECT 1800.925 1700.000 1801.205 1704.000 ;
        RECT 1749.020 1690.150 1749.280 1690.470 ;
        RECT 1749.080 20.730 1749.220 1690.150 ;
        RECT 1801.060 1690.130 1801.200 1700.000 ;
        RECT 1801.000 1689.810 1801.260 1690.130 ;
        RECT 1727.400 20.410 1727.660 20.730 ;
        RECT 1749.020 20.410 1749.280 20.730 ;
        RECT 1727.460 2.400 1727.600 20.410 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1755.890 1686.640 1756.210 1686.700 ;
        RECT 1807.410 1686.640 1807.730 1686.700 ;
        RECT 1755.890 1686.500 1807.730 1686.640 ;
        RECT 1755.890 1686.440 1756.210 1686.500 ;
        RECT 1807.410 1686.440 1807.730 1686.500 ;
        RECT 1745.310 16.560 1745.630 16.620 ;
        RECT 1755.890 16.560 1756.210 16.620 ;
        RECT 1745.310 16.420 1756.210 16.560 ;
        RECT 1745.310 16.360 1745.630 16.420 ;
        RECT 1755.890 16.360 1756.210 16.420 ;
      LAYER via ;
        RECT 1755.920 1686.440 1756.180 1686.700 ;
        RECT 1807.440 1686.440 1807.700 1686.700 ;
        RECT 1745.340 16.360 1745.600 16.620 ;
        RECT 1755.920 16.360 1756.180 16.620 ;
      LAYER met2 ;
        RECT 1807.365 1700.000 1807.645 1704.000 ;
        RECT 1807.500 1686.730 1807.640 1700.000 ;
        RECT 1755.920 1686.410 1756.180 1686.730 ;
        RECT 1807.440 1686.410 1807.700 1686.730 ;
        RECT 1755.980 16.650 1756.120 1686.410 ;
        RECT 1745.340 16.330 1745.600 16.650 ;
        RECT 1755.920 16.330 1756.180 16.650 ;
        RECT 1745.400 2.400 1745.540 16.330 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1767.465 1687.505 1767.635 1688.695 ;
        RECT 1783.105 1687.165 1783.275 1688.695 ;
      LAYER mcon ;
        RECT 1767.465 1688.525 1767.635 1688.695 ;
        RECT 1783.105 1688.525 1783.275 1688.695 ;
      LAYER met1 ;
        RECT 1767.405 1688.680 1767.695 1688.725 ;
        RECT 1783.045 1688.680 1783.335 1688.725 ;
        RECT 1767.405 1688.540 1783.335 1688.680 ;
        RECT 1767.405 1688.495 1767.695 1688.540 ;
        RECT 1783.045 1688.495 1783.335 1688.540 ;
        RECT 1766.010 1687.660 1766.330 1687.720 ;
        RECT 1767.405 1687.660 1767.695 1687.705 ;
        RECT 1766.010 1687.520 1767.695 1687.660 ;
        RECT 1766.010 1687.460 1766.330 1687.520 ;
        RECT 1767.405 1687.475 1767.695 1687.520 ;
        RECT 1783.045 1687.320 1783.335 1687.365 ;
        RECT 1814.310 1687.320 1814.630 1687.380 ;
        RECT 1783.045 1687.180 1814.630 1687.320 ;
        RECT 1783.045 1687.135 1783.335 1687.180 ;
        RECT 1814.310 1687.120 1814.630 1687.180 ;
        RECT 1762.790 17.580 1763.110 17.640 ;
        RECT 1766.010 17.580 1766.330 17.640 ;
        RECT 1762.790 17.440 1766.330 17.580 ;
        RECT 1762.790 17.380 1763.110 17.440 ;
        RECT 1766.010 17.380 1766.330 17.440 ;
      LAYER via ;
        RECT 1766.040 1687.460 1766.300 1687.720 ;
        RECT 1814.340 1687.120 1814.600 1687.380 ;
        RECT 1762.820 17.380 1763.080 17.640 ;
        RECT 1766.040 17.380 1766.300 17.640 ;
      LAYER met2 ;
        RECT 1814.265 1700.000 1814.545 1704.000 ;
        RECT 1766.040 1687.430 1766.300 1687.750 ;
        RECT 1766.100 17.670 1766.240 1687.430 ;
        RECT 1814.400 1687.410 1814.540 1700.000 ;
        RECT 1814.340 1687.090 1814.600 1687.410 ;
        RECT 1762.820 17.350 1763.080 17.670 ;
        RECT 1766.040 17.350 1766.300 17.670 ;
        RECT 1762.880 2.400 1763.020 17.350 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1816.225 1594.005 1816.395 1642.115 ;
        RECT 1815.765 1352.605 1815.935 1400.715 ;
        RECT 1815.765 1256.045 1815.935 1304.155 ;
        RECT 1814.845 386.325 1815.015 434.775 ;
        RECT 1814.845 351.305 1815.015 385.815 ;
        RECT 1815.765 241.485 1815.935 289.595 ;
        RECT 1815.765 144.925 1815.935 193.035 ;
        RECT 1816.225 48.365 1816.395 96.475 ;
      LAYER mcon ;
        RECT 1816.225 1641.945 1816.395 1642.115 ;
        RECT 1815.765 1400.545 1815.935 1400.715 ;
        RECT 1815.765 1303.985 1815.935 1304.155 ;
        RECT 1814.845 434.605 1815.015 434.775 ;
        RECT 1814.845 385.645 1815.015 385.815 ;
        RECT 1815.765 289.425 1815.935 289.595 ;
        RECT 1815.765 192.865 1815.935 193.035 ;
        RECT 1816.225 96.305 1816.395 96.475 ;
      LAYER met1 ;
        RECT 1815.230 1700.580 1815.550 1700.640 ;
        RECT 1819.370 1700.580 1819.690 1700.640 ;
        RECT 1815.230 1700.440 1819.690 1700.580 ;
        RECT 1815.230 1700.380 1815.550 1700.440 ;
        RECT 1819.370 1700.380 1819.690 1700.440 ;
        RECT 1815.230 1690.380 1815.550 1690.440 ;
        RECT 1815.690 1690.380 1816.010 1690.440 ;
        RECT 1815.230 1690.240 1816.010 1690.380 ;
        RECT 1815.230 1690.180 1815.550 1690.240 ;
        RECT 1815.690 1690.180 1816.010 1690.240 ;
        RECT 1816.150 1642.100 1816.470 1642.160 ;
        RECT 1815.955 1641.960 1816.470 1642.100 ;
        RECT 1816.150 1641.900 1816.470 1641.960 ;
        RECT 1816.165 1594.160 1816.455 1594.205 ;
        RECT 1816.610 1594.160 1816.930 1594.220 ;
        RECT 1816.165 1594.020 1816.930 1594.160 ;
        RECT 1816.165 1593.975 1816.455 1594.020 ;
        RECT 1816.610 1593.960 1816.930 1594.020 ;
        RECT 1814.770 1545.880 1815.090 1545.940 ;
        RECT 1816.610 1545.880 1816.930 1545.940 ;
        RECT 1814.770 1545.740 1816.930 1545.880 ;
        RECT 1814.770 1545.680 1815.090 1545.740 ;
        RECT 1816.610 1545.680 1816.930 1545.740 ;
        RECT 1814.770 1510.520 1815.090 1510.580 ;
        RECT 1816.150 1510.520 1816.470 1510.580 ;
        RECT 1814.770 1510.380 1816.470 1510.520 ;
        RECT 1814.770 1510.320 1815.090 1510.380 ;
        RECT 1816.150 1510.320 1816.470 1510.380 ;
        RECT 1815.690 1400.700 1816.010 1400.760 ;
        RECT 1815.495 1400.560 1816.010 1400.700 ;
        RECT 1815.690 1400.500 1816.010 1400.560 ;
        RECT 1815.705 1352.760 1815.995 1352.805 ;
        RECT 1816.150 1352.760 1816.470 1352.820 ;
        RECT 1815.705 1352.620 1816.470 1352.760 ;
        RECT 1815.705 1352.575 1815.995 1352.620 ;
        RECT 1816.150 1352.560 1816.470 1352.620 ;
        RECT 1815.690 1304.140 1816.010 1304.200 ;
        RECT 1815.495 1304.000 1816.010 1304.140 ;
        RECT 1815.690 1303.940 1816.010 1304.000 ;
        RECT 1815.705 1256.200 1815.995 1256.245 ;
        RECT 1816.150 1256.200 1816.470 1256.260 ;
        RECT 1815.705 1256.060 1816.470 1256.200 ;
        RECT 1815.705 1256.015 1815.995 1256.060 ;
        RECT 1816.150 1256.000 1816.470 1256.060 ;
        RECT 1814.770 1159.300 1815.090 1159.360 ;
        RECT 1816.150 1159.300 1816.470 1159.360 ;
        RECT 1814.770 1159.160 1816.470 1159.300 ;
        RECT 1814.770 1159.100 1815.090 1159.160 ;
        RECT 1816.150 1159.100 1816.470 1159.160 ;
        RECT 1814.770 1062.740 1815.090 1062.800 ;
        RECT 1816.150 1062.740 1816.470 1062.800 ;
        RECT 1814.770 1062.600 1816.470 1062.740 ;
        RECT 1814.770 1062.540 1815.090 1062.600 ;
        RECT 1816.150 1062.540 1816.470 1062.600 ;
        RECT 1814.770 966.180 1815.090 966.240 ;
        RECT 1816.150 966.180 1816.470 966.240 ;
        RECT 1814.770 966.040 1816.470 966.180 ;
        RECT 1814.770 965.980 1815.090 966.040 ;
        RECT 1816.150 965.980 1816.470 966.040 ;
        RECT 1814.770 869.620 1815.090 869.680 ;
        RECT 1816.150 869.620 1816.470 869.680 ;
        RECT 1814.770 869.480 1816.470 869.620 ;
        RECT 1814.770 869.420 1815.090 869.480 ;
        RECT 1816.150 869.420 1816.470 869.480 ;
        RECT 1814.770 821.000 1815.090 821.060 ;
        RECT 1815.690 821.000 1816.010 821.060 ;
        RECT 1814.770 820.860 1816.010 821.000 ;
        RECT 1814.770 820.800 1815.090 820.860 ;
        RECT 1815.690 820.800 1816.010 820.860 ;
        RECT 1814.785 434.760 1815.075 434.805 ;
        RECT 1815.230 434.760 1815.550 434.820 ;
        RECT 1814.785 434.620 1815.550 434.760 ;
        RECT 1814.785 434.575 1815.075 434.620 ;
        RECT 1815.230 434.560 1815.550 434.620 ;
        RECT 1814.770 386.480 1815.090 386.540 ;
        RECT 1814.575 386.340 1815.090 386.480 ;
        RECT 1814.770 386.280 1815.090 386.340 ;
        RECT 1814.770 385.800 1815.090 385.860 ;
        RECT 1814.575 385.660 1815.090 385.800 ;
        RECT 1814.770 385.600 1815.090 385.660 ;
        RECT 1814.785 351.460 1815.075 351.505 ;
        RECT 1815.230 351.460 1815.550 351.520 ;
        RECT 1814.785 351.320 1815.550 351.460 ;
        RECT 1814.785 351.275 1815.075 351.320 ;
        RECT 1815.230 351.260 1815.550 351.320 ;
        RECT 1815.230 303.520 1815.550 303.580 ;
        RECT 1816.150 303.520 1816.470 303.580 ;
        RECT 1815.230 303.380 1816.470 303.520 ;
        RECT 1815.230 303.320 1815.550 303.380 ;
        RECT 1816.150 303.320 1816.470 303.380 ;
        RECT 1815.705 289.580 1815.995 289.625 ;
        RECT 1816.150 289.580 1816.470 289.640 ;
        RECT 1815.705 289.440 1816.470 289.580 ;
        RECT 1815.705 289.395 1815.995 289.440 ;
        RECT 1816.150 289.380 1816.470 289.440 ;
        RECT 1815.690 241.640 1816.010 241.700 ;
        RECT 1815.495 241.500 1816.010 241.640 ;
        RECT 1815.690 241.440 1816.010 241.500 ;
        RECT 1815.230 206.960 1815.550 207.020 ;
        RECT 1816.150 206.960 1816.470 207.020 ;
        RECT 1815.230 206.820 1816.470 206.960 ;
        RECT 1815.230 206.760 1815.550 206.820 ;
        RECT 1816.150 206.760 1816.470 206.820 ;
        RECT 1815.705 193.020 1815.995 193.065 ;
        RECT 1816.150 193.020 1816.470 193.080 ;
        RECT 1815.705 192.880 1816.470 193.020 ;
        RECT 1815.705 192.835 1815.995 192.880 ;
        RECT 1816.150 192.820 1816.470 192.880 ;
        RECT 1815.690 145.080 1816.010 145.140 ;
        RECT 1815.495 144.940 1816.010 145.080 ;
        RECT 1815.690 144.880 1816.010 144.940 ;
        RECT 1815.230 110.400 1815.550 110.460 ;
        RECT 1816.150 110.400 1816.470 110.460 ;
        RECT 1815.230 110.260 1816.470 110.400 ;
        RECT 1815.230 110.200 1815.550 110.260 ;
        RECT 1816.150 110.200 1816.470 110.260 ;
        RECT 1816.150 96.460 1816.470 96.520 ;
        RECT 1815.955 96.320 1816.470 96.460 ;
        RECT 1816.150 96.260 1816.470 96.320 ;
        RECT 1816.150 48.520 1816.470 48.580 ;
        RECT 1815.955 48.380 1816.470 48.520 ;
        RECT 1816.150 48.320 1816.470 48.380 ;
        RECT 1780.730 16.560 1781.050 16.620 ;
        RECT 1816.150 16.560 1816.470 16.620 ;
        RECT 1780.730 16.420 1816.470 16.560 ;
        RECT 1780.730 16.360 1781.050 16.420 ;
        RECT 1816.150 16.360 1816.470 16.420 ;
      LAYER via ;
        RECT 1815.260 1700.380 1815.520 1700.640 ;
        RECT 1819.400 1700.380 1819.660 1700.640 ;
        RECT 1815.260 1690.180 1815.520 1690.440 ;
        RECT 1815.720 1690.180 1815.980 1690.440 ;
        RECT 1816.180 1641.900 1816.440 1642.160 ;
        RECT 1816.640 1593.960 1816.900 1594.220 ;
        RECT 1814.800 1545.680 1815.060 1545.940 ;
        RECT 1816.640 1545.680 1816.900 1545.940 ;
        RECT 1814.800 1510.320 1815.060 1510.580 ;
        RECT 1816.180 1510.320 1816.440 1510.580 ;
        RECT 1815.720 1400.500 1815.980 1400.760 ;
        RECT 1816.180 1352.560 1816.440 1352.820 ;
        RECT 1815.720 1303.940 1815.980 1304.200 ;
        RECT 1816.180 1256.000 1816.440 1256.260 ;
        RECT 1814.800 1159.100 1815.060 1159.360 ;
        RECT 1816.180 1159.100 1816.440 1159.360 ;
        RECT 1814.800 1062.540 1815.060 1062.800 ;
        RECT 1816.180 1062.540 1816.440 1062.800 ;
        RECT 1814.800 965.980 1815.060 966.240 ;
        RECT 1816.180 965.980 1816.440 966.240 ;
        RECT 1814.800 869.420 1815.060 869.680 ;
        RECT 1816.180 869.420 1816.440 869.680 ;
        RECT 1814.800 820.800 1815.060 821.060 ;
        RECT 1815.720 820.800 1815.980 821.060 ;
        RECT 1815.260 434.560 1815.520 434.820 ;
        RECT 1814.800 386.280 1815.060 386.540 ;
        RECT 1814.800 385.600 1815.060 385.860 ;
        RECT 1815.260 351.260 1815.520 351.520 ;
        RECT 1815.260 303.320 1815.520 303.580 ;
        RECT 1816.180 303.320 1816.440 303.580 ;
        RECT 1816.180 289.380 1816.440 289.640 ;
        RECT 1815.720 241.440 1815.980 241.700 ;
        RECT 1815.260 206.760 1815.520 207.020 ;
        RECT 1816.180 206.760 1816.440 207.020 ;
        RECT 1816.180 192.820 1816.440 193.080 ;
        RECT 1815.720 144.880 1815.980 145.140 ;
        RECT 1815.260 110.200 1815.520 110.460 ;
        RECT 1816.180 110.200 1816.440 110.460 ;
        RECT 1816.180 96.260 1816.440 96.520 ;
        RECT 1816.180 48.320 1816.440 48.580 ;
        RECT 1780.760 16.360 1781.020 16.620 ;
        RECT 1816.180 16.360 1816.440 16.620 ;
      LAYER met2 ;
        RECT 1820.705 1701.090 1820.985 1704.000 ;
        RECT 1819.460 1700.950 1820.985 1701.090 ;
        RECT 1819.460 1700.670 1819.600 1700.950 ;
        RECT 1815.260 1700.350 1815.520 1700.670 ;
        RECT 1819.400 1700.350 1819.660 1700.670 ;
        RECT 1815.320 1690.470 1815.460 1700.350 ;
        RECT 1820.705 1700.000 1820.985 1700.950 ;
        RECT 1815.260 1690.150 1815.520 1690.470 ;
        RECT 1815.720 1690.150 1815.980 1690.470 ;
        RECT 1815.780 1686.980 1815.920 1690.150 ;
        RECT 1815.780 1686.840 1816.380 1686.980 ;
        RECT 1816.240 1642.190 1816.380 1686.840 ;
        RECT 1816.180 1641.870 1816.440 1642.190 ;
        RECT 1816.640 1593.930 1816.900 1594.250 ;
        RECT 1816.700 1545.970 1816.840 1593.930 ;
        RECT 1814.800 1545.650 1815.060 1545.970 ;
        RECT 1816.640 1545.650 1816.900 1545.970 ;
        RECT 1814.860 1510.610 1815.000 1545.650 ;
        RECT 1814.800 1510.290 1815.060 1510.610 ;
        RECT 1816.180 1510.290 1816.440 1510.610 ;
        RECT 1816.240 1425.010 1816.380 1510.290 ;
        RECT 1815.780 1424.870 1816.380 1425.010 ;
        RECT 1815.780 1400.790 1815.920 1424.870 ;
        RECT 1815.720 1400.470 1815.980 1400.790 ;
        RECT 1816.180 1352.530 1816.440 1352.850 ;
        RECT 1816.240 1317.570 1816.380 1352.530 ;
        RECT 1815.780 1317.430 1816.380 1317.570 ;
        RECT 1815.780 1304.230 1815.920 1317.430 ;
        RECT 1815.720 1303.910 1815.980 1304.230 ;
        RECT 1816.180 1255.970 1816.440 1256.290 ;
        RECT 1816.240 1221.010 1816.380 1255.970 ;
        RECT 1815.780 1220.870 1816.380 1221.010 ;
        RECT 1815.780 1207.525 1815.920 1220.870 ;
        RECT 1814.790 1207.155 1815.070 1207.525 ;
        RECT 1815.710 1207.155 1815.990 1207.525 ;
        RECT 1814.860 1159.390 1815.000 1207.155 ;
        RECT 1814.800 1159.070 1815.060 1159.390 ;
        RECT 1816.180 1159.070 1816.440 1159.390 ;
        RECT 1816.240 1124.450 1816.380 1159.070 ;
        RECT 1815.780 1124.310 1816.380 1124.450 ;
        RECT 1815.780 1110.965 1815.920 1124.310 ;
        RECT 1814.790 1110.595 1815.070 1110.965 ;
        RECT 1815.710 1110.595 1815.990 1110.965 ;
        RECT 1814.860 1062.830 1815.000 1110.595 ;
        RECT 1814.800 1062.510 1815.060 1062.830 ;
        RECT 1816.180 1062.510 1816.440 1062.830 ;
        RECT 1816.240 1027.890 1816.380 1062.510 ;
        RECT 1815.780 1027.750 1816.380 1027.890 ;
        RECT 1815.780 1014.405 1815.920 1027.750 ;
        RECT 1814.790 1014.035 1815.070 1014.405 ;
        RECT 1815.710 1014.035 1815.990 1014.405 ;
        RECT 1814.860 966.270 1815.000 1014.035 ;
        RECT 1814.800 965.950 1815.060 966.270 ;
        RECT 1816.180 965.950 1816.440 966.270 ;
        RECT 1816.240 931.330 1816.380 965.950 ;
        RECT 1815.780 931.190 1816.380 931.330 ;
        RECT 1815.780 917.845 1815.920 931.190 ;
        RECT 1814.790 917.475 1815.070 917.845 ;
        RECT 1815.710 917.475 1815.990 917.845 ;
        RECT 1814.860 869.710 1815.000 917.475 ;
        RECT 1814.800 869.390 1815.060 869.710 ;
        RECT 1816.180 869.390 1816.440 869.710 ;
        RECT 1816.240 834.770 1816.380 869.390 ;
        RECT 1815.780 834.630 1816.380 834.770 ;
        RECT 1815.780 821.090 1815.920 834.630 ;
        RECT 1814.800 820.770 1815.060 821.090 ;
        RECT 1815.720 820.770 1815.980 821.090 ;
        RECT 1814.860 773.005 1815.000 820.770 ;
        RECT 1814.790 772.635 1815.070 773.005 ;
        RECT 1816.170 772.635 1816.450 773.005 ;
        RECT 1816.240 738.210 1816.380 772.635 ;
        RECT 1815.780 738.070 1816.380 738.210 ;
        RECT 1815.780 700.130 1815.920 738.070 ;
        RECT 1814.860 699.990 1815.920 700.130 ;
        RECT 1814.860 676.445 1815.000 699.990 ;
        RECT 1814.790 676.075 1815.070 676.445 ;
        RECT 1816.170 676.075 1816.450 676.445 ;
        RECT 1816.240 641.650 1816.380 676.075 ;
        RECT 1815.780 641.510 1816.380 641.650 ;
        RECT 1815.780 603.570 1815.920 641.510 ;
        RECT 1814.860 603.430 1815.920 603.570 ;
        RECT 1814.860 579.885 1815.000 603.430 ;
        RECT 1814.790 579.515 1815.070 579.885 ;
        RECT 1816.170 579.515 1816.450 579.885 ;
        RECT 1816.240 545.090 1816.380 579.515 ;
        RECT 1815.780 544.950 1816.380 545.090 ;
        RECT 1815.780 507.010 1815.920 544.950 ;
        RECT 1814.860 506.870 1815.920 507.010 ;
        RECT 1814.860 483.325 1815.000 506.870 ;
        RECT 1814.790 482.955 1815.070 483.325 ;
        RECT 1816.170 482.955 1816.450 483.325 ;
        RECT 1816.240 448.530 1816.380 482.955 ;
        RECT 1815.320 448.390 1816.380 448.530 ;
        RECT 1815.320 434.850 1815.460 448.390 ;
        RECT 1815.260 434.530 1815.520 434.850 ;
        RECT 1814.800 386.250 1815.060 386.570 ;
        RECT 1814.860 385.890 1815.000 386.250 ;
        RECT 1814.800 385.570 1815.060 385.890 ;
        RECT 1815.260 351.230 1815.520 351.550 ;
        RECT 1815.320 303.610 1815.460 351.230 ;
        RECT 1815.260 303.290 1815.520 303.610 ;
        RECT 1816.180 303.290 1816.440 303.610 ;
        RECT 1816.240 289.670 1816.380 303.290 ;
        RECT 1816.180 289.350 1816.440 289.670 ;
        RECT 1815.720 241.410 1815.980 241.730 ;
        RECT 1815.780 207.130 1815.920 241.410 ;
        RECT 1815.320 207.050 1815.920 207.130 ;
        RECT 1815.260 206.990 1815.920 207.050 ;
        RECT 1815.260 206.730 1815.520 206.990 ;
        RECT 1816.180 206.730 1816.440 207.050 ;
        RECT 1816.240 193.110 1816.380 206.730 ;
        RECT 1816.180 192.790 1816.440 193.110 ;
        RECT 1815.720 144.850 1815.980 145.170 ;
        RECT 1815.780 110.570 1815.920 144.850 ;
        RECT 1815.320 110.490 1815.920 110.570 ;
        RECT 1815.260 110.430 1815.920 110.490 ;
        RECT 1815.260 110.170 1815.520 110.430 ;
        RECT 1816.180 110.170 1816.440 110.490 ;
        RECT 1816.240 96.550 1816.380 110.170 ;
        RECT 1816.180 96.230 1816.440 96.550 ;
        RECT 1816.180 48.290 1816.440 48.610 ;
        RECT 1816.240 16.650 1816.380 48.290 ;
        RECT 1780.760 16.330 1781.020 16.650 ;
        RECT 1816.180 16.330 1816.440 16.650 ;
        RECT 1780.820 2.400 1780.960 16.330 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
      LAYER via2 ;
        RECT 1814.790 1207.200 1815.070 1207.480 ;
        RECT 1815.710 1207.200 1815.990 1207.480 ;
        RECT 1814.790 1110.640 1815.070 1110.920 ;
        RECT 1815.710 1110.640 1815.990 1110.920 ;
        RECT 1814.790 1014.080 1815.070 1014.360 ;
        RECT 1815.710 1014.080 1815.990 1014.360 ;
        RECT 1814.790 917.520 1815.070 917.800 ;
        RECT 1815.710 917.520 1815.990 917.800 ;
        RECT 1814.790 772.680 1815.070 772.960 ;
        RECT 1816.170 772.680 1816.450 772.960 ;
        RECT 1814.790 676.120 1815.070 676.400 ;
        RECT 1816.170 676.120 1816.450 676.400 ;
        RECT 1814.790 579.560 1815.070 579.840 ;
        RECT 1816.170 579.560 1816.450 579.840 ;
        RECT 1814.790 483.000 1815.070 483.280 ;
        RECT 1816.170 483.000 1816.450 483.280 ;
      LAYER met3 ;
        RECT 1814.765 1207.490 1815.095 1207.505 ;
        RECT 1815.685 1207.490 1816.015 1207.505 ;
        RECT 1814.765 1207.190 1816.015 1207.490 ;
        RECT 1814.765 1207.175 1815.095 1207.190 ;
        RECT 1815.685 1207.175 1816.015 1207.190 ;
        RECT 1814.765 1110.930 1815.095 1110.945 ;
        RECT 1815.685 1110.930 1816.015 1110.945 ;
        RECT 1814.765 1110.630 1816.015 1110.930 ;
        RECT 1814.765 1110.615 1815.095 1110.630 ;
        RECT 1815.685 1110.615 1816.015 1110.630 ;
        RECT 1814.765 1014.370 1815.095 1014.385 ;
        RECT 1815.685 1014.370 1816.015 1014.385 ;
        RECT 1814.765 1014.070 1816.015 1014.370 ;
        RECT 1814.765 1014.055 1815.095 1014.070 ;
        RECT 1815.685 1014.055 1816.015 1014.070 ;
        RECT 1814.765 917.810 1815.095 917.825 ;
        RECT 1815.685 917.810 1816.015 917.825 ;
        RECT 1814.765 917.510 1816.015 917.810 ;
        RECT 1814.765 917.495 1815.095 917.510 ;
        RECT 1815.685 917.495 1816.015 917.510 ;
        RECT 1814.765 772.970 1815.095 772.985 ;
        RECT 1816.145 772.970 1816.475 772.985 ;
        RECT 1814.765 772.670 1816.475 772.970 ;
        RECT 1814.765 772.655 1815.095 772.670 ;
        RECT 1816.145 772.655 1816.475 772.670 ;
        RECT 1814.765 676.410 1815.095 676.425 ;
        RECT 1816.145 676.410 1816.475 676.425 ;
        RECT 1814.765 676.110 1816.475 676.410 ;
        RECT 1814.765 676.095 1815.095 676.110 ;
        RECT 1816.145 676.095 1816.475 676.110 ;
        RECT 1814.765 579.850 1815.095 579.865 ;
        RECT 1816.145 579.850 1816.475 579.865 ;
        RECT 1814.765 579.550 1816.475 579.850 ;
        RECT 1814.765 579.535 1815.095 579.550 ;
        RECT 1816.145 579.535 1816.475 579.550 ;
        RECT 1814.765 483.290 1815.095 483.305 ;
        RECT 1816.145 483.290 1816.475 483.305 ;
        RECT 1814.765 482.990 1816.475 483.290 ;
        RECT 1814.765 482.975 1815.095 482.990 ;
        RECT 1816.145 482.975 1816.475 482.990 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1814.385 1684.785 1814.555 1685.975 ;
      LAYER mcon ;
        RECT 1814.385 1685.805 1814.555 1685.975 ;
      LAYER met1 ;
        RECT 1814.325 1685.960 1814.615 1686.005 ;
        RECT 1827.650 1685.960 1827.970 1686.020 ;
        RECT 1814.325 1685.820 1827.970 1685.960 ;
        RECT 1814.325 1685.775 1814.615 1685.820 ;
        RECT 1827.650 1685.760 1827.970 1685.820 ;
        RECT 1800.510 1684.940 1800.830 1685.000 ;
        RECT 1814.325 1684.940 1814.615 1684.985 ;
        RECT 1800.510 1684.800 1814.615 1684.940 ;
        RECT 1800.510 1684.740 1800.830 1684.800 ;
        RECT 1814.325 1684.755 1814.615 1684.800 ;
      LAYER via ;
        RECT 1827.680 1685.760 1827.940 1686.020 ;
        RECT 1800.540 1684.740 1800.800 1685.000 ;
      LAYER met2 ;
        RECT 1827.605 1700.000 1827.885 1704.000 ;
        RECT 1827.740 1686.050 1827.880 1700.000 ;
        RECT 1827.680 1685.730 1827.940 1686.050 ;
        RECT 1800.540 1684.710 1800.800 1685.030 ;
        RECT 1800.600 3.130 1800.740 1684.710 ;
        RECT 1798.760 2.990 1800.740 3.130 ;
        RECT 1798.760 2.400 1798.900 2.990 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1821.210 1684.940 1821.530 1685.000 ;
        RECT 1834.550 1684.940 1834.870 1685.000 ;
        RECT 1821.210 1684.800 1834.870 1684.940 ;
        RECT 1821.210 1684.740 1821.530 1684.800 ;
        RECT 1834.550 1684.740 1834.870 1684.800 ;
        RECT 1816.610 17.580 1816.930 17.640 ;
        RECT 1821.210 17.580 1821.530 17.640 ;
        RECT 1816.610 17.440 1821.530 17.580 ;
        RECT 1816.610 17.380 1816.930 17.440 ;
        RECT 1821.210 17.380 1821.530 17.440 ;
      LAYER via ;
        RECT 1821.240 1684.740 1821.500 1685.000 ;
        RECT 1834.580 1684.740 1834.840 1685.000 ;
        RECT 1816.640 17.380 1816.900 17.640 ;
        RECT 1821.240 17.380 1821.500 17.640 ;
      LAYER met2 ;
        RECT 1834.505 1700.000 1834.785 1704.000 ;
        RECT 1834.640 1685.030 1834.780 1700.000 ;
        RECT 1821.240 1684.710 1821.500 1685.030 ;
        RECT 1834.580 1684.710 1834.840 1685.030 ;
        RECT 1821.300 17.670 1821.440 1684.710 ;
        RECT 1816.640 17.350 1816.900 17.670 ;
        RECT 1821.240 17.350 1821.500 17.670 ;
        RECT 1816.700 2.400 1816.840 17.350 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.010 1683.920 1835.330 1683.980 ;
        RECT 1840.990 1683.920 1841.310 1683.980 ;
        RECT 1835.010 1683.780 1841.310 1683.920 ;
        RECT 1835.010 1683.720 1835.330 1683.780 ;
        RECT 1840.990 1683.720 1841.310 1683.780 ;
      LAYER via ;
        RECT 1835.040 1683.720 1835.300 1683.980 ;
        RECT 1841.020 1683.720 1841.280 1683.980 ;
      LAYER met2 ;
        RECT 1840.945 1700.000 1841.225 1704.000 ;
        RECT 1841.080 1684.010 1841.220 1700.000 ;
        RECT 1835.040 1683.690 1835.300 1684.010 ;
        RECT 1841.020 1683.690 1841.280 1684.010 ;
        RECT 1835.100 16.050 1835.240 1683.690 ;
        RECT 1834.640 15.910 1835.240 16.050 ;
        RECT 1834.640 2.400 1834.780 15.910 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1847.845 1700.410 1848.125 1704.000 ;
        RECT 1847.845 1700.270 1849.040 1700.410 ;
        RECT 1847.845 1700.000 1848.125 1700.270 ;
        RECT 1848.900 1688.850 1849.040 1700.270 ;
        RECT 1848.900 1688.710 1850.420 1688.850 ;
        RECT 1850.280 16.730 1850.420 1688.710 ;
        RECT 1850.280 16.590 1852.260 16.730 ;
        RECT 1852.120 2.400 1852.260 16.590 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 20.640 1856.030 20.700 ;
        RECT 1869.970 20.640 1870.290 20.700 ;
        RECT 1855.710 20.500 1870.290 20.640 ;
        RECT 1855.710 20.440 1856.030 20.500 ;
        RECT 1869.970 20.440 1870.290 20.500 ;
      LAYER via ;
        RECT 1855.740 20.440 1856.000 20.700 ;
        RECT 1870.000 20.440 1870.260 20.700 ;
      LAYER met2 ;
        RECT 1854.745 1700.410 1855.025 1704.000 ;
        RECT 1854.745 1700.270 1855.940 1700.410 ;
        RECT 1854.745 1700.000 1855.025 1700.270 ;
        RECT 1855.800 20.730 1855.940 1700.270 ;
        RECT 1855.740 20.410 1856.000 20.730 ;
        RECT 1870.000 20.410 1870.260 20.730 ;
        RECT 1870.060 2.400 1870.200 20.410 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 746.190 36.620 746.510 36.680 ;
        RECT 1430.210 36.620 1430.530 36.680 ;
        RECT 746.190 36.480 1430.530 36.620 ;
        RECT 746.190 36.420 746.510 36.480 ;
        RECT 1430.210 36.420 1430.530 36.480 ;
      LAYER via ;
        RECT 746.220 36.420 746.480 36.680 ;
        RECT 1430.240 36.420 1430.500 36.680 ;
      LAYER met2 ;
        RECT 1430.165 1700.000 1430.445 1704.000 ;
        RECT 1430.300 36.710 1430.440 1700.000 ;
        RECT 746.220 36.390 746.480 36.710 ;
        RECT 1430.240 36.390 1430.500 36.710 ;
        RECT 746.280 2.400 746.420 36.390 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1861.230 1688.680 1861.550 1688.740 ;
        RECT 1866.290 1688.680 1866.610 1688.740 ;
        RECT 1861.230 1688.540 1866.610 1688.680 ;
        RECT 1861.230 1688.480 1861.550 1688.540 ;
        RECT 1866.290 1688.480 1866.610 1688.540 ;
        RECT 1866.290 17.580 1866.610 17.640 ;
        RECT 1887.910 17.580 1888.230 17.640 ;
        RECT 1866.290 17.440 1888.230 17.580 ;
        RECT 1866.290 17.380 1866.610 17.440 ;
        RECT 1887.910 17.380 1888.230 17.440 ;
      LAYER via ;
        RECT 1861.260 1688.480 1861.520 1688.740 ;
        RECT 1866.320 1688.480 1866.580 1688.740 ;
        RECT 1866.320 17.380 1866.580 17.640 ;
        RECT 1887.940 17.380 1888.200 17.640 ;
      LAYER met2 ;
        RECT 1861.185 1700.000 1861.465 1704.000 ;
        RECT 1861.320 1688.770 1861.460 1700.000 ;
        RECT 1861.260 1688.450 1861.520 1688.770 ;
        RECT 1866.320 1688.450 1866.580 1688.770 ;
        RECT 1866.380 17.670 1866.520 1688.450 ;
        RECT 1866.320 17.350 1866.580 17.670 ;
        RECT 1887.940 17.350 1888.200 17.670 ;
        RECT 1888.000 2.400 1888.140 17.350 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1868.130 1684.600 1868.450 1684.660 ;
        RECT 1873.190 1684.600 1873.510 1684.660 ;
        RECT 1868.130 1684.460 1873.510 1684.600 ;
        RECT 1868.130 1684.400 1868.450 1684.460 ;
        RECT 1873.190 1684.400 1873.510 1684.460 ;
        RECT 1873.190 18.940 1873.510 19.000 ;
        RECT 1905.850 18.940 1906.170 19.000 ;
        RECT 1873.190 18.800 1906.170 18.940 ;
        RECT 1873.190 18.740 1873.510 18.800 ;
        RECT 1905.850 18.740 1906.170 18.800 ;
      LAYER via ;
        RECT 1868.160 1684.400 1868.420 1684.660 ;
        RECT 1873.220 1684.400 1873.480 1684.660 ;
        RECT 1873.220 18.740 1873.480 19.000 ;
        RECT 1905.880 18.740 1906.140 19.000 ;
      LAYER met2 ;
        RECT 1868.085 1700.000 1868.365 1704.000 ;
        RECT 1868.220 1684.690 1868.360 1700.000 ;
        RECT 1868.160 1684.370 1868.420 1684.690 ;
        RECT 1873.220 1684.370 1873.480 1684.690 ;
        RECT 1873.280 19.030 1873.420 1684.370 ;
        RECT 1873.220 18.710 1873.480 19.030 ;
        RECT 1905.880 18.710 1906.140 19.030 ;
        RECT 1905.940 2.400 1906.080 18.710 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1875.030 1686.640 1875.350 1686.700 ;
        RECT 1907.690 1686.640 1908.010 1686.700 ;
        RECT 1875.030 1686.500 1908.010 1686.640 ;
        RECT 1875.030 1686.440 1875.350 1686.500 ;
        RECT 1907.690 1686.440 1908.010 1686.500 ;
        RECT 1907.690 20.640 1908.010 20.700 ;
        RECT 1923.330 20.640 1923.650 20.700 ;
        RECT 1907.690 20.500 1923.650 20.640 ;
        RECT 1907.690 20.440 1908.010 20.500 ;
        RECT 1923.330 20.440 1923.650 20.500 ;
      LAYER via ;
        RECT 1875.060 1686.440 1875.320 1686.700 ;
        RECT 1907.720 1686.440 1907.980 1686.700 ;
        RECT 1907.720 20.440 1907.980 20.700 ;
        RECT 1923.360 20.440 1923.620 20.700 ;
      LAYER met2 ;
        RECT 1874.985 1700.000 1875.265 1704.000 ;
        RECT 1875.120 1686.730 1875.260 1700.000 ;
        RECT 1875.060 1686.410 1875.320 1686.730 ;
        RECT 1907.720 1686.410 1907.980 1686.730 ;
        RECT 1907.780 20.730 1907.920 1686.410 ;
        RECT 1907.720 20.410 1907.980 20.730 ;
        RECT 1923.360 20.410 1923.620 20.730 ;
        RECT 1923.420 2.400 1923.560 20.410 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1909.145 1687.505 1909.315 1690.055 ;
      LAYER mcon ;
        RECT 1909.145 1689.885 1909.315 1690.055 ;
      LAYER met1 ;
        RECT 1881.470 1690.040 1881.790 1690.100 ;
        RECT 1909.085 1690.040 1909.375 1690.085 ;
        RECT 1881.470 1689.900 1909.375 1690.040 ;
        RECT 1881.470 1689.840 1881.790 1689.900 ;
        RECT 1909.085 1689.855 1909.375 1689.900 ;
        RECT 1909.085 1687.660 1909.375 1687.705 ;
        RECT 1921.490 1687.660 1921.810 1687.720 ;
        RECT 1909.085 1687.520 1921.810 1687.660 ;
        RECT 1909.085 1687.475 1909.375 1687.520 ;
        RECT 1921.490 1687.460 1921.810 1687.520 ;
        RECT 1921.490 16.220 1921.810 16.280 ;
        RECT 1941.270 16.220 1941.590 16.280 ;
        RECT 1921.490 16.080 1941.590 16.220 ;
        RECT 1921.490 16.020 1921.810 16.080 ;
        RECT 1941.270 16.020 1941.590 16.080 ;
      LAYER via ;
        RECT 1881.500 1689.840 1881.760 1690.100 ;
        RECT 1921.520 1687.460 1921.780 1687.720 ;
        RECT 1921.520 16.020 1921.780 16.280 ;
        RECT 1941.300 16.020 1941.560 16.280 ;
      LAYER met2 ;
        RECT 1881.425 1700.000 1881.705 1704.000 ;
        RECT 1881.560 1690.130 1881.700 1700.000 ;
        RECT 1881.500 1689.810 1881.760 1690.130 ;
        RECT 1921.520 1687.430 1921.780 1687.750 ;
        RECT 1921.580 16.310 1921.720 1687.430 ;
        RECT 1921.520 15.990 1921.780 16.310 ;
        RECT 1941.300 15.990 1941.560 16.310 ;
        RECT 1941.360 2.400 1941.500 15.990 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1888.370 1690.380 1888.690 1690.440 ;
        RECT 1888.370 1690.240 1917.120 1690.380 ;
        RECT 1888.370 1690.180 1888.690 1690.240 ;
        RECT 1916.980 1689.700 1917.120 1690.240 ;
        RECT 1916.980 1689.560 1930.460 1689.700 ;
        RECT 1930.320 1689.360 1930.460 1689.560 ;
        RECT 1942.190 1689.360 1942.510 1689.420 ;
        RECT 1930.320 1689.220 1942.510 1689.360 ;
        RECT 1942.190 1689.160 1942.510 1689.220 ;
        RECT 1942.190 17.580 1942.510 17.640 ;
        RECT 1959.210 17.580 1959.530 17.640 ;
        RECT 1942.190 17.440 1959.530 17.580 ;
        RECT 1942.190 17.380 1942.510 17.440 ;
        RECT 1959.210 17.380 1959.530 17.440 ;
      LAYER via ;
        RECT 1888.400 1690.180 1888.660 1690.440 ;
        RECT 1942.220 1689.160 1942.480 1689.420 ;
        RECT 1942.220 17.380 1942.480 17.640 ;
        RECT 1959.240 17.380 1959.500 17.640 ;
      LAYER met2 ;
        RECT 1888.325 1700.000 1888.605 1704.000 ;
        RECT 1888.460 1690.470 1888.600 1700.000 ;
        RECT 1888.400 1690.150 1888.660 1690.470 ;
        RECT 1942.220 1689.130 1942.480 1689.450 ;
        RECT 1942.280 17.670 1942.420 1689.130 ;
        RECT 1942.220 17.350 1942.480 17.670 ;
        RECT 1959.240 17.350 1959.500 17.670 ;
        RECT 1959.300 2.400 1959.440 17.350 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1895.270 1688.000 1895.590 1688.060 ;
        RECT 1908.150 1688.000 1908.470 1688.060 ;
        RECT 1895.270 1687.860 1908.470 1688.000 ;
        RECT 1895.270 1687.800 1895.590 1687.860 ;
        RECT 1908.150 1687.800 1908.470 1687.860 ;
        RECT 1908.150 14.860 1908.470 14.920 ;
        RECT 1977.150 14.860 1977.470 14.920 ;
        RECT 1908.150 14.720 1977.470 14.860 ;
        RECT 1908.150 14.660 1908.470 14.720 ;
        RECT 1977.150 14.660 1977.470 14.720 ;
      LAYER via ;
        RECT 1895.300 1687.800 1895.560 1688.060 ;
        RECT 1908.180 1687.800 1908.440 1688.060 ;
        RECT 1908.180 14.660 1908.440 14.920 ;
        RECT 1977.180 14.660 1977.440 14.920 ;
      LAYER met2 ;
        RECT 1895.225 1700.000 1895.505 1704.000 ;
        RECT 1895.360 1688.090 1895.500 1700.000 ;
        RECT 1895.300 1687.770 1895.560 1688.090 ;
        RECT 1908.180 1687.770 1908.440 1688.090 ;
        RECT 1908.240 14.950 1908.380 1687.770 ;
        RECT 1908.180 14.630 1908.440 14.950 ;
        RECT 1977.180 14.630 1977.440 14.950 ;
        RECT 1977.240 2.400 1977.380 14.630 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.550 1689.020 1995.870 1689.080 ;
        RECT 1980.000 1688.880 1995.870 1689.020 ;
        RECT 1901.710 1688.340 1902.030 1688.400 ;
        RECT 1980.000 1688.340 1980.140 1688.880 ;
        RECT 1995.550 1688.820 1995.870 1688.880 ;
        RECT 1901.710 1688.200 1980.140 1688.340 ;
        RECT 1901.710 1688.140 1902.030 1688.200 ;
      LAYER via ;
        RECT 1901.740 1688.140 1902.000 1688.400 ;
        RECT 1995.580 1688.820 1995.840 1689.080 ;
      LAYER met2 ;
        RECT 1901.665 1700.000 1901.945 1704.000 ;
        RECT 1901.800 1688.430 1901.940 1700.000 ;
        RECT 1995.580 1688.790 1995.840 1689.110 ;
        RECT 1901.740 1688.110 1902.000 1688.430 ;
        RECT 1995.640 3.130 1995.780 1688.790 ;
        RECT 1995.180 2.990 1995.780 3.130 ;
        RECT 1995.180 2.400 1995.320 2.990 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1908.610 1687.320 1908.930 1687.380 ;
        RECT 1908.610 1687.180 1973.240 1687.320 ;
        RECT 1908.610 1687.120 1908.930 1687.180 ;
        RECT 1973.100 1686.640 1973.240 1687.180 ;
        RECT 2009.350 1686.640 2009.670 1686.700 ;
        RECT 1973.100 1686.500 2009.670 1686.640 ;
        RECT 2009.350 1686.440 2009.670 1686.500 ;
      LAYER via ;
        RECT 1908.640 1687.120 1908.900 1687.380 ;
        RECT 2009.380 1686.440 2009.640 1686.700 ;
      LAYER met2 ;
        RECT 1908.565 1700.000 1908.845 1704.000 ;
        RECT 1908.700 1687.410 1908.840 1700.000 ;
        RECT 1908.640 1687.090 1908.900 1687.410 ;
        RECT 2009.380 1686.410 2009.640 1686.730 ;
        RECT 2009.440 16.730 2009.580 1686.410 ;
        RECT 2009.440 16.590 2012.800 16.730 ;
        RECT 2012.660 2.400 2012.800 16.590 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1972.625 1686.825 1974.175 1686.995 ;
      LAYER mcon ;
        RECT 1974.005 1686.825 1974.175 1686.995 ;
      LAYER met1 ;
        RECT 1915.050 1686.980 1915.370 1687.040 ;
        RECT 1972.565 1686.980 1972.855 1687.025 ;
        RECT 1915.050 1686.840 1972.855 1686.980 ;
        RECT 1915.050 1686.780 1915.370 1686.840 ;
        RECT 1972.565 1686.795 1972.855 1686.840 ;
        RECT 1973.945 1686.980 1974.235 1687.025 ;
        RECT 2024.990 1686.980 2025.310 1687.040 ;
        RECT 1973.945 1686.840 2025.310 1686.980 ;
        RECT 1973.945 1686.795 1974.235 1686.840 ;
        RECT 2024.990 1686.780 2025.310 1686.840 ;
        RECT 2024.990 16.900 2025.310 16.960 ;
        RECT 2030.510 16.900 2030.830 16.960 ;
        RECT 2024.990 16.760 2030.830 16.900 ;
        RECT 2024.990 16.700 2025.310 16.760 ;
        RECT 2030.510 16.700 2030.830 16.760 ;
      LAYER via ;
        RECT 1915.080 1686.780 1915.340 1687.040 ;
        RECT 2025.020 1686.780 2025.280 1687.040 ;
        RECT 2025.020 16.700 2025.280 16.960 ;
        RECT 2030.540 16.700 2030.800 16.960 ;
      LAYER met2 ;
        RECT 1915.005 1700.000 1915.285 1704.000 ;
        RECT 1915.140 1687.070 1915.280 1700.000 ;
        RECT 1915.080 1686.750 1915.340 1687.070 ;
        RECT 2025.020 1686.750 2025.280 1687.070 ;
        RECT 2025.080 16.990 2025.220 1686.750 ;
        RECT 2025.020 16.670 2025.280 16.990 ;
        RECT 2030.540 16.670 2030.800 16.990 ;
        RECT 2030.600 2.400 2030.740 16.670 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1971.705 16.915 1971.875 18.955 ;
        RECT 1971.705 16.745 1972.335 16.915 ;
        RECT 2024.605 15.725 2024.775 16.915 ;
      LAYER mcon ;
        RECT 1971.705 18.785 1971.875 18.955 ;
        RECT 1972.165 16.745 1972.335 16.915 ;
        RECT 2024.605 16.745 2024.775 16.915 ;
      LAYER met1 ;
        RECT 1924.250 18.940 1924.570 19.000 ;
        RECT 1971.645 18.940 1971.935 18.985 ;
        RECT 1924.250 18.800 1971.935 18.940 ;
        RECT 1924.250 18.740 1924.570 18.800 ;
        RECT 1971.645 18.755 1971.935 18.800 ;
        RECT 1972.105 16.900 1972.395 16.945 ;
        RECT 2024.545 16.900 2024.835 16.945 ;
        RECT 1972.105 16.760 2024.835 16.900 ;
        RECT 1972.105 16.715 1972.395 16.760 ;
        RECT 2024.545 16.715 2024.835 16.760 ;
        RECT 2024.545 15.880 2024.835 15.925 ;
        RECT 2048.450 15.880 2048.770 15.940 ;
        RECT 2024.545 15.740 2048.770 15.880 ;
        RECT 2024.545 15.695 2024.835 15.740 ;
        RECT 2048.450 15.680 2048.770 15.740 ;
      LAYER via ;
        RECT 1924.280 18.740 1924.540 19.000 ;
        RECT 2048.480 15.680 2048.740 15.940 ;
      LAYER met2 ;
        RECT 1921.905 1701.090 1922.185 1704.000 ;
        RECT 1921.905 1700.950 1924.020 1701.090 ;
        RECT 1921.905 1700.000 1922.185 1700.950 ;
        RECT 1923.880 1688.850 1924.020 1700.950 ;
        RECT 1923.880 1688.710 1924.480 1688.850 ;
        RECT 1924.340 19.030 1924.480 1688.710 ;
        RECT 1924.280 18.710 1924.540 19.030 ;
        RECT 2048.480 15.650 2048.740 15.970 ;
        RECT 2048.540 2.400 2048.680 15.650 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 763.670 36.280 763.990 36.340 ;
        RECT 1435.270 36.280 1435.590 36.340 ;
        RECT 763.670 36.140 1435.590 36.280 ;
        RECT 763.670 36.080 763.990 36.140 ;
        RECT 1435.270 36.080 1435.590 36.140 ;
      LAYER via ;
        RECT 763.700 36.080 763.960 36.340 ;
        RECT 1435.300 36.080 1435.560 36.340 ;
      LAYER met2 ;
        RECT 1437.065 1700.410 1437.345 1704.000 ;
        RECT 1435.360 1700.270 1437.345 1700.410 ;
        RECT 1435.360 36.370 1435.500 1700.270 ;
        RECT 1437.065 1700.000 1437.345 1700.270 ;
        RECT 763.700 36.050 763.960 36.370 ;
        RECT 1435.300 36.050 1435.560 36.370 ;
        RECT 763.760 2.400 763.900 36.050 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1931.150 23.020 1931.470 23.080 ;
        RECT 2066.390 23.020 2066.710 23.080 ;
        RECT 1931.150 22.880 2066.710 23.020 ;
        RECT 1931.150 22.820 1931.470 22.880 ;
        RECT 2066.390 22.820 2066.710 22.880 ;
      LAYER via ;
        RECT 1931.180 22.820 1931.440 23.080 ;
        RECT 2066.420 22.820 2066.680 23.080 ;
      LAYER met2 ;
        RECT 1928.805 1700.410 1929.085 1704.000 ;
        RECT 1928.805 1700.270 1930.460 1700.410 ;
        RECT 1928.805 1700.000 1929.085 1700.270 ;
        RECT 1930.320 1688.850 1930.460 1700.270 ;
        RECT 1930.320 1688.710 1931.380 1688.850 ;
        RECT 1931.240 23.110 1931.380 1688.710 ;
        RECT 1931.180 22.790 1931.440 23.110 ;
        RECT 2066.420 22.790 2066.680 23.110 ;
        RECT 2066.480 2.400 2066.620 22.790 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1938.050 20.300 1938.370 20.360 ;
        RECT 1938.050 20.160 1970.020 20.300 ;
        RECT 1938.050 20.100 1938.370 20.160 ;
        RECT 1969.880 19.960 1970.020 20.160 ;
        RECT 2084.330 19.960 2084.650 20.020 ;
        RECT 1969.880 19.820 2084.650 19.960 ;
        RECT 2084.330 19.760 2084.650 19.820 ;
      LAYER via ;
        RECT 1938.080 20.100 1938.340 20.360 ;
        RECT 2084.360 19.760 2084.620 20.020 ;
      LAYER met2 ;
        RECT 1935.245 1700.410 1935.525 1704.000 ;
        RECT 1935.245 1700.270 1937.360 1700.410 ;
        RECT 1935.245 1700.000 1935.525 1700.270 ;
        RECT 1937.220 1688.850 1937.360 1700.270 ;
        RECT 1937.220 1688.710 1938.280 1688.850 ;
        RECT 1938.140 20.390 1938.280 1688.710 ;
        RECT 1938.080 20.070 1938.340 20.390 ;
        RECT 2084.360 19.730 2084.620 20.050 ;
        RECT 2084.420 2.400 2084.560 19.730 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1968.485 19.465 1970.035 19.635 ;
      LAYER mcon ;
        RECT 1969.865 19.465 1970.035 19.635 ;
      LAYER met1 ;
        RECT 1944.950 19.620 1945.270 19.680 ;
        RECT 1968.425 19.620 1968.715 19.665 ;
        RECT 1944.950 19.480 1968.715 19.620 ;
        RECT 1944.950 19.420 1945.270 19.480 ;
        RECT 1968.425 19.435 1968.715 19.480 ;
        RECT 1969.805 19.620 1970.095 19.665 ;
        RECT 2101.810 19.620 2102.130 19.680 ;
        RECT 1969.805 19.480 2102.130 19.620 ;
        RECT 1969.805 19.435 1970.095 19.480 ;
        RECT 2101.810 19.420 2102.130 19.480 ;
      LAYER via ;
        RECT 1944.980 19.420 1945.240 19.680 ;
        RECT 2101.840 19.420 2102.100 19.680 ;
      LAYER met2 ;
        RECT 1942.145 1701.090 1942.425 1704.000 ;
        RECT 1942.145 1700.950 1944.260 1701.090 ;
        RECT 1942.145 1700.000 1942.425 1700.950 ;
        RECT 1944.120 1688.850 1944.260 1700.950 ;
        RECT 1944.120 1688.710 1945.180 1688.850 ;
        RECT 1945.040 19.710 1945.180 1688.710 ;
        RECT 1944.980 19.390 1945.240 19.710 ;
        RECT 2101.840 19.390 2102.100 19.710 ;
        RECT 2101.900 2.400 2102.040 19.390 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1949.090 1685.280 1949.410 1685.340 ;
        RECT 1951.850 1685.280 1952.170 1685.340 ;
        RECT 1949.090 1685.140 1952.170 1685.280 ;
        RECT 1949.090 1685.080 1949.410 1685.140 ;
        RECT 1951.850 1685.080 1952.170 1685.140 ;
        RECT 1951.850 27.440 1952.170 27.500 ;
        RECT 2119.750 27.440 2120.070 27.500 ;
        RECT 1951.850 27.300 2120.070 27.440 ;
        RECT 1951.850 27.240 1952.170 27.300 ;
        RECT 2119.750 27.240 2120.070 27.300 ;
      LAYER via ;
        RECT 1949.120 1685.080 1949.380 1685.340 ;
        RECT 1951.880 1685.080 1952.140 1685.340 ;
        RECT 1951.880 27.240 1952.140 27.500 ;
        RECT 2119.780 27.240 2120.040 27.500 ;
      LAYER met2 ;
        RECT 1949.045 1700.000 1949.325 1704.000 ;
        RECT 1949.180 1685.370 1949.320 1700.000 ;
        RECT 1949.120 1685.050 1949.380 1685.370 ;
        RECT 1951.880 1685.050 1952.140 1685.370 ;
        RECT 1951.940 27.530 1952.080 1685.050 ;
        RECT 1951.880 27.210 1952.140 27.530 ;
        RECT 2119.780 27.210 2120.040 27.530 ;
        RECT 2119.840 2.400 2119.980 27.210 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1972.625 17.085 1972.795 18.955 ;
      LAYER mcon ;
        RECT 1972.625 18.785 1972.795 18.955 ;
      LAYER met1 ;
        RECT 1957.370 41.040 1957.690 41.100 ;
        RECT 1958.750 41.040 1959.070 41.100 ;
        RECT 1957.370 40.900 1959.070 41.040 ;
        RECT 1957.370 40.840 1957.690 40.900 ;
        RECT 1958.750 40.840 1959.070 40.900 ;
        RECT 1972.565 18.940 1972.855 18.985 ;
        RECT 2137.690 18.940 2138.010 19.000 ;
        RECT 1972.565 18.800 2138.010 18.940 ;
        RECT 1972.565 18.755 1972.855 18.800 ;
        RECT 2137.690 18.740 2138.010 18.800 ;
        RECT 1972.565 17.240 1972.855 17.285 ;
        RECT 1971.720 17.100 1972.855 17.240 ;
        RECT 1957.370 16.900 1957.690 16.960 ;
        RECT 1971.720 16.900 1971.860 17.100 ;
        RECT 1972.565 17.055 1972.855 17.100 ;
        RECT 1957.370 16.760 1971.860 16.900 ;
        RECT 1957.370 16.700 1957.690 16.760 ;
      LAYER via ;
        RECT 1957.400 40.840 1957.660 41.100 ;
        RECT 1958.780 40.840 1959.040 41.100 ;
        RECT 2137.720 18.740 2137.980 19.000 ;
        RECT 1957.400 16.700 1957.660 16.960 ;
      LAYER met2 ;
        RECT 1955.485 1700.410 1955.765 1704.000 ;
        RECT 1955.485 1700.270 1957.600 1700.410 ;
        RECT 1955.485 1700.000 1955.765 1700.270 ;
        RECT 1957.460 1688.850 1957.600 1700.270 ;
        RECT 1957.460 1688.710 1958.980 1688.850 ;
        RECT 1958.840 41.130 1958.980 1688.710 ;
        RECT 1957.400 40.810 1957.660 41.130 ;
        RECT 1958.780 40.810 1959.040 41.130 ;
        RECT 1957.460 16.990 1957.600 40.810 ;
        RECT 2137.720 18.710 2137.980 19.030 ;
        RECT 1957.400 16.670 1957.660 16.990 ;
        RECT 2137.780 2.400 2137.920 18.710 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1965.650 18.600 1965.970 18.660 ;
        RECT 1965.650 18.460 1970.940 18.600 ;
        RECT 1965.650 18.400 1965.970 18.460 ;
        RECT 1970.800 18.260 1970.940 18.460 ;
        RECT 2155.630 18.260 2155.950 18.320 ;
        RECT 1970.800 18.120 2155.950 18.260 ;
        RECT 2155.630 18.060 2155.950 18.120 ;
      LAYER via ;
        RECT 1965.680 18.400 1965.940 18.660 ;
        RECT 2155.660 18.060 2155.920 18.320 ;
      LAYER met2 ;
        RECT 1962.385 1700.410 1962.665 1704.000 ;
        RECT 1962.385 1700.270 1964.500 1700.410 ;
        RECT 1962.385 1700.000 1962.665 1700.270 ;
        RECT 1964.360 1688.850 1964.500 1700.270 ;
        RECT 1964.360 1688.710 1965.880 1688.850 ;
        RECT 1965.740 18.690 1965.880 1688.710 ;
        RECT 1965.680 18.370 1965.940 18.690 ;
        RECT 2155.660 18.030 2155.920 18.350 ;
        RECT 2155.720 2.400 2155.860 18.030 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1969.330 1689.020 1969.650 1689.080 ;
        RECT 1972.090 1689.020 1972.410 1689.080 ;
        RECT 1969.330 1688.880 1972.410 1689.020 ;
        RECT 1969.330 1688.820 1969.650 1688.880 ;
        RECT 1972.090 1688.820 1972.410 1688.880 ;
        RECT 1972.090 26.080 1972.410 26.140 ;
        RECT 2173.110 26.080 2173.430 26.140 ;
        RECT 1972.090 25.940 2173.430 26.080 ;
        RECT 1972.090 25.880 1972.410 25.940 ;
        RECT 2173.110 25.880 2173.430 25.940 ;
      LAYER via ;
        RECT 1969.360 1688.820 1969.620 1689.080 ;
        RECT 1972.120 1688.820 1972.380 1689.080 ;
        RECT 1972.120 25.880 1972.380 26.140 ;
        RECT 2173.140 25.880 2173.400 26.140 ;
      LAYER met2 ;
        RECT 1969.285 1700.000 1969.565 1704.000 ;
        RECT 1969.420 1689.110 1969.560 1700.000 ;
        RECT 1969.360 1688.790 1969.620 1689.110 ;
        RECT 1972.120 1688.790 1972.380 1689.110 ;
        RECT 1972.180 26.170 1972.320 1688.790 ;
        RECT 1972.120 25.850 1972.380 26.170 ;
        RECT 2173.140 25.850 2173.400 26.170 ;
        RECT 2173.200 2.400 2173.340 25.850 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1979.450 25.400 1979.770 25.460 ;
        RECT 2191.050 25.400 2191.370 25.460 ;
        RECT 1979.450 25.260 2191.370 25.400 ;
        RECT 1979.450 25.200 1979.770 25.260 ;
        RECT 2191.050 25.200 2191.370 25.260 ;
      LAYER via ;
        RECT 1979.480 25.200 1979.740 25.460 ;
        RECT 2191.080 25.200 2191.340 25.460 ;
      LAYER met2 ;
        RECT 1975.725 1700.410 1976.005 1704.000 ;
        RECT 1975.725 1700.270 1977.840 1700.410 ;
        RECT 1975.725 1700.000 1976.005 1700.270 ;
        RECT 1977.700 1688.680 1977.840 1700.270 ;
        RECT 1977.700 1688.540 1979.680 1688.680 ;
        RECT 1979.540 25.490 1979.680 1688.540 ;
        RECT 1979.480 25.170 1979.740 25.490 ;
        RECT 2191.080 25.170 2191.340 25.490 ;
        RECT 2191.140 2.400 2191.280 25.170 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1982.670 1688.680 1982.990 1688.740 ;
        RECT 1986.350 1688.680 1986.670 1688.740 ;
        RECT 1982.670 1688.540 1986.670 1688.680 ;
        RECT 1982.670 1688.480 1982.990 1688.540 ;
        RECT 1986.350 1688.480 1986.670 1688.540 ;
        RECT 1986.350 24.380 1986.670 24.440 ;
        RECT 2208.990 24.380 2209.310 24.440 ;
        RECT 1986.350 24.240 2209.310 24.380 ;
        RECT 1986.350 24.180 1986.670 24.240 ;
        RECT 2208.990 24.180 2209.310 24.240 ;
      LAYER via ;
        RECT 1982.700 1688.480 1982.960 1688.740 ;
        RECT 1986.380 1688.480 1986.640 1688.740 ;
        RECT 1986.380 24.180 1986.640 24.440 ;
        RECT 2209.020 24.180 2209.280 24.440 ;
      LAYER met2 ;
        RECT 1982.625 1700.000 1982.905 1704.000 ;
        RECT 1982.760 1688.770 1982.900 1700.000 ;
        RECT 1982.700 1688.450 1982.960 1688.770 ;
        RECT 1986.380 1688.450 1986.640 1688.770 ;
        RECT 1986.440 24.470 1986.580 1688.450 ;
        RECT 1986.380 24.150 1986.640 24.470 ;
        RECT 2209.020 24.150 2209.280 24.470 ;
        RECT 2209.080 2.400 2209.220 24.150 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1989.110 1688.680 1989.430 1688.740 ;
        RECT 1992.790 1688.680 1993.110 1688.740 ;
        RECT 1989.110 1688.540 1993.110 1688.680 ;
        RECT 1989.110 1688.480 1989.430 1688.540 ;
        RECT 1992.790 1688.480 1993.110 1688.540 ;
        RECT 1992.790 35.600 1993.110 35.660 ;
        RECT 2226.930 35.600 2227.250 35.660 ;
        RECT 1992.790 35.460 2227.250 35.600 ;
        RECT 1992.790 35.400 1993.110 35.460 ;
        RECT 2226.930 35.400 2227.250 35.460 ;
      LAYER via ;
        RECT 1989.140 1688.480 1989.400 1688.740 ;
        RECT 1992.820 1688.480 1993.080 1688.740 ;
        RECT 1992.820 35.400 1993.080 35.660 ;
        RECT 2226.960 35.400 2227.220 35.660 ;
      LAYER met2 ;
        RECT 1989.065 1700.000 1989.345 1704.000 ;
        RECT 1989.200 1688.770 1989.340 1700.000 ;
        RECT 1989.140 1688.450 1989.400 1688.770 ;
        RECT 1992.820 1688.450 1993.080 1688.770 ;
        RECT 1992.880 35.690 1993.020 1688.450 ;
        RECT 1992.820 35.370 1993.080 35.690 ;
        RECT 2226.960 35.370 2227.220 35.690 ;
        RECT 2227.020 2.400 2227.160 35.370 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 781.610 35.940 781.930 36.000 ;
        RECT 1442.170 35.940 1442.490 36.000 ;
        RECT 781.610 35.800 1442.490 35.940 ;
        RECT 781.610 35.740 781.930 35.800 ;
        RECT 1442.170 35.740 1442.490 35.800 ;
      LAYER via ;
        RECT 781.640 35.740 781.900 36.000 ;
        RECT 1442.200 35.740 1442.460 36.000 ;
      LAYER met2 ;
        RECT 1443.965 1700.410 1444.245 1704.000 ;
        RECT 1442.260 1700.270 1444.245 1700.410 ;
        RECT 1442.260 36.030 1442.400 1700.270 ;
        RECT 1443.965 1700.000 1444.245 1700.270 ;
        RECT 781.640 35.710 781.900 36.030 ;
        RECT 1442.200 35.710 1442.460 36.030 ;
        RECT 781.700 2.400 781.840 35.710 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1996.010 1688.680 1996.330 1688.740 ;
        RECT 2000.150 1688.680 2000.470 1688.740 ;
        RECT 1996.010 1688.540 2000.470 1688.680 ;
        RECT 1996.010 1688.480 1996.330 1688.540 ;
        RECT 2000.150 1688.480 2000.470 1688.540 ;
        RECT 2000.150 44.780 2000.470 44.840 ;
        RECT 2244.870 44.780 2245.190 44.840 ;
        RECT 2000.150 44.640 2245.190 44.780 ;
        RECT 2000.150 44.580 2000.470 44.640 ;
        RECT 2244.870 44.580 2245.190 44.640 ;
      LAYER via ;
        RECT 1996.040 1688.480 1996.300 1688.740 ;
        RECT 2000.180 1688.480 2000.440 1688.740 ;
        RECT 2000.180 44.580 2000.440 44.840 ;
        RECT 2244.900 44.580 2245.160 44.840 ;
      LAYER met2 ;
        RECT 1995.965 1700.000 1996.245 1704.000 ;
        RECT 1996.100 1688.770 1996.240 1700.000 ;
        RECT 1996.040 1688.450 1996.300 1688.770 ;
        RECT 2000.180 1688.450 2000.440 1688.770 ;
        RECT 2000.240 44.870 2000.380 1688.450 ;
        RECT 2000.180 44.550 2000.440 44.870 ;
        RECT 2244.900 44.550 2245.160 44.870 ;
        RECT 2244.960 2.400 2245.100 44.550 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2002.910 1688.680 2003.230 1688.740 ;
        RECT 2007.050 1688.680 2007.370 1688.740 ;
        RECT 2002.910 1688.540 2007.370 1688.680 ;
        RECT 2002.910 1688.480 2003.230 1688.540 ;
        RECT 2007.050 1688.480 2007.370 1688.540 ;
        RECT 2007.050 43.760 2007.370 43.820 ;
        RECT 2262.350 43.760 2262.670 43.820 ;
        RECT 2007.050 43.620 2262.670 43.760 ;
        RECT 2007.050 43.560 2007.370 43.620 ;
        RECT 2262.350 43.560 2262.670 43.620 ;
      LAYER via ;
        RECT 2002.940 1688.480 2003.200 1688.740 ;
        RECT 2007.080 1688.480 2007.340 1688.740 ;
        RECT 2007.080 43.560 2007.340 43.820 ;
        RECT 2262.380 43.560 2262.640 43.820 ;
      LAYER met2 ;
        RECT 2002.865 1700.000 2003.145 1704.000 ;
        RECT 2003.000 1688.770 2003.140 1700.000 ;
        RECT 2002.940 1688.450 2003.200 1688.770 ;
        RECT 2007.080 1688.450 2007.340 1688.770 ;
        RECT 2007.140 43.850 2007.280 1688.450 ;
        RECT 2007.080 43.530 2007.340 43.850 ;
        RECT 2262.380 43.530 2262.640 43.850 ;
        RECT 2262.440 2.400 2262.580 43.530 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2009.350 1688.680 2009.670 1688.740 ;
        RECT 2013.950 1688.680 2014.270 1688.740 ;
        RECT 2009.350 1688.540 2014.270 1688.680 ;
        RECT 2009.350 1688.480 2009.670 1688.540 ;
        RECT 2013.950 1688.480 2014.270 1688.540 ;
        RECT 2013.950 44.100 2014.270 44.160 ;
        RECT 2280.290 44.100 2280.610 44.160 ;
        RECT 2013.950 43.960 2280.610 44.100 ;
        RECT 2013.950 43.900 2014.270 43.960 ;
        RECT 2280.290 43.900 2280.610 43.960 ;
      LAYER via ;
        RECT 2009.380 1688.480 2009.640 1688.740 ;
        RECT 2013.980 1688.480 2014.240 1688.740 ;
        RECT 2013.980 43.900 2014.240 44.160 ;
        RECT 2280.320 43.900 2280.580 44.160 ;
      LAYER met2 ;
        RECT 2009.305 1700.000 2009.585 1704.000 ;
        RECT 2009.440 1688.770 2009.580 1700.000 ;
        RECT 2009.380 1688.450 2009.640 1688.770 ;
        RECT 2013.980 1688.450 2014.240 1688.770 ;
        RECT 2014.040 44.190 2014.180 1688.450 ;
        RECT 2013.980 43.870 2014.240 44.190 ;
        RECT 2280.320 43.870 2280.580 44.190 ;
        RECT 2280.380 2.400 2280.520 43.870 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2016.250 1688.680 2016.570 1688.740 ;
        RECT 2020.850 1688.680 2021.170 1688.740 ;
        RECT 2016.250 1688.540 2021.170 1688.680 ;
        RECT 2016.250 1688.480 2016.570 1688.540 ;
        RECT 2020.850 1688.480 2021.170 1688.540 ;
        RECT 2020.850 44.440 2021.170 44.500 ;
        RECT 2298.230 44.440 2298.550 44.500 ;
        RECT 2020.850 44.300 2298.550 44.440 ;
        RECT 2020.850 44.240 2021.170 44.300 ;
        RECT 2298.230 44.240 2298.550 44.300 ;
      LAYER via ;
        RECT 2016.280 1688.480 2016.540 1688.740 ;
        RECT 2020.880 1688.480 2021.140 1688.740 ;
        RECT 2020.880 44.240 2021.140 44.500 ;
        RECT 2298.260 44.240 2298.520 44.500 ;
      LAYER met2 ;
        RECT 2016.205 1700.000 2016.485 1704.000 ;
        RECT 2016.340 1688.770 2016.480 1700.000 ;
        RECT 2016.280 1688.450 2016.540 1688.770 ;
        RECT 2020.880 1688.450 2021.140 1688.770 ;
        RECT 2020.940 44.530 2021.080 1688.450 ;
        RECT 2020.880 44.210 2021.140 44.530 ;
        RECT 2298.260 44.210 2298.520 44.530 ;
        RECT 2298.320 2.400 2298.460 44.210 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2023.150 1688.680 2023.470 1688.740 ;
        RECT 2027.750 1688.680 2028.070 1688.740 ;
        RECT 2023.150 1688.540 2028.070 1688.680 ;
        RECT 2023.150 1688.480 2023.470 1688.540 ;
        RECT 2027.750 1688.480 2028.070 1688.540 ;
        RECT 2027.750 48.180 2028.070 48.240 ;
        RECT 2316.170 48.180 2316.490 48.240 ;
        RECT 2027.750 48.040 2316.490 48.180 ;
        RECT 2027.750 47.980 2028.070 48.040 ;
        RECT 2316.170 47.980 2316.490 48.040 ;
      LAYER via ;
        RECT 2023.180 1688.480 2023.440 1688.740 ;
        RECT 2027.780 1688.480 2028.040 1688.740 ;
        RECT 2027.780 47.980 2028.040 48.240 ;
        RECT 2316.200 47.980 2316.460 48.240 ;
      LAYER met2 ;
        RECT 2023.105 1700.000 2023.385 1704.000 ;
        RECT 2023.240 1688.770 2023.380 1700.000 ;
        RECT 2023.180 1688.450 2023.440 1688.770 ;
        RECT 2027.780 1688.450 2028.040 1688.770 ;
        RECT 2027.840 48.270 2027.980 1688.450 ;
        RECT 2027.780 47.950 2028.040 48.270 ;
        RECT 2316.200 47.950 2316.460 48.270 ;
        RECT 2316.260 2.400 2316.400 47.950 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2029.590 1688.680 2029.910 1688.740 ;
        RECT 2034.650 1688.680 2034.970 1688.740 ;
        RECT 2029.590 1688.540 2034.970 1688.680 ;
        RECT 2029.590 1688.480 2029.910 1688.540 ;
        RECT 2034.650 1688.480 2034.970 1688.540 ;
        RECT 2034.650 47.840 2034.970 47.900 ;
        RECT 2334.110 47.840 2334.430 47.900 ;
        RECT 2034.650 47.700 2334.430 47.840 ;
        RECT 2034.650 47.640 2034.970 47.700 ;
        RECT 2334.110 47.640 2334.430 47.700 ;
      LAYER via ;
        RECT 2029.620 1688.480 2029.880 1688.740 ;
        RECT 2034.680 1688.480 2034.940 1688.740 ;
        RECT 2034.680 47.640 2034.940 47.900 ;
        RECT 2334.140 47.640 2334.400 47.900 ;
      LAYER met2 ;
        RECT 2029.545 1700.000 2029.825 1704.000 ;
        RECT 2029.680 1688.770 2029.820 1700.000 ;
        RECT 2029.620 1688.450 2029.880 1688.770 ;
        RECT 2034.680 1688.450 2034.940 1688.770 ;
        RECT 2034.740 47.930 2034.880 1688.450 ;
        RECT 2034.680 47.610 2034.940 47.930 ;
        RECT 2334.140 47.610 2334.400 47.930 ;
        RECT 2334.200 2.400 2334.340 47.610 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2036.490 1688.680 2036.810 1688.740 ;
        RECT 2041.550 1688.680 2041.870 1688.740 ;
        RECT 2036.490 1688.540 2041.870 1688.680 ;
        RECT 2036.490 1688.480 2036.810 1688.540 ;
        RECT 2041.550 1688.480 2041.870 1688.540 ;
        RECT 2041.550 47.500 2041.870 47.560 ;
        RECT 2351.590 47.500 2351.910 47.560 ;
        RECT 2041.550 47.360 2351.910 47.500 ;
        RECT 2041.550 47.300 2041.870 47.360 ;
        RECT 2351.590 47.300 2351.910 47.360 ;
      LAYER via ;
        RECT 2036.520 1688.480 2036.780 1688.740 ;
        RECT 2041.580 1688.480 2041.840 1688.740 ;
        RECT 2041.580 47.300 2041.840 47.560 ;
        RECT 2351.620 47.300 2351.880 47.560 ;
      LAYER met2 ;
        RECT 2036.445 1700.000 2036.725 1704.000 ;
        RECT 2036.580 1688.770 2036.720 1700.000 ;
        RECT 2036.520 1688.450 2036.780 1688.770 ;
        RECT 2041.580 1688.450 2041.840 1688.770 ;
        RECT 2041.640 47.590 2041.780 1688.450 ;
        RECT 2041.580 47.270 2041.840 47.590 ;
        RECT 2351.620 47.270 2351.880 47.590 ;
        RECT 2351.680 2.400 2351.820 47.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2176.405 1682.405 2176.575 1688.015 ;
        RECT 2231.605 13.685 2231.775 14.535 ;
      LAYER mcon ;
        RECT 2176.405 1687.845 2176.575 1688.015 ;
        RECT 2231.605 14.365 2231.775 14.535 ;
      LAYER met1 ;
        RECT 2043.390 1688.000 2043.710 1688.060 ;
        RECT 2176.345 1688.000 2176.635 1688.045 ;
        RECT 2043.390 1687.860 2176.635 1688.000 ;
        RECT 2043.390 1687.800 2043.710 1687.860 ;
        RECT 2176.345 1687.815 2176.635 1687.860 ;
        RECT 2176.345 1682.560 2176.635 1682.605 ;
        RECT 2211.290 1682.560 2211.610 1682.620 ;
        RECT 2176.345 1682.420 2211.610 1682.560 ;
        RECT 2176.345 1682.375 2176.635 1682.420 ;
        RECT 2211.290 1682.360 2211.610 1682.420 ;
        RECT 2211.290 14.520 2211.610 14.580 ;
        RECT 2231.545 14.520 2231.835 14.565 ;
        RECT 2211.290 14.380 2231.835 14.520 ;
        RECT 2211.290 14.320 2211.610 14.380 ;
        RECT 2231.545 14.335 2231.835 14.380 ;
        RECT 2369.530 14.180 2369.850 14.240 ;
        RECT 2240.360 14.040 2369.850 14.180 ;
        RECT 2231.545 13.840 2231.835 13.885 ;
        RECT 2240.360 13.840 2240.500 14.040 ;
        RECT 2369.530 13.980 2369.850 14.040 ;
        RECT 2231.545 13.700 2240.500 13.840 ;
        RECT 2231.545 13.655 2231.835 13.700 ;
      LAYER via ;
        RECT 2043.420 1687.800 2043.680 1688.060 ;
        RECT 2211.320 1682.360 2211.580 1682.620 ;
        RECT 2211.320 14.320 2211.580 14.580 ;
        RECT 2369.560 13.980 2369.820 14.240 ;
      LAYER met2 ;
        RECT 2043.345 1700.000 2043.625 1704.000 ;
        RECT 2043.480 1688.090 2043.620 1700.000 ;
        RECT 2043.420 1687.770 2043.680 1688.090 ;
        RECT 2211.320 1682.330 2211.580 1682.650 ;
        RECT 2211.380 14.610 2211.520 1682.330 ;
        RECT 2211.320 14.290 2211.580 14.610 ;
        RECT 2369.560 13.950 2369.820 14.270 ;
        RECT 2369.620 2.400 2369.760 13.950 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2049.830 1685.280 2050.150 1685.340 ;
        RECT 2387.930 1685.280 2388.250 1685.340 ;
        RECT 2049.830 1685.140 2388.250 1685.280 ;
        RECT 2049.830 1685.080 2050.150 1685.140 ;
        RECT 2387.930 1685.080 2388.250 1685.140 ;
      LAYER via ;
        RECT 2049.860 1685.080 2050.120 1685.340 ;
        RECT 2387.960 1685.080 2388.220 1685.340 ;
      LAYER met2 ;
        RECT 2049.785 1700.000 2050.065 1704.000 ;
        RECT 2049.920 1685.370 2050.060 1700.000 ;
        RECT 2049.860 1685.050 2050.120 1685.370 ;
        RECT 2387.960 1685.050 2388.220 1685.370 ;
        RECT 2388.020 17.410 2388.160 1685.050 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2141.445 1686.825 2141.615 1687.675 ;
      LAYER mcon ;
        RECT 2141.445 1687.505 2141.615 1687.675 ;
      LAYER met1 ;
        RECT 2141.385 1687.660 2141.675 1687.705 ;
        RECT 2169.890 1687.660 2170.210 1687.720 ;
        RECT 2141.385 1687.520 2170.210 1687.660 ;
        RECT 2141.385 1687.475 2141.675 1687.520 ;
        RECT 2169.890 1687.460 2170.210 1687.520 ;
        RECT 2056.730 1686.980 2057.050 1687.040 ;
        RECT 2141.385 1686.980 2141.675 1687.025 ;
        RECT 2056.730 1686.840 2141.675 1686.980 ;
        RECT 2056.730 1686.780 2057.050 1686.840 ;
        RECT 2141.385 1686.795 2141.675 1686.840 ;
        RECT 2169.890 15.200 2170.210 15.260 ;
        RECT 2405.410 15.200 2405.730 15.260 ;
        RECT 2169.890 15.060 2405.730 15.200 ;
        RECT 2169.890 15.000 2170.210 15.060 ;
        RECT 2405.410 15.000 2405.730 15.060 ;
      LAYER via ;
        RECT 2169.920 1687.460 2170.180 1687.720 ;
        RECT 2056.760 1686.780 2057.020 1687.040 ;
        RECT 2169.920 15.000 2170.180 15.260 ;
        RECT 2405.440 15.000 2405.700 15.260 ;
      LAYER met2 ;
        RECT 2056.685 1700.000 2056.965 1704.000 ;
        RECT 2056.820 1687.070 2056.960 1700.000 ;
        RECT 2169.920 1687.430 2170.180 1687.750 ;
        RECT 2056.760 1686.750 2057.020 1687.070 ;
        RECT 2169.980 15.290 2170.120 1687.430 ;
        RECT 2169.920 14.970 2170.180 15.290 ;
        RECT 2405.440 14.970 2405.700 15.290 ;
        RECT 2405.500 2.400 2405.640 14.970 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1449.070 35.600 1449.390 35.660 ;
        RECT 800.560 35.460 1449.390 35.600 ;
        RECT 799.550 35.260 799.870 35.320 ;
        RECT 800.560 35.260 800.700 35.460 ;
        RECT 1449.070 35.400 1449.390 35.460 ;
        RECT 799.550 35.120 800.700 35.260 ;
        RECT 799.550 35.060 799.870 35.120 ;
      LAYER via ;
        RECT 799.580 35.060 799.840 35.320 ;
        RECT 1449.100 35.400 1449.360 35.660 ;
      LAYER met2 ;
        RECT 1450.405 1700.410 1450.685 1704.000 ;
        RECT 1449.160 1700.270 1450.685 1700.410 ;
        RECT 1449.160 35.690 1449.300 1700.270 ;
        RECT 1450.405 1700.000 1450.685 1700.270 ;
        RECT 1449.100 35.370 1449.360 35.690 ;
        RECT 799.580 35.030 799.840 35.350 ;
        RECT 799.640 2.400 799.780 35.030 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1255.945 39.865 1256.115 41.395 ;
        RECT 1272.965 39.865 1273.135 41.395 ;
      LAYER mcon ;
        RECT 1255.945 41.225 1256.115 41.395 ;
        RECT 1272.965 41.225 1273.135 41.395 ;
      LAYER met1 ;
        RECT 1386.970 1678.480 1387.290 1678.540 ;
        RECT 1390.650 1678.480 1390.970 1678.540 ;
        RECT 1386.970 1678.340 1390.970 1678.480 ;
        RECT 1386.970 1678.280 1387.290 1678.340 ;
        RECT 1390.650 1678.280 1390.970 1678.340 ;
        RECT 644.990 41.380 645.310 41.440 ;
        RECT 1255.885 41.380 1256.175 41.425 ;
        RECT 644.990 41.240 1256.175 41.380 ;
        RECT 644.990 41.180 645.310 41.240 ;
        RECT 1255.885 41.195 1256.175 41.240 ;
        RECT 1272.905 41.380 1273.195 41.425 ;
        RECT 1386.970 41.380 1387.290 41.440 ;
        RECT 1272.905 41.240 1387.290 41.380 ;
        RECT 1272.905 41.195 1273.195 41.240 ;
        RECT 1386.970 41.180 1387.290 41.240 ;
        RECT 1255.885 40.020 1256.175 40.065 ;
        RECT 1272.905 40.020 1273.195 40.065 ;
        RECT 1255.885 39.880 1273.195 40.020 ;
        RECT 1255.885 39.835 1256.175 39.880 ;
        RECT 1272.905 39.835 1273.195 39.880 ;
      LAYER via ;
        RECT 1387.000 1678.280 1387.260 1678.540 ;
        RECT 1390.680 1678.280 1390.940 1678.540 ;
        RECT 645.020 41.180 645.280 41.440 ;
        RECT 1387.000 41.180 1387.260 41.440 ;
      LAYER met2 ;
        RECT 1391.985 1700.410 1392.265 1704.000 ;
        RECT 1390.740 1700.270 1392.265 1700.410 ;
        RECT 1390.740 1678.570 1390.880 1700.270 ;
        RECT 1391.985 1700.000 1392.265 1700.270 ;
        RECT 1387.000 1678.250 1387.260 1678.570 ;
        RECT 1390.680 1678.250 1390.940 1678.570 ;
        RECT 1387.060 41.470 1387.200 1678.250 ;
        RECT 645.020 41.150 645.280 41.470 ;
        RECT 1387.000 41.150 1387.260 41.470 ;
        RECT 645.080 2.400 645.220 41.150 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2065.470 1685.960 2065.790 1686.020 ;
        RECT 2428.870 1685.960 2429.190 1686.020 ;
        RECT 2065.470 1685.820 2429.190 1685.960 ;
        RECT 2065.470 1685.760 2065.790 1685.820 ;
        RECT 2428.870 1685.760 2429.190 1685.820 ;
      LAYER via ;
        RECT 2065.500 1685.760 2065.760 1686.020 ;
        RECT 2428.900 1685.760 2429.160 1686.020 ;
      LAYER met2 ;
        RECT 2065.425 1700.000 2065.705 1704.000 ;
        RECT 2065.560 1686.050 2065.700 1700.000 ;
        RECT 2065.500 1685.730 2065.760 1686.050 ;
        RECT 2428.900 1685.730 2429.160 1686.050 ;
        RECT 2428.960 2.400 2429.100 1685.730 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2085.325 1687.165 2085.495 1688.355 ;
        RECT 2140.525 1683.425 2140.695 1687.335 ;
        RECT 2211.365 16.065 2211.535 17.935 ;
      LAYER mcon ;
        RECT 2085.325 1688.185 2085.495 1688.355 ;
        RECT 2140.525 1687.165 2140.695 1687.335 ;
        RECT 2211.365 17.765 2211.535 17.935 ;
      LAYER met1 ;
        RECT 2072.370 1688.340 2072.690 1688.400 ;
        RECT 2085.265 1688.340 2085.555 1688.385 ;
        RECT 2072.370 1688.200 2085.555 1688.340 ;
        RECT 2072.370 1688.140 2072.690 1688.200 ;
        RECT 2085.265 1688.155 2085.555 1688.200 ;
        RECT 2085.265 1687.320 2085.555 1687.365 ;
        RECT 2140.465 1687.320 2140.755 1687.365 ;
        RECT 2085.265 1687.180 2140.755 1687.320 ;
        RECT 2085.265 1687.135 2085.555 1687.180 ;
        RECT 2140.465 1687.135 2140.755 1687.180 ;
        RECT 2140.465 1683.580 2140.755 1683.625 ;
        RECT 2176.790 1683.580 2177.110 1683.640 ;
        RECT 2140.465 1683.440 2177.110 1683.580 ;
        RECT 2140.465 1683.395 2140.755 1683.440 ;
        RECT 2176.790 1683.380 2177.110 1683.440 ;
        RECT 2177.250 738.520 2177.570 738.780 ;
        RECT 2177.340 738.100 2177.480 738.520 ;
        RECT 2177.250 737.840 2177.570 738.100 ;
        RECT 2177.250 17.920 2177.570 17.980 ;
        RECT 2211.305 17.920 2211.595 17.965 ;
        RECT 2177.250 17.780 2211.595 17.920 ;
        RECT 2177.250 17.720 2177.570 17.780 ;
        RECT 2211.305 17.735 2211.595 17.780 ;
        RECT 2211.305 16.220 2211.595 16.265 ;
        RECT 2446.810 16.220 2447.130 16.280 ;
        RECT 2211.305 16.080 2447.130 16.220 ;
        RECT 2211.305 16.035 2211.595 16.080 ;
        RECT 2446.810 16.020 2447.130 16.080 ;
      LAYER via ;
        RECT 2072.400 1688.140 2072.660 1688.400 ;
        RECT 2176.820 1683.380 2177.080 1683.640 ;
        RECT 2177.280 738.520 2177.540 738.780 ;
        RECT 2177.280 737.840 2177.540 738.100 ;
        RECT 2177.280 17.720 2177.540 17.980 ;
        RECT 2446.840 16.020 2447.100 16.280 ;
      LAYER met2 ;
        RECT 2072.325 1700.000 2072.605 1704.000 ;
        RECT 2072.460 1688.430 2072.600 1700.000 ;
        RECT 2072.400 1688.110 2072.660 1688.430 ;
        RECT 2176.820 1683.350 2177.080 1683.670 ;
        RECT 2176.880 1677.290 2177.020 1683.350 ;
        RECT 2176.880 1677.150 2177.480 1677.290 ;
        RECT 2177.340 738.810 2177.480 1677.150 ;
        RECT 2177.280 738.490 2177.540 738.810 ;
        RECT 2177.280 737.810 2177.540 738.130 ;
        RECT 2177.340 18.010 2177.480 737.810 ;
        RECT 2177.280 17.690 2177.540 18.010 ;
        RECT 2446.840 15.990 2447.100 16.310 ;
        RECT 2446.900 2.400 2447.040 15.990 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2135.465 1686.145 2135.635 1689.715 ;
      LAYER mcon ;
        RECT 2135.465 1689.545 2135.635 1689.715 ;
      LAYER met1 ;
        RECT 2079.270 1689.700 2079.590 1689.760 ;
        RECT 2135.405 1689.700 2135.695 1689.745 ;
        RECT 2079.270 1689.560 2135.695 1689.700 ;
        RECT 2079.270 1689.500 2079.590 1689.560 ;
        RECT 2135.405 1689.515 2135.695 1689.560 ;
        RECT 2135.405 1686.300 2135.695 1686.345 ;
        RECT 2463.370 1686.300 2463.690 1686.360 ;
        RECT 2135.405 1686.160 2463.690 1686.300 ;
        RECT 2135.405 1686.115 2135.695 1686.160 ;
        RECT 2463.370 1686.100 2463.690 1686.160 ;
        RECT 2463.370 2.960 2463.690 3.020 ;
        RECT 2464.750 2.960 2465.070 3.020 ;
        RECT 2463.370 2.820 2465.070 2.960 ;
        RECT 2463.370 2.760 2463.690 2.820 ;
        RECT 2464.750 2.760 2465.070 2.820 ;
      LAYER via ;
        RECT 2079.300 1689.500 2079.560 1689.760 ;
        RECT 2463.400 1686.100 2463.660 1686.360 ;
        RECT 2463.400 2.760 2463.660 3.020 ;
        RECT 2464.780 2.760 2465.040 3.020 ;
      LAYER met2 ;
        RECT 2079.225 1700.000 2079.505 1704.000 ;
        RECT 2079.360 1689.790 2079.500 1700.000 ;
        RECT 2079.300 1689.470 2079.560 1689.790 ;
        RECT 2463.400 1686.070 2463.660 1686.390 ;
        RECT 2463.460 3.050 2463.600 1686.070 ;
        RECT 2463.400 2.730 2463.660 3.050 ;
        RECT 2464.780 2.730 2465.040 3.050 ;
        RECT 2464.840 2.400 2464.980 2.730 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2128.105 1688.525 2128.275 1690.735 ;
      LAYER mcon ;
        RECT 2128.105 1690.565 2128.275 1690.735 ;
      LAYER met1 ;
        RECT 2128.045 1690.720 2128.335 1690.765 ;
        RECT 2128.045 1690.580 2135.620 1690.720 ;
        RECT 2128.045 1690.535 2128.335 1690.580 ;
        RECT 2135.480 1690.380 2135.620 1690.580 ;
        RECT 2156.090 1690.380 2156.410 1690.440 ;
        RECT 2135.480 1690.240 2156.410 1690.380 ;
        RECT 2156.090 1690.180 2156.410 1690.240 ;
        RECT 2128.045 1688.680 2128.335 1688.725 ;
        RECT 2125.820 1688.540 2128.335 1688.680 ;
        RECT 2085.710 1688.340 2086.030 1688.400 ;
        RECT 2125.820 1688.340 2125.960 1688.540 ;
        RECT 2128.045 1688.495 2128.335 1688.540 ;
        RECT 2085.710 1688.200 2125.960 1688.340 ;
        RECT 2085.710 1688.140 2086.030 1688.200 ;
        RECT 2156.090 16.900 2156.410 16.960 ;
        RECT 2482.690 16.900 2483.010 16.960 ;
        RECT 2156.090 16.760 2483.010 16.900 ;
        RECT 2156.090 16.700 2156.410 16.760 ;
        RECT 2482.690 16.700 2483.010 16.760 ;
      LAYER via ;
        RECT 2156.120 1690.180 2156.380 1690.440 ;
        RECT 2085.740 1688.140 2086.000 1688.400 ;
        RECT 2156.120 16.700 2156.380 16.960 ;
        RECT 2482.720 16.700 2482.980 16.960 ;
      LAYER met2 ;
        RECT 2085.665 1700.000 2085.945 1704.000 ;
        RECT 2085.800 1688.430 2085.940 1700.000 ;
        RECT 2156.120 1690.150 2156.380 1690.470 ;
        RECT 2085.740 1688.110 2086.000 1688.430 ;
        RECT 2156.180 16.990 2156.320 1690.150 ;
        RECT 2156.120 16.670 2156.380 16.990 ;
        RECT 2482.720 16.670 2482.980 16.990 ;
        RECT 2482.780 2.400 2482.920 16.670 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2135.005 1686.485 2135.175 1690.395 ;
      LAYER mcon ;
        RECT 2135.005 1690.225 2135.175 1690.395 ;
      LAYER met1 ;
        RECT 2092.610 1690.380 2092.930 1690.440 ;
        RECT 2134.945 1690.380 2135.235 1690.425 ;
        RECT 2092.610 1690.240 2135.235 1690.380 ;
        RECT 2092.610 1690.180 2092.930 1690.240 ;
        RECT 2134.945 1690.195 2135.235 1690.240 ;
        RECT 2134.945 1686.640 2135.235 1686.685 ;
        RECT 2480.390 1686.640 2480.710 1686.700 ;
        RECT 2134.945 1686.500 2480.710 1686.640 ;
        RECT 2134.945 1686.455 2135.235 1686.500 ;
        RECT 2480.390 1686.440 2480.710 1686.500 ;
        RECT 2480.390 15.880 2480.710 15.940 ;
        RECT 2500.630 15.880 2500.950 15.940 ;
        RECT 2480.390 15.740 2500.950 15.880 ;
        RECT 2480.390 15.680 2480.710 15.740 ;
        RECT 2500.630 15.680 2500.950 15.740 ;
      LAYER via ;
        RECT 2092.640 1690.180 2092.900 1690.440 ;
        RECT 2480.420 1686.440 2480.680 1686.700 ;
        RECT 2480.420 15.680 2480.680 15.940 ;
        RECT 2500.660 15.680 2500.920 15.940 ;
      LAYER met2 ;
        RECT 2092.565 1700.000 2092.845 1704.000 ;
        RECT 2092.700 1690.470 2092.840 1700.000 ;
        RECT 2092.640 1690.150 2092.900 1690.470 ;
        RECT 2480.420 1686.410 2480.680 1686.730 ;
        RECT 2480.480 15.970 2480.620 1686.410 ;
        RECT 2480.420 15.650 2480.680 15.970 ;
        RECT 2500.660 15.650 2500.920 15.970 ;
        RECT 2500.720 2.400 2500.860 15.650 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2099.510 1686.300 2099.830 1686.360 ;
        RECT 2107.790 1686.300 2108.110 1686.360 ;
        RECT 2099.510 1686.160 2108.110 1686.300 ;
        RECT 2099.510 1686.100 2099.830 1686.160 ;
        RECT 2107.790 1686.100 2108.110 1686.160 ;
        RECT 2107.790 20.640 2108.110 20.700 ;
        RECT 2518.110 20.640 2518.430 20.700 ;
        RECT 2107.790 20.500 2518.430 20.640 ;
        RECT 2107.790 20.440 2108.110 20.500 ;
        RECT 2518.110 20.440 2518.430 20.500 ;
      LAYER via ;
        RECT 2099.540 1686.100 2099.800 1686.360 ;
        RECT 2107.820 1686.100 2108.080 1686.360 ;
        RECT 2107.820 20.440 2108.080 20.700 ;
        RECT 2518.140 20.440 2518.400 20.700 ;
      LAYER met2 ;
        RECT 2099.465 1700.000 2099.745 1704.000 ;
        RECT 2099.600 1686.390 2099.740 1700.000 ;
        RECT 2099.540 1686.070 2099.800 1686.390 ;
        RECT 2107.820 1686.070 2108.080 1686.390 ;
        RECT 2107.880 20.730 2108.020 1686.070 ;
        RECT 2107.820 20.410 2108.080 20.730 ;
        RECT 2518.140 20.410 2518.400 20.730 ;
        RECT 2518.200 2.400 2518.340 20.410 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2105.950 1690.040 2106.270 1690.100 ;
        RECT 2501.090 1690.040 2501.410 1690.100 ;
        RECT 2105.950 1689.900 2501.410 1690.040 ;
        RECT 2105.950 1689.840 2106.270 1689.900 ;
        RECT 2501.090 1689.840 2501.410 1689.900 ;
        RECT 2501.090 16.900 2501.410 16.960 ;
        RECT 2536.050 16.900 2536.370 16.960 ;
        RECT 2501.090 16.760 2536.370 16.900 ;
        RECT 2501.090 16.700 2501.410 16.760 ;
        RECT 2536.050 16.700 2536.370 16.760 ;
      LAYER via ;
        RECT 2105.980 1689.840 2106.240 1690.100 ;
        RECT 2501.120 1689.840 2501.380 1690.100 ;
        RECT 2501.120 16.700 2501.380 16.960 ;
        RECT 2536.080 16.700 2536.340 16.960 ;
      LAYER met2 ;
        RECT 2105.905 1700.000 2106.185 1704.000 ;
        RECT 2106.040 1690.130 2106.180 1700.000 ;
        RECT 2105.980 1689.810 2106.240 1690.130 ;
        RECT 2501.120 1689.810 2501.380 1690.130 ;
        RECT 2501.180 16.990 2501.320 1689.810 ;
        RECT 2501.120 16.670 2501.380 16.990 ;
        RECT 2536.080 16.670 2536.340 16.990 ;
        RECT 2536.140 2.400 2536.280 16.670 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2135.850 1689.700 2136.170 1689.760 ;
        RECT 2142.290 1689.700 2142.610 1689.760 ;
        RECT 2135.850 1689.560 2142.610 1689.700 ;
        RECT 2135.850 1689.500 2136.170 1689.560 ;
        RECT 2142.290 1689.500 2142.610 1689.560 ;
        RECT 2112.850 1689.020 2113.170 1689.080 ;
        RECT 2112.850 1688.880 2132.860 1689.020 ;
        RECT 2112.850 1688.820 2113.170 1688.880 ;
        RECT 2132.720 1688.680 2132.860 1688.880 ;
        RECT 2134.930 1688.680 2135.250 1688.740 ;
        RECT 2132.720 1688.540 2135.250 1688.680 ;
        RECT 2134.930 1688.480 2135.250 1688.540 ;
        RECT 2142.290 20.300 2142.610 20.360 ;
        RECT 2553.990 20.300 2554.310 20.360 ;
        RECT 2142.290 20.160 2554.310 20.300 ;
        RECT 2142.290 20.100 2142.610 20.160 ;
        RECT 2553.990 20.100 2554.310 20.160 ;
      LAYER via ;
        RECT 2135.880 1689.500 2136.140 1689.760 ;
        RECT 2142.320 1689.500 2142.580 1689.760 ;
        RECT 2112.880 1688.820 2113.140 1689.080 ;
        RECT 2134.960 1688.480 2135.220 1688.740 ;
        RECT 2142.320 20.100 2142.580 20.360 ;
        RECT 2554.020 20.100 2554.280 20.360 ;
      LAYER met2 ;
        RECT 2112.805 1700.000 2113.085 1704.000 ;
        RECT 2112.940 1689.110 2113.080 1700.000 ;
        RECT 2135.880 1689.470 2136.140 1689.790 ;
        RECT 2142.320 1689.470 2142.580 1689.790 ;
        RECT 2112.880 1688.790 2113.140 1689.110 ;
        RECT 2134.960 1688.450 2135.220 1688.770 ;
        RECT 2135.020 1688.170 2135.160 1688.450 ;
        RECT 2135.940 1688.170 2136.080 1689.470 ;
        RECT 2135.020 1688.030 2136.080 1688.170 ;
        RECT 2142.380 20.390 2142.520 1689.470 ;
        RECT 2142.320 20.070 2142.580 20.390 ;
        RECT 2554.020 20.070 2554.280 20.390 ;
        RECT 2554.080 2.400 2554.220 20.070 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2162.605 1689.205 2162.775 1690.395 ;
      LAYER mcon ;
        RECT 2162.605 1690.225 2162.775 1690.395 ;
      LAYER met1 ;
        RECT 2162.545 1690.380 2162.835 1690.425 ;
        RECT 2514.890 1690.380 2515.210 1690.440 ;
        RECT 2162.545 1690.240 2515.210 1690.380 ;
        RECT 2162.545 1690.195 2162.835 1690.240 ;
        RECT 2514.890 1690.180 2515.210 1690.240 ;
        RECT 2119.290 1689.360 2119.610 1689.420 ;
        RECT 2162.545 1689.360 2162.835 1689.405 ;
        RECT 2119.290 1689.220 2162.835 1689.360 ;
        RECT 2119.290 1689.160 2119.610 1689.220 ;
        RECT 2162.545 1689.175 2162.835 1689.220 ;
        RECT 2571.930 16.900 2572.250 16.960 ;
        RECT 2536.600 16.760 2572.250 16.900 ;
        RECT 2514.890 16.220 2515.210 16.280 ;
        RECT 2536.600 16.220 2536.740 16.760 ;
        RECT 2571.930 16.700 2572.250 16.760 ;
        RECT 2514.890 16.080 2536.740 16.220 ;
        RECT 2514.890 16.020 2515.210 16.080 ;
      LAYER via ;
        RECT 2514.920 1690.180 2515.180 1690.440 ;
        RECT 2119.320 1689.160 2119.580 1689.420 ;
        RECT 2514.920 16.020 2515.180 16.280 ;
        RECT 2571.960 16.700 2572.220 16.960 ;
      LAYER met2 ;
        RECT 2119.245 1700.000 2119.525 1704.000 ;
        RECT 2119.380 1689.450 2119.520 1700.000 ;
        RECT 2514.920 1690.150 2515.180 1690.470 ;
        RECT 2119.320 1689.130 2119.580 1689.450 ;
        RECT 2514.980 16.310 2515.120 1690.150 ;
        RECT 2571.960 16.670 2572.220 16.990 ;
        RECT 2514.920 15.990 2515.180 16.310 ;
        RECT 2572.020 2.400 2572.160 16.670 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2126.190 1688.340 2126.510 1688.400 ;
        RECT 2149.190 1688.340 2149.510 1688.400 ;
        RECT 2126.190 1688.200 2149.510 1688.340 ;
        RECT 2126.190 1688.140 2126.510 1688.200 ;
        RECT 2149.190 1688.140 2149.510 1688.200 ;
        RECT 2149.190 19.960 2149.510 20.020 ;
        RECT 2589.410 19.960 2589.730 20.020 ;
        RECT 2149.190 19.820 2589.730 19.960 ;
        RECT 2149.190 19.760 2149.510 19.820 ;
        RECT 2589.410 19.760 2589.730 19.820 ;
      LAYER via ;
        RECT 2126.220 1688.140 2126.480 1688.400 ;
        RECT 2149.220 1688.140 2149.480 1688.400 ;
        RECT 2149.220 19.760 2149.480 20.020 ;
        RECT 2589.440 19.760 2589.700 20.020 ;
      LAYER met2 ;
        RECT 2126.145 1700.000 2126.425 1704.000 ;
        RECT 2126.280 1688.430 2126.420 1700.000 ;
        RECT 2126.220 1688.110 2126.480 1688.430 ;
        RECT 2149.220 1688.110 2149.480 1688.430 ;
        RECT 2149.280 20.050 2149.420 1688.110 ;
        RECT 2149.220 19.730 2149.480 20.050 ;
        RECT 2589.440 19.730 2589.700 20.050 ;
        RECT 2589.500 2.400 2589.640 19.730 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 823.470 35.260 823.790 35.320 ;
        RECT 1456.430 35.260 1456.750 35.320 ;
        RECT 823.470 35.120 1456.750 35.260 ;
        RECT 823.470 35.060 823.790 35.120 ;
        RECT 1456.430 35.060 1456.750 35.120 ;
      LAYER via ;
        RECT 823.500 35.060 823.760 35.320 ;
        RECT 1456.460 35.060 1456.720 35.320 ;
      LAYER met2 ;
        RECT 1459.605 1700.410 1459.885 1704.000 ;
        RECT 1457.900 1700.270 1459.885 1700.410 ;
        RECT 1457.900 1677.970 1458.040 1700.270 ;
        RECT 1459.605 1700.000 1459.885 1700.270 ;
        RECT 1456.520 1677.830 1458.040 1677.970 ;
        RECT 1456.520 35.350 1456.660 1677.830 ;
        RECT 823.500 35.030 823.760 35.350 ;
        RECT 1456.460 35.030 1456.720 35.350 ;
        RECT 823.560 2.400 823.700 35.030 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2535.590 1689.700 2535.910 1689.760 ;
        RECT 2163.080 1689.560 2535.910 1689.700 ;
        RECT 2133.090 1689.020 2133.410 1689.080 ;
        RECT 2163.080 1689.020 2163.220 1689.560 ;
        RECT 2535.590 1689.500 2535.910 1689.560 ;
        RECT 2133.090 1688.880 2163.220 1689.020 ;
        RECT 2133.090 1688.820 2133.410 1688.880 ;
        RECT 2535.590 20.640 2535.910 20.700 ;
        RECT 2607.350 20.640 2607.670 20.700 ;
        RECT 2535.590 20.500 2607.670 20.640 ;
        RECT 2535.590 20.440 2535.910 20.500 ;
        RECT 2607.350 20.440 2607.670 20.500 ;
      LAYER via ;
        RECT 2133.120 1688.820 2133.380 1689.080 ;
        RECT 2535.620 1689.500 2535.880 1689.760 ;
        RECT 2535.620 20.440 2535.880 20.700 ;
        RECT 2607.380 20.440 2607.640 20.700 ;
      LAYER met2 ;
        RECT 2133.045 1700.000 2133.325 1704.000 ;
        RECT 2133.180 1689.110 2133.320 1700.000 ;
        RECT 2535.620 1689.470 2535.880 1689.790 ;
        RECT 2133.120 1688.790 2133.380 1689.110 ;
        RECT 2535.680 20.730 2535.820 1689.470 ;
        RECT 2535.620 20.410 2535.880 20.730 ;
        RECT 2607.380 20.410 2607.640 20.730 ;
        RECT 2607.440 2.400 2607.580 20.410 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2162.145 1689.545 2162.315 1690.395 ;
      LAYER mcon ;
        RECT 2162.145 1690.225 2162.315 1690.395 ;
      LAYER met1 ;
        RECT 2170.350 1690.720 2170.670 1690.780 ;
        RECT 2162.160 1690.580 2170.670 1690.720 ;
        RECT 2162.160 1690.425 2162.300 1690.580 ;
        RECT 2170.350 1690.520 2170.670 1690.580 ;
        RECT 2162.085 1690.195 2162.375 1690.425 ;
        RECT 2145.510 1689.700 2145.830 1689.760 ;
        RECT 2162.085 1689.700 2162.375 1689.745 ;
        RECT 2145.510 1689.560 2162.375 1689.700 ;
        RECT 2145.510 1689.500 2145.830 1689.560 ;
        RECT 2162.085 1689.515 2162.375 1689.560 ;
        RECT 2139.530 1688.680 2139.850 1688.740 ;
        RECT 2145.510 1688.680 2145.830 1688.740 ;
        RECT 2139.530 1688.540 2145.830 1688.680 ;
        RECT 2139.530 1688.480 2139.850 1688.540 ;
        RECT 2145.510 1688.480 2145.830 1688.540 ;
        RECT 2170.350 19.620 2170.670 19.680 ;
        RECT 2625.290 19.620 2625.610 19.680 ;
        RECT 2170.350 19.480 2625.610 19.620 ;
        RECT 2170.350 19.420 2170.670 19.480 ;
        RECT 2625.290 19.420 2625.610 19.480 ;
      LAYER via ;
        RECT 2170.380 1690.520 2170.640 1690.780 ;
        RECT 2145.540 1689.500 2145.800 1689.760 ;
        RECT 2139.560 1688.480 2139.820 1688.740 ;
        RECT 2145.540 1688.480 2145.800 1688.740 ;
        RECT 2170.380 19.420 2170.640 19.680 ;
        RECT 2625.320 19.420 2625.580 19.680 ;
      LAYER met2 ;
        RECT 2139.485 1700.000 2139.765 1704.000 ;
        RECT 2139.620 1688.770 2139.760 1700.000 ;
        RECT 2170.380 1690.490 2170.640 1690.810 ;
        RECT 2145.540 1689.470 2145.800 1689.790 ;
        RECT 2145.600 1688.770 2145.740 1689.470 ;
        RECT 2139.560 1688.450 2139.820 1688.770 ;
        RECT 2145.540 1688.450 2145.800 1688.770 ;
        RECT 2170.440 19.710 2170.580 1690.490 ;
        RECT 2170.380 19.390 2170.640 19.710 ;
        RECT 2625.320 19.390 2625.580 19.710 ;
        RECT 2625.380 2.400 2625.520 19.390 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2166.745 1688.185 2166.915 1689.035 ;
      LAYER mcon ;
        RECT 2166.745 1688.865 2166.915 1689.035 ;
      LAYER met1 ;
        RECT 2166.685 1689.020 2166.975 1689.065 ;
        RECT 2556.290 1689.020 2556.610 1689.080 ;
        RECT 2166.685 1688.880 2556.610 1689.020 ;
        RECT 2166.685 1688.835 2166.975 1688.880 ;
        RECT 2556.290 1688.820 2556.610 1688.880 ;
        RECT 2146.430 1688.680 2146.750 1688.740 ;
        RECT 2146.430 1688.540 2159.540 1688.680 ;
        RECT 2146.430 1688.480 2146.750 1688.540 ;
        RECT 2159.400 1688.340 2159.540 1688.540 ;
        RECT 2166.685 1688.340 2166.975 1688.385 ;
        RECT 2159.400 1688.200 2166.975 1688.340 ;
        RECT 2166.685 1688.155 2166.975 1688.200 ;
        RECT 2556.290 15.540 2556.610 15.600 ;
        RECT 2643.230 15.540 2643.550 15.600 ;
        RECT 2556.290 15.400 2643.550 15.540 ;
        RECT 2556.290 15.340 2556.610 15.400 ;
        RECT 2643.230 15.340 2643.550 15.400 ;
      LAYER via ;
        RECT 2556.320 1688.820 2556.580 1689.080 ;
        RECT 2146.460 1688.480 2146.720 1688.740 ;
        RECT 2556.320 15.340 2556.580 15.600 ;
        RECT 2643.260 15.340 2643.520 15.600 ;
      LAYER met2 ;
        RECT 2146.385 1700.000 2146.665 1704.000 ;
        RECT 2146.520 1688.770 2146.660 1700.000 ;
        RECT 2556.320 1688.790 2556.580 1689.110 ;
        RECT 2146.460 1688.450 2146.720 1688.770 ;
        RECT 2556.380 15.630 2556.520 1688.790 ;
        RECT 2556.320 15.310 2556.580 15.630 ;
        RECT 2643.260 15.310 2643.520 15.630 ;
        RECT 2643.320 2.400 2643.460 15.310 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2167.205 1688.185 2167.375 1691.075 ;
      LAYER mcon ;
        RECT 2167.205 1690.905 2167.375 1691.075 ;
      LAYER met1 ;
        RECT 2167.145 1691.060 2167.435 1691.105 ;
        RECT 2161.700 1690.920 2167.435 1691.060 ;
        RECT 2155.170 1690.720 2155.490 1690.780 ;
        RECT 2155.170 1690.580 2156.780 1690.720 ;
        RECT 2155.170 1690.520 2155.490 1690.580 ;
        RECT 2156.640 1690.380 2156.780 1690.580 ;
        RECT 2161.700 1690.380 2161.840 1690.920 ;
        RECT 2167.145 1690.875 2167.435 1690.920 ;
        RECT 2156.640 1690.240 2161.840 1690.380 ;
        RECT 2167.145 1688.340 2167.435 1688.385 ;
        RECT 2181.850 1688.340 2182.170 1688.400 ;
        RECT 2167.145 1688.200 2182.170 1688.340 ;
        RECT 2167.145 1688.155 2167.435 1688.200 ;
        RECT 2181.850 1688.140 2182.170 1688.200 ;
        RECT 2183.690 19.280 2184.010 19.340 ;
        RECT 2661.170 19.280 2661.490 19.340 ;
        RECT 2183.690 19.140 2661.490 19.280 ;
        RECT 2183.690 19.080 2184.010 19.140 ;
        RECT 2661.170 19.080 2661.490 19.140 ;
      LAYER via ;
        RECT 2155.200 1690.520 2155.460 1690.780 ;
        RECT 2181.880 1688.140 2182.140 1688.400 ;
        RECT 2183.720 19.080 2183.980 19.340 ;
        RECT 2661.200 19.080 2661.460 19.340 ;
      LAYER met2 ;
        RECT 2153.285 1700.410 2153.565 1704.000 ;
        RECT 2153.285 1700.270 2155.400 1700.410 ;
        RECT 2153.285 1700.000 2153.565 1700.270 ;
        RECT 2155.260 1690.810 2155.400 1700.270 ;
        RECT 2155.200 1690.490 2155.460 1690.810 ;
        RECT 2181.880 1688.110 2182.140 1688.430 ;
        RECT 2181.940 1677.970 2182.080 1688.110 ;
        RECT 2181.940 1677.830 2183.920 1677.970 ;
        RECT 2183.780 19.370 2183.920 1677.830 ;
        RECT 2183.720 19.050 2183.980 19.370 ;
        RECT 2661.200 19.050 2661.460 19.370 ;
        RECT 2661.260 2.400 2661.400 19.050 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2185.145 1687.165 2185.315 1688.695 ;
        RECT 2211.365 1687.165 2211.535 1689.375 ;
      LAYER mcon ;
        RECT 2211.365 1689.205 2211.535 1689.375 ;
        RECT 2185.145 1688.525 2185.315 1688.695 ;
      LAYER met1 ;
        RECT 2211.305 1689.360 2211.595 1689.405 ;
        RECT 2570.090 1689.360 2570.410 1689.420 ;
        RECT 2211.305 1689.220 2570.410 1689.360 ;
        RECT 2211.305 1689.175 2211.595 1689.220 ;
        RECT 2570.090 1689.160 2570.410 1689.220 ;
        RECT 2159.770 1688.680 2160.090 1688.740 ;
        RECT 2185.085 1688.680 2185.375 1688.725 ;
        RECT 2159.770 1688.540 2185.375 1688.680 ;
        RECT 2159.770 1688.480 2160.090 1688.540 ;
        RECT 2185.085 1688.495 2185.375 1688.540 ;
        RECT 2185.085 1687.320 2185.375 1687.365 ;
        RECT 2211.305 1687.320 2211.595 1687.365 ;
        RECT 2185.085 1687.180 2211.595 1687.320 ;
        RECT 2185.085 1687.135 2185.375 1687.180 ;
        RECT 2211.305 1687.135 2211.595 1687.180 ;
        RECT 2570.090 15.880 2570.410 15.940 ;
        RECT 2678.650 15.880 2678.970 15.940 ;
        RECT 2570.090 15.740 2678.970 15.880 ;
        RECT 2570.090 15.680 2570.410 15.740 ;
        RECT 2678.650 15.680 2678.970 15.740 ;
      LAYER via ;
        RECT 2570.120 1689.160 2570.380 1689.420 ;
        RECT 2159.800 1688.480 2160.060 1688.740 ;
        RECT 2570.120 15.680 2570.380 15.940 ;
        RECT 2678.680 15.680 2678.940 15.940 ;
      LAYER met2 ;
        RECT 2159.725 1700.000 2160.005 1704.000 ;
        RECT 2159.860 1688.770 2160.000 1700.000 ;
        RECT 2570.120 1689.130 2570.380 1689.450 ;
        RECT 2159.800 1688.450 2160.060 1688.770 ;
        RECT 2570.180 15.970 2570.320 1689.130 ;
        RECT 2570.120 15.650 2570.380 15.970 ;
        RECT 2678.680 15.650 2678.940 15.970 ;
        RECT 2678.740 2.400 2678.880 15.650 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2176.405 1256.385 2176.575 1304.155 ;
        RECT 2175.485 1207.425 2175.655 1255.875 ;
        RECT 2175.485 1110.865 2175.655 1124.975 ;
        RECT 2175.945 379.525 2176.115 427.635 ;
        RECT 2175.945 255.085 2176.115 331.075 ;
        RECT 2176.405 193.205 2176.575 241.315 ;
        RECT 2176.405 96.645 2176.575 144.755 ;
      LAYER mcon ;
        RECT 2176.405 1303.985 2176.575 1304.155 ;
        RECT 2175.485 1255.705 2175.655 1255.875 ;
        RECT 2175.485 1124.805 2175.655 1124.975 ;
        RECT 2175.945 427.465 2176.115 427.635 ;
        RECT 2175.945 330.905 2176.115 331.075 ;
        RECT 2176.405 241.145 2176.575 241.315 ;
        RECT 2176.405 144.585 2176.575 144.755 ;
      LAYER met1 ;
        RECT 2166.670 1687.320 2166.990 1687.380 ;
        RECT 2175.410 1687.320 2175.730 1687.380 ;
        RECT 2166.670 1687.180 2175.730 1687.320 ;
        RECT 2166.670 1687.120 2166.990 1687.180 ;
        RECT 2175.410 1687.120 2175.730 1687.180 ;
        RECT 2176.790 1583.620 2177.110 1583.680 ;
        RECT 2177.710 1583.620 2178.030 1583.680 ;
        RECT 2176.790 1583.480 2178.030 1583.620 ;
        RECT 2176.790 1583.420 2177.110 1583.480 ;
        RECT 2177.710 1583.420 2178.030 1583.480 ;
        RECT 2176.790 1511.200 2177.110 1511.260 ;
        RECT 2177.710 1511.200 2178.030 1511.260 ;
        RECT 2176.790 1511.060 2178.030 1511.200 ;
        RECT 2176.790 1511.000 2177.110 1511.060 ;
        RECT 2177.710 1511.000 2178.030 1511.060 ;
        RECT 2176.790 1487.060 2177.110 1487.120 ;
        RECT 2177.710 1487.060 2178.030 1487.120 ;
        RECT 2176.790 1486.920 2178.030 1487.060 ;
        RECT 2176.790 1486.860 2177.110 1486.920 ;
        RECT 2177.710 1486.860 2178.030 1486.920 ;
        RECT 2176.790 1414.640 2177.110 1414.700 ;
        RECT 2177.710 1414.640 2178.030 1414.700 ;
        RECT 2176.790 1414.500 2178.030 1414.640 ;
        RECT 2176.790 1414.440 2177.110 1414.500 ;
        RECT 2177.710 1414.440 2178.030 1414.500 ;
        RECT 2176.790 1390.500 2177.110 1390.560 ;
        RECT 2177.710 1390.500 2178.030 1390.560 ;
        RECT 2176.790 1390.360 2178.030 1390.500 ;
        RECT 2176.790 1390.300 2177.110 1390.360 ;
        RECT 2177.710 1390.300 2178.030 1390.360 ;
        RECT 2176.790 1318.080 2177.110 1318.140 ;
        RECT 2177.710 1318.080 2178.030 1318.140 ;
        RECT 2176.790 1317.940 2178.030 1318.080 ;
        RECT 2176.790 1317.880 2177.110 1317.940 ;
        RECT 2177.710 1317.880 2178.030 1317.940 ;
        RECT 2176.330 1304.140 2176.650 1304.200 ;
        RECT 2176.135 1304.000 2176.650 1304.140 ;
        RECT 2176.330 1303.940 2176.650 1304.000 ;
        RECT 2176.330 1256.540 2176.650 1256.600 ;
        RECT 2176.135 1256.400 2176.650 1256.540 ;
        RECT 2176.330 1256.340 2176.650 1256.400 ;
        RECT 2175.425 1255.860 2175.715 1255.905 ;
        RECT 2175.870 1255.860 2176.190 1255.920 ;
        RECT 2175.425 1255.720 2176.190 1255.860 ;
        RECT 2175.425 1255.675 2175.715 1255.720 ;
        RECT 2175.870 1255.660 2176.190 1255.720 ;
        RECT 2175.410 1207.580 2175.730 1207.640 ;
        RECT 2175.215 1207.440 2175.730 1207.580 ;
        RECT 2175.410 1207.380 2175.730 1207.440 ;
        RECT 2175.410 1173.040 2175.730 1173.300 ;
        RECT 2175.500 1172.560 2175.640 1173.040 ;
        RECT 2175.870 1172.560 2176.190 1172.620 ;
        RECT 2175.500 1172.420 2176.190 1172.560 ;
        RECT 2175.870 1172.360 2176.190 1172.420 ;
        RECT 2175.410 1124.960 2175.730 1125.020 ;
        RECT 2175.215 1124.820 2175.730 1124.960 ;
        RECT 2175.410 1124.760 2175.730 1124.820 ;
        RECT 2175.410 1111.020 2175.730 1111.080 ;
        RECT 2175.215 1110.880 2175.730 1111.020 ;
        RECT 2175.410 1110.820 2175.730 1110.880 ;
        RECT 2175.410 1076.480 2175.730 1076.740 ;
        RECT 2175.500 1076.000 2175.640 1076.480 ;
        RECT 2175.870 1076.000 2176.190 1076.060 ;
        RECT 2175.500 1075.860 2176.190 1076.000 ;
        RECT 2175.870 1075.800 2176.190 1075.860 ;
        RECT 2175.870 979.440 2176.190 979.500 ;
        RECT 2176.790 979.440 2177.110 979.500 ;
        RECT 2175.870 979.300 2177.110 979.440 ;
        RECT 2175.870 979.240 2176.190 979.300 ;
        RECT 2176.790 979.240 2177.110 979.300 ;
        RECT 2175.870 835.280 2176.190 835.340 ;
        RECT 2176.790 835.280 2177.110 835.340 ;
        RECT 2175.870 835.140 2177.110 835.280 ;
        RECT 2175.870 835.080 2176.190 835.140 ;
        RECT 2176.790 835.080 2177.110 835.140 ;
        RECT 2175.870 825.420 2176.190 825.480 ;
        RECT 2177.710 825.420 2178.030 825.480 ;
        RECT 2175.870 825.280 2178.030 825.420 ;
        RECT 2175.870 825.220 2176.190 825.280 ;
        RECT 2177.710 825.220 2178.030 825.280 ;
        RECT 2177.710 738.860 2178.030 739.120 ;
        RECT 2177.800 738.100 2177.940 738.860 ;
        RECT 2177.710 737.840 2178.030 738.100 ;
        RECT 2176.790 690.100 2177.110 690.160 ;
        RECT 2177.710 690.100 2178.030 690.160 ;
        RECT 2176.790 689.960 2178.030 690.100 ;
        RECT 2176.790 689.900 2177.110 689.960 ;
        RECT 2177.710 689.900 2178.030 689.960 ;
        RECT 2176.790 627.880 2177.110 627.940 ;
        RECT 2177.710 627.880 2178.030 627.940 ;
        RECT 2176.790 627.740 2178.030 627.880 ;
        RECT 2176.790 627.680 2177.110 627.740 ;
        RECT 2177.710 627.680 2178.030 627.740 ;
        RECT 2176.790 545.260 2177.110 545.320 ;
        RECT 2177.710 545.260 2178.030 545.320 ;
        RECT 2176.790 545.120 2178.030 545.260 ;
        RECT 2176.790 545.060 2177.110 545.120 ;
        RECT 2177.710 545.060 2178.030 545.120 ;
        RECT 2175.870 427.620 2176.190 427.680 ;
        RECT 2175.675 427.480 2176.190 427.620 ;
        RECT 2175.870 427.420 2176.190 427.480 ;
        RECT 2175.870 379.680 2176.190 379.740 ;
        RECT 2175.675 379.540 2176.190 379.680 ;
        RECT 2175.870 379.480 2176.190 379.540 ;
        RECT 2175.870 338.680 2176.190 338.940 ;
        RECT 2175.960 338.260 2176.100 338.680 ;
        RECT 2175.870 338.000 2176.190 338.260 ;
        RECT 2175.870 331.060 2176.190 331.120 ;
        RECT 2175.675 330.920 2176.190 331.060 ;
        RECT 2175.870 330.860 2176.190 330.920 ;
        RECT 2175.870 255.240 2176.190 255.300 ;
        RECT 2175.675 255.100 2176.190 255.240 ;
        RECT 2175.870 255.040 2176.190 255.100 ;
        RECT 2176.330 241.300 2176.650 241.360 ;
        RECT 2176.135 241.160 2176.650 241.300 ;
        RECT 2176.330 241.100 2176.650 241.160 ;
        RECT 2176.345 193.360 2176.635 193.405 ;
        RECT 2176.790 193.360 2177.110 193.420 ;
        RECT 2176.345 193.220 2177.110 193.360 ;
        RECT 2176.345 193.175 2176.635 193.220 ;
        RECT 2176.790 193.160 2177.110 193.220 ;
        RECT 2176.345 144.740 2176.635 144.785 ;
        RECT 2176.790 144.740 2177.110 144.800 ;
        RECT 2176.345 144.600 2177.110 144.740 ;
        RECT 2176.345 144.555 2176.635 144.600 ;
        RECT 2176.790 144.540 2177.110 144.600 ;
        RECT 2176.330 96.800 2176.650 96.860 ;
        RECT 2176.135 96.660 2176.650 96.800 ;
        RECT 2176.330 96.600 2176.650 96.660 ;
        RECT 2175.870 18.940 2176.190 19.000 ;
        RECT 2696.590 18.940 2696.910 19.000 ;
        RECT 2175.870 18.800 2696.910 18.940 ;
        RECT 2175.870 18.740 2176.190 18.800 ;
        RECT 2696.590 18.740 2696.910 18.800 ;
      LAYER via ;
        RECT 2166.700 1687.120 2166.960 1687.380 ;
        RECT 2175.440 1687.120 2175.700 1687.380 ;
        RECT 2176.820 1583.420 2177.080 1583.680 ;
        RECT 2177.740 1583.420 2178.000 1583.680 ;
        RECT 2176.820 1511.000 2177.080 1511.260 ;
        RECT 2177.740 1511.000 2178.000 1511.260 ;
        RECT 2176.820 1486.860 2177.080 1487.120 ;
        RECT 2177.740 1486.860 2178.000 1487.120 ;
        RECT 2176.820 1414.440 2177.080 1414.700 ;
        RECT 2177.740 1414.440 2178.000 1414.700 ;
        RECT 2176.820 1390.300 2177.080 1390.560 ;
        RECT 2177.740 1390.300 2178.000 1390.560 ;
        RECT 2176.820 1317.880 2177.080 1318.140 ;
        RECT 2177.740 1317.880 2178.000 1318.140 ;
        RECT 2176.360 1303.940 2176.620 1304.200 ;
        RECT 2176.360 1256.340 2176.620 1256.600 ;
        RECT 2175.900 1255.660 2176.160 1255.920 ;
        RECT 2175.440 1207.380 2175.700 1207.640 ;
        RECT 2175.440 1173.040 2175.700 1173.300 ;
        RECT 2175.900 1172.360 2176.160 1172.620 ;
        RECT 2175.440 1124.760 2175.700 1125.020 ;
        RECT 2175.440 1110.820 2175.700 1111.080 ;
        RECT 2175.440 1076.480 2175.700 1076.740 ;
        RECT 2175.900 1075.800 2176.160 1076.060 ;
        RECT 2175.900 979.240 2176.160 979.500 ;
        RECT 2176.820 979.240 2177.080 979.500 ;
        RECT 2175.900 835.080 2176.160 835.340 ;
        RECT 2176.820 835.080 2177.080 835.340 ;
        RECT 2175.900 825.220 2176.160 825.480 ;
        RECT 2177.740 825.220 2178.000 825.480 ;
        RECT 2177.740 738.860 2178.000 739.120 ;
        RECT 2177.740 737.840 2178.000 738.100 ;
        RECT 2176.820 689.900 2177.080 690.160 ;
        RECT 2177.740 689.900 2178.000 690.160 ;
        RECT 2176.820 627.680 2177.080 627.940 ;
        RECT 2177.740 627.680 2178.000 627.940 ;
        RECT 2176.820 545.060 2177.080 545.320 ;
        RECT 2177.740 545.060 2178.000 545.320 ;
        RECT 2175.900 427.420 2176.160 427.680 ;
        RECT 2175.900 379.480 2176.160 379.740 ;
        RECT 2175.900 338.680 2176.160 338.940 ;
        RECT 2175.900 338.000 2176.160 338.260 ;
        RECT 2175.900 330.860 2176.160 331.120 ;
        RECT 2175.900 255.040 2176.160 255.300 ;
        RECT 2176.360 241.100 2176.620 241.360 ;
        RECT 2176.820 193.160 2177.080 193.420 ;
        RECT 2176.820 144.540 2177.080 144.800 ;
        RECT 2176.360 96.600 2176.620 96.860 ;
        RECT 2175.900 18.740 2176.160 19.000 ;
        RECT 2696.620 18.740 2696.880 19.000 ;
      LAYER met2 ;
        RECT 2166.625 1700.000 2166.905 1704.000 ;
        RECT 2166.760 1687.410 2166.900 1700.000 ;
        RECT 2166.700 1687.090 2166.960 1687.410 ;
        RECT 2175.440 1687.090 2175.700 1687.410 ;
        RECT 2175.500 1607.930 2175.640 1687.090 ;
        RECT 2175.500 1607.790 2177.020 1607.930 ;
        RECT 2176.880 1583.710 2177.020 1607.790 ;
        RECT 2176.820 1583.390 2177.080 1583.710 ;
        RECT 2177.740 1583.390 2178.000 1583.710 ;
        RECT 2177.800 1511.290 2177.940 1583.390 ;
        RECT 2176.820 1510.970 2177.080 1511.290 ;
        RECT 2177.740 1510.970 2178.000 1511.290 ;
        RECT 2176.880 1487.150 2177.020 1510.970 ;
        RECT 2176.820 1486.830 2177.080 1487.150 ;
        RECT 2177.740 1486.830 2178.000 1487.150 ;
        RECT 2177.800 1414.730 2177.940 1486.830 ;
        RECT 2176.820 1414.410 2177.080 1414.730 ;
        RECT 2177.740 1414.410 2178.000 1414.730 ;
        RECT 2176.880 1390.590 2177.020 1414.410 ;
        RECT 2176.820 1390.270 2177.080 1390.590 ;
        RECT 2177.740 1390.270 2178.000 1390.590 ;
        RECT 2177.800 1318.170 2177.940 1390.270 ;
        RECT 2176.820 1317.850 2177.080 1318.170 ;
        RECT 2177.740 1317.850 2178.000 1318.170 ;
        RECT 2176.880 1317.570 2177.020 1317.850 ;
        RECT 2176.420 1317.430 2177.020 1317.570 ;
        RECT 2176.420 1304.230 2176.560 1317.430 ;
        RECT 2176.360 1303.910 2176.620 1304.230 ;
        RECT 2176.360 1256.370 2176.620 1256.630 ;
        RECT 2175.960 1256.310 2176.620 1256.370 ;
        RECT 2175.960 1256.230 2176.560 1256.310 ;
        RECT 2175.960 1255.950 2176.100 1256.230 ;
        RECT 2175.900 1255.630 2176.160 1255.950 ;
        RECT 2175.440 1207.350 2175.700 1207.670 ;
        RECT 2175.500 1173.330 2175.640 1207.350 ;
        RECT 2175.440 1173.010 2175.700 1173.330 ;
        RECT 2175.900 1172.330 2176.160 1172.650 ;
        RECT 2175.960 1159.130 2176.100 1172.330 ;
        RECT 2175.500 1158.990 2176.100 1159.130 ;
        RECT 2175.500 1125.050 2175.640 1158.990 ;
        RECT 2175.440 1124.730 2175.700 1125.050 ;
        RECT 2175.440 1110.790 2175.700 1111.110 ;
        RECT 2175.500 1076.770 2175.640 1110.790 ;
        RECT 2175.440 1076.450 2175.700 1076.770 ;
        RECT 2175.900 1075.770 2176.160 1076.090 ;
        RECT 2175.960 1062.685 2176.100 1075.770 ;
        RECT 2175.890 1062.315 2176.170 1062.685 ;
        RECT 2176.810 1062.315 2177.090 1062.685 ;
        RECT 2176.880 1014.460 2177.020 1062.315 ;
        RECT 2175.960 1014.405 2177.020 1014.460 ;
        RECT 2175.890 1014.320 2177.090 1014.405 ;
        RECT 2175.890 1014.035 2176.170 1014.320 ;
        RECT 2176.810 1014.035 2177.090 1014.320 ;
        RECT 2176.880 979.530 2177.020 1014.035 ;
        RECT 2175.900 979.210 2176.160 979.530 ;
        RECT 2176.820 979.210 2177.080 979.530 ;
        RECT 2175.960 931.330 2176.100 979.210 ;
        RECT 2175.960 931.190 2177.020 931.330 ;
        RECT 2176.880 835.370 2177.020 931.190 ;
        RECT 2175.900 835.050 2176.160 835.370 ;
        RECT 2176.820 835.050 2177.080 835.370 ;
        RECT 2175.960 825.510 2176.100 835.050 ;
        RECT 2175.900 825.190 2176.160 825.510 ;
        RECT 2177.740 825.190 2178.000 825.510 ;
        RECT 2177.800 739.150 2177.940 825.190 ;
        RECT 2177.740 738.830 2178.000 739.150 ;
        RECT 2177.740 737.810 2178.000 738.130 ;
        RECT 2177.800 690.190 2177.940 737.810 ;
        RECT 2176.820 689.870 2177.080 690.190 ;
        RECT 2177.740 689.870 2178.000 690.190 ;
        RECT 2176.880 627.970 2177.020 689.870 ;
        RECT 2176.820 627.650 2177.080 627.970 ;
        RECT 2177.740 627.650 2178.000 627.970 ;
        RECT 2177.800 545.350 2177.940 627.650 ;
        RECT 2176.820 545.090 2177.080 545.350 ;
        RECT 2176.420 545.030 2177.080 545.090 ;
        RECT 2177.740 545.030 2178.000 545.350 ;
        RECT 2176.420 544.950 2177.020 545.030 ;
        RECT 2176.420 497.490 2176.560 544.950 ;
        RECT 2176.420 497.350 2177.020 497.490 ;
        RECT 2176.880 496.130 2177.020 497.350 ;
        RECT 2175.960 495.990 2177.020 496.130 ;
        RECT 2175.960 435.725 2176.100 495.990 ;
        RECT 2175.890 435.355 2176.170 435.725 ;
        RECT 2175.890 434.675 2176.170 435.045 ;
        RECT 2175.960 427.710 2176.100 434.675 ;
        RECT 2175.900 427.390 2176.160 427.710 ;
        RECT 2175.900 379.450 2176.160 379.770 ;
        RECT 2175.960 338.970 2176.100 379.450 ;
        RECT 2175.900 338.650 2176.160 338.970 ;
        RECT 2175.900 337.970 2176.160 338.290 ;
        RECT 2175.960 331.150 2176.100 337.970 ;
        RECT 2175.900 330.830 2176.160 331.150 ;
        RECT 2175.900 255.010 2176.160 255.330 ;
        RECT 2175.960 241.810 2176.100 255.010 ;
        RECT 2175.960 241.670 2176.560 241.810 ;
        RECT 2176.420 241.390 2176.560 241.670 ;
        RECT 2176.360 241.070 2176.620 241.390 ;
        RECT 2176.820 193.130 2177.080 193.450 ;
        RECT 2176.880 144.830 2177.020 193.130 ;
        RECT 2176.820 144.510 2177.080 144.830 ;
        RECT 2176.360 96.570 2176.620 96.890 ;
        RECT 2176.420 62.290 2176.560 96.570 ;
        RECT 2175.960 62.150 2176.560 62.290 ;
        RECT 2175.960 19.030 2176.100 62.150 ;
        RECT 2175.900 18.710 2176.160 19.030 ;
        RECT 2696.620 18.710 2696.880 19.030 ;
        RECT 2696.680 2.400 2696.820 18.710 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 2175.890 1062.360 2176.170 1062.640 ;
        RECT 2176.810 1062.360 2177.090 1062.640 ;
        RECT 2175.890 1014.080 2176.170 1014.360 ;
        RECT 2176.810 1014.080 2177.090 1014.360 ;
        RECT 2175.890 435.400 2176.170 435.680 ;
        RECT 2175.890 434.720 2176.170 435.000 ;
      LAYER met3 ;
        RECT 2175.865 1062.650 2176.195 1062.665 ;
        RECT 2176.785 1062.650 2177.115 1062.665 ;
        RECT 2175.865 1062.350 2177.115 1062.650 ;
        RECT 2175.865 1062.335 2176.195 1062.350 ;
        RECT 2176.785 1062.335 2177.115 1062.350 ;
        RECT 2175.865 1014.370 2176.195 1014.385 ;
        RECT 2176.785 1014.370 2177.115 1014.385 ;
        RECT 2175.865 1014.070 2177.115 1014.370 ;
        RECT 2175.865 1014.055 2176.195 1014.070 ;
        RECT 2176.785 1014.055 2177.115 1014.070 ;
        RECT 2175.865 435.690 2176.195 435.705 ;
        RECT 2175.865 435.375 2176.410 435.690 ;
        RECT 2176.110 435.025 2176.410 435.375 ;
        RECT 2175.865 434.710 2176.410 435.025 ;
        RECT 2175.865 434.695 2176.195 434.710 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2590.790 1688.680 2591.110 1688.740 ;
        RECT 2235.760 1688.540 2591.110 1688.680 ;
        RECT 2191.050 1688.000 2191.370 1688.060 ;
        RECT 2235.760 1688.000 2235.900 1688.540 ;
        RECT 2590.790 1688.480 2591.110 1688.540 ;
        RECT 2191.050 1687.860 2235.900 1688.000 ;
        RECT 2191.050 1687.800 2191.370 1687.860 ;
        RECT 2590.790 16.220 2591.110 16.280 ;
        RECT 2714.530 16.220 2714.850 16.280 ;
        RECT 2590.790 16.080 2714.850 16.220 ;
        RECT 2590.790 16.020 2591.110 16.080 ;
        RECT 2714.530 16.020 2714.850 16.080 ;
      LAYER via ;
        RECT 2191.080 1687.800 2191.340 1688.060 ;
        RECT 2590.820 1688.480 2591.080 1688.740 ;
        RECT 2590.820 16.020 2591.080 16.280 ;
        RECT 2714.560 16.020 2714.820 16.280 ;
      LAYER met2 ;
        RECT 2173.525 1700.410 2173.805 1704.000 ;
        RECT 2173.525 1700.270 2175.180 1700.410 ;
        RECT 2173.525 1700.000 2173.805 1700.270 ;
        RECT 2175.040 1689.645 2175.180 1700.270 ;
        RECT 2174.970 1689.275 2175.250 1689.645 ;
        RECT 2191.070 1689.275 2191.350 1689.645 ;
        RECT 2191.140 1688.090 2191.280 1689.275 ;
        RECT 2590.820 1688.450 2591.080 1688.770 ;
        RECT 2191.080 1687.770 2191.340 1688.090 ;
        RECT 2590.880 16.310 2591.020 1688.450 ;
        RECT 2590.820 15.990 2591.080 16.310 ;
        RECT 2714.560 15.990 2714.820 16.310 ;
        RECT 2714.620 2.400 2714.760 15.990 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
      LAYER via2 ;
        RECT 2174.970 1689.320 2175.250 1689.600 ;
        RECT 2191.070 1689.320 2191.350 1689.600 ;
      LAYER met3 ;
        RECT 2174.945 1689.610 2175.275 1689.625 ;
        RECT 2191.045 1689.610 2191.375 1689.625 ;
        RECT 2174.945 1689.310 2191.375 1689.610 ;
        RECT 2174.945 1689.295 2175.275 1689.310 ;
        RECT 2191.045 1689.295 2191.375 1689.310 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 1686.980 2180.330 1687.040 ;
        RECT 2184.150 1686.980 2184.470 1687.040 ;
        RECT 2180.010 1686.840 2184.470 1686.980 ;
        RECT 2180.010 1686.780 2180.330 1686.840 ;
        RECT 2184.150 1686.780 2184.470 1686.840 ;
        RECT 2184.150 18.600 2184.470 18.660 ;
        RECT 2732.470 18.600 2732.790 18.660 ;
        RECT 2184.150 18.460 2732.790 18.600 ;
        RECT 2184.150 18.400 2184.470 18.460 ;
        RECT 2732.470 18.400 2732.790 18.460 ;
      LAYER via ;
        RECT 2180.040 1686.780 2180.300 1687.040 ;
        RECT 2184.180 1686.780 2184.440 1687.040 ;
        RECT 2184.180 18.400 2184.440 18.660 ;
        RECT 2732.500 18.400 2732.760 18.660 ;
      LAYER met2 ;
        RECT 2179.965 1700.000 2180.245 1704.000 ;
        RECT 2180.100 1687.070 2180.240 1700.000 ;
        RECT 2180.040 1686.750 2180.300 1687.070 ;
        RECT 2184.180 1686.750 2184.440 1687.070 ;
        RECT 2184.240 18.690 2184.380 1686.750 ;
        RECT 2184.180 18.370 2184.440 18.690 ;
        RECT 2732.500 18.370 2732.760 18.690 ;
        RECT 2732.560 2.400 2732.700 18.370 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2210.905 1687.505 2211.075 1689.375 ;
      LAYER mcon ;
        RECT 2210.905 1689.205 2211.075 1689.375 ;
      LAYER met1 ;
        RECT 2186.910 1689.360 2187.230 1689.420 ;
        RECT 2210.845 1689.360 2211.135 1689.405 ;
        RECT 2186.910 1689.220 2211.135 1689.360 ;
        RECT 2186.910 1689.160 2187.230 1689.220 ;
        RECT 2210.845 1689.175 2211.135 1689.220 ;
        RECT 2210.845 1687.660 2211.135 1687.705 ;
        RECT 2210.845 1687.520 2211.980 1687.660 ;
        RECT 2210.845 1687.475 2211.135 1687.520 ;
        RECT 2211.840 1687.320 2211.980 1687.520 ;
        RECT 2604.590 1687.320 2604.910 1687.380 ;
        RECT 2211.840 1687.180 2604.910 1687.320 ;
        RECT 2604.590 1687.120 2604.910 1687.180 ;
        RECT 2604.590 16.560 2604.910 16.620 ;
        RECT 2750.410 16.560 2750.730 16.620 ;
        RECT 2604.590 16.420 2750.730 16.560 ;
        RECT 2604.590 16.360 2604.910 16.420 ;
        RECT 2750.410 16.360 2750.730 16.420 ;
      LAYER via ;
        RECT 2186.940 1689.160 2187.200 1689.420 ;
        RECT 2604.620 1687.120 2604.880 1687.380 ;
        RECT 2604.620 16.360 2604.880 16.620 ;
        RECT 2750.440 16.360 2750.700 16.620 ;
      LAYER met2 ;
        RECT 2186.865 1700.000 2187.145 1704.000 ;
        RECT 2187.000 1689.450 2187.140 1700.000 ;
        RECT 2186.940 1689.130 2187.200 1689.450 ;
        RECT 2604.620 1687.090 2604.880 1687.410 ;
        RECT 2604.680 16.650 2604.820 1687.090 ;
        RECT 2604.620 16.330 2604.880 16.650 ;
        RECT 2750.440 16.330 2750.700 16.650 ;
        RECT 2750.500 2.400 2750.640 16.330 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2214.585 1687.505 2214.755 1688.695 ;
        RECT 2224.705 1687.675 2224.875 1688.355 ;
        RECT 2223.785 1687.505 2224.875 1687.675 ;
        RECT 2228.385 1686.825 2228.555 1688.355 ;
      LAYER mcon ;
        RECT 2214.585 1688.525 2214.755 1688.695 ;
        RECT 2224.705 1688.185 2224.875 1688.355 ;
        RECT 2228.385 1688.185 2228.555 1688.355 ;
      LAYER met1 ;
        RECT 2193.810 1688.680 2194.130 1688.740 ;
        RECT 2214.525 1688.680 2214.815 1688.725 ;
        RECT 2193.810 1688.540 2214.815 1688.680 ;
        RECT 2193.810 1688.480 2194.130 1688.540 ;
        RECT 2214.525 1688.495 2214.815 1688.540 ;
        RECT 2224.645 1688.340 2224.935 1688.385 ;
        RECT 2228.325 1688.340 2228.615 1688.385 ;
        RECT 2224.645 1688.200 2228.615 1688.340 ;
        RECT 2224.645 1688.155 2224.935 1688.200 ;
        RECT 2228.325 1688.155 2228.615 1688.200 ;
        RECT 2214.525 1687.660 2214.815 1687.705 ;
        RECT 2223.725 1687.660 2224.015 1687.705 ;
        RECT 2214.525 1687.520 2224.015 1687.660 ;
        RECT 2214.525 1687.475 2214.815 1687.520 ;
        RECT 2223.725 1687.475 2224.015 1687.520 ;
        RECT 2228.325 1686.980 2228.615 1687.025 ;
        RECT 2618.390 1686.980 2618.710 1687.040 ;
        RECT 2228.325 1686.840 2618.710 1686.980 ;
        RECT 2228.325 1686.795 2228.615 1686.840 ;
        RECT 2618.390 1686.780 2618.710 1686.840 ;
        RECT 2618.390 16.900 2618.710 16.960 ;
        RECT 2767.890 16.900 2768.210 16.960 ;
        RECT 2618.390 16.760 2768.210 16.900 ;
        RECT 2618.390 16.700 2618.710 16.760 ;
        RECT 2767.890 16.700 2768.210 16.760 ;
      LAYER via ;
        RECT 2193.840 1688.480 2194.100 1688.740 ;
        RECT 2618.420 1686.780 2618.680 1687.040 ;
        RECT 2618.420 16.700 2618.680 16.960 ;
        RECT 2767.920 16.700 2768.180 16.960 ;
      LAYER met2 ;
        RECT 2193.765 1700.000 2194.045 1704.000 ;
        RECT 2193.900 1688.770 2194.040 1700.000 ;
        RECT 2193.840 1688.450 2194.100 1688.770 ;
        RECT 2618.420 1686.750 2618.680 1687.070 ;
        RECT 2618.480 16.990 2618.620 1686.750 ;
        RECT 2618.420 16.670 2618.680 16.990 ;
        RECT 2767.920 16.670 2768.180 16.990 ;
        RECT 2767.980 2.400 2768.120 16.670 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 34.920 841.270 34.980 ;
        RECT 1463.330 34.920 1463.650 34.980 ;
        RECT 840.950 34.780 1463.650 34.920 ;
        RECT 840.950 34.720 841.270 34.780 ;
        RECT 1463.330 34.720 1463.650 34.780 ;
      LAYER via ;
        RECT 840.980 34.720 841.240 34.980 ;
        RECT 1463.360 34.720 1463.620 34.980 ;
      LAYER met2 ;
        RECT 1466.505 1700.410 1466.785 1704.000 ;
        RECT 1464.800 1700.270 1466.785 1700.410 ;
        RECT 1464.800 1678.140 1464.940 1700.270 ;
        RECT 1466.505 1700.000 1466.785 1700.270 ;
        RECT 1463.420 1678.000 1464.940 1678.140 ;
        RECT 1463.420 35.010 1463.560 1678.000 ;
        RECT 840.980 34.690 841.240 35.010 ;
        RECT 1463.360 34.690 1463.620 35.010 ;
        RECT 841.040 2.400 841.180 34.690 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2200.710 18.260 2201.030 18.320 ;
        RECT 2785.830 18.260 2786.150 18.320 ;
        RECT 2200.710 18.120 2786.150 18.260 ;
        RECT 2200.710 18.060 2201.030 18.120 ;
        RECT 2785.830 18.060 2786.150 18.120 ;
      LAYER via ;
        RECT 2200.740 18.060 2201.000 18.320 ;
        RECT 2785.860 18.060 2786.120 18.320 ;
      LAYER met2 ;
        RECT 2200.205 1700.410 2200.485 1704.000 ;
        RECT 2200.205 1700.270 2200.940 1700.410 ;
        RECT 2200.205 1700.000 2200.485 1700.270 ;
        RECT 2200.800 18.350 2200.940 1700.270 ;
        RECT 2200.740 18.030 2201.000 18.350 ;
        RECT 2785.860 18.030 2786.120 18.350 ;
        RECT 2785.920 2.400 2786.060 18.030 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2207.150 1688.340 2207.470 1688.400 ;
        RECT 2224.170 1688.340 2224.490 1688.400 ;
        RECT 2207.150 1688.200 2224.490 1688.340 ;
        RECT 2207.150 1688.140 2207.470 1688.200 ;
        RECT 2224.170 1688.140 2224.490 1688.200 ;
        RECT 2224.170 1687.660 2224.490 1687.720 ;
        RECT 2625.290 1687.660 2625.610 1687.720 ;
        RECT 2224.170 1687.520 2625.610 1687.660 ;
        RECT 2224.170 1687.460 2224.490 1687.520 ;
        RECT 2625.290 1687.460 2625.610 1687.520 ;
        RECT 2625.290 20.640 2625.610 20.700 ;
        RECT 2803.770 20.640 2804.090 20.700 ;
        RECT 2625.290 20.500 2804.090 20.640 ;
        RECT 2625.290 20.440 2625.610 20.500 ;
        RECT 2803.770 20.440 2804.090 20.500 ;
      LAYER via ;
        RECT 2207.180 1688.140 2207.440 1688.400 ;
        RECT 2224.200 1688.140 2224.460 1688.400 ;
        RECT 2224.200 1687.460 2224.460 1687.720 ;
        RECT 2625.320 1687.460 2625.580 1687.720 ;
        RECT 2625.320 20.440 2625.580 20.700 ;
        RECT 2803.800 20.440 2804.060 20.700 ;
      LAYER met2 ;
        RECT 2207.105 1700.000 2207.385 1704.000 ;
        RECT 2207.240 1688.430 2207.380 1700.000 ;
        RECT 2207.180 1688.110 2207.440 1688.430 ;
        RECT 2224.200 1688.110 2224.460 1688.430 ;
        RECT 2224.260 1687.750 2224.400 1688.110 ;
        RECT 2224.200 1687.430 2224.460 1687.750 ;
        RECT 2625.320 1687.430 2625.580 1687.750 ;
        RECT 2625.380 20.730 2625.520 1687.430 ;
        RECT 2625.320 20.410 2625.580 20.730 ;
        RECT 2803.800 20.410 2804.060 20.730 ;
        RECT 2803.860 2.400 2804.000 20.410 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.510 17.920 2214.830 17.980 ;
        RECT 2821.710 17.920 2822.030 17.980 ;
        RECT 2214.510 17.780 2822.030 17.920 ;
        RECT 2214.510 17.720 2214.830 17.780 ;
        RECT 2821.710 17.720 2822.030 17.780 ;
      LAYER via ;
        RECT 2214.540 17.720 2214.800 17.980 ;
        RECT 2821.740 17.720 2822.000 17.980 ;
      LAYER met2 ;
        RECT 2213.545 1700.410 2213.825 1704.000 ;
        RECT 2213.545 1700.270 2214.740 1700.410 ;
        RECT 2213.545 1700.000 2213.825 1700.270 ;
        RECT 2214.600 18.010 2214.740 1700.270 ;
        RECT 2214.540 17.690 2214.800 18.010 ;
        RECT 2821.740 17.690 2822.000 18.010 ;
        RECT 2821.800 2.400 2821.940 17.690 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2234.825 1683.935 2234.995 1688.695 ;
        RECT 2234.825 1683.765 2235.455 1683.935 ;
        RECT 2250.005 1683.765 2250.175 1688.015 ;
      LAYER mcon ;
        RECT 2234.825 1688.525 2234.995 1688.695 ;
        RECT 2250.005 1687.845 2250.175 1688.015 ;
        RECT 2235.285 1683.765 2235.455 1683.935 ;
      LAYER met1 ;
        RECT 2220.490 1688.680 2220.810 1688.740 ;
        RECT 2234.765 1688.680 2235.055 1688.725 ;
        RECT 2220.490 1688.540 2235.055 1688.680 ;
        RECT 2220.490 1688.480 2220.810 1688.540 ;
        RECT 2234.765 1688.495 2235.055 1688.540 ;
        RECT 2249.945 1688.000 2250.235 1688.045 ;
        RECT 2639.090 1688.000 2639.410 1688.060 ;
        RECT 2249.945 1687.860 2639.410 1688.000 ;
        RECT 2249.945 1687.815 2250.235 1687.860 ;
        RECT 2639.090 1687.800 2639.410 1687.860 ;
        RECT 2235.225 1683.920 2235.515 1683.965 ;
        RECT 2249.945 1683.920 2250.235 1683.965 ;
        RECT 2235.225 1683.780 2250.235 1683.920 ;
        RECT 2235.225 1683.735 2235.515 1683.780 ;
        RECT 2249.945 1683.735 2250.235 1683.780 ;
        RECT 2639.090 20.300 2639.410 20.360 ;
        RECT 2839.190 20.300 2839.510 20.360 ;
        RECT 2639.090 20.160 2839.510 20.300 ;
        RECT 2639.090 20.100 2639.410 20.160 ;
        RECT 2839.190 20.100 2839.510 20.160 ;
      LAYER via ;
        RECT 2220.520 1688.480 2220.780 1688.740 ;
        RECT 2639.120 1687.800 2639.380 1688.060 ;
        RECT 2639.120 20.100 2639.380 20.360 ;
        RECT 2839.220 20.100 2839.480 20.360 ;
      LAYER met2 ;
        RECT 2220.445 1700.000 2220.725 1704.000 ;
        RECT 2220.580 1688.770 2220.720 1700.000 ;
        RECT 2220.520 1688.450 2220.780 1688.770 ;
        RECT 2639.120 1687.770 2639.380 1688.090 ;
        RECT 2639.180 20.390 2639.320 1687.770 ;
        RECT 2639.120 20.070 2639.380 20.390 ;
        RECT 2839.220 20.070 2839.480 20.390 ;
        RECT 2839.280 2.400 2839.420 20.070 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2280.825 14.365 2280.995 17.595 ;
      LAYER mcon ;
        RECT 2280.825 17.425 2280.995 17.595 ;
      LAYER met1 ;
        RECT 2280.765 17.580 2281.055 17.625 ;
        RECT 2857.130 17.580 2857.450 17.640 ;
        RECT 2280.765 17.440 2857.450 17.580 ;
        RECT 2280.765 17.395 2281.055 17.440 ;
        RECT 2857.130 17.380 2857.450 17.440 ;
        RECT 2280.765 14.520 2281.055 14.565 ;
        RECT 2239.900 14.380 2281.055 14.520 ;
        RECT 2228.310 14.180 2228.630 14.240 ;
        RECT 2239.900 14.180 2240.040 14.380 ;
        RECT 2280.765 14.335 2281.055 14.380 ;
        RECT 2228.310 14.040 2240.040 14.180 ;
        RECT 2228.310 13.980 2228.630 14.040 ;
      LAYER via ;
        RECT 2857.160 17.380 2857.420 17.640 ;
        RECT 2228.340 13.980 2228.600 14.240 ;
      LAYER met2 ;
        RECT 2227.345 1700.410 2227.625 1704.000 ;
        RECT 2227.345 1700.270 2228.540 1700.410 ;
        RECT 2227.345 1700.000 2227.625 1700.270 ;
        RECT 2228.400 14.270 2228.540 1700.270 ;
        RECT 2857.160 17.350 2857.420 17.670 ;
        RECT 2228.340 13.950 2228.600 14.270 ;
        RECT 2857.220 2.400 2857.360 17.350 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2645.990 1688.340 2646.310 1688.400 ;
        RECT 2249.560 1688.200 2646.310 1688.340 ;
        RECT 2236.590 1688.000 2236.910 1688.060 ;
        RECT 2249.560 1688.000 2249.700 1688.200 ;
        RECT 2645.990 1688.140 2646.310 1688.200 ;
        RECT 2236.590 1687.860 2249.700 1688.000 ;
        RECT 2236.590 1687.800 2236.910 1687.860 ;
        RECT 2645.990 19.960 2646.310 20.020 ;
        RECT 2875.070 19.960 2875.390 20.020 ;
        RECT 2645.990 19.820 2875.390 19.960 ;
        RECT 2645.990 19.760 2646.310 19.820 ;
        RECT 2875.070 19.760 2875.390 19.820 ;
      LAYER via ;
        RECT 2236.620 1687.800 2236.880 1688.060 ;
        RECT 2646.020 1688.140 2646.280 1688.400 ;
        RECT 2646.020 19.760 2646.280 20.020 ;
        RECT 2875.100 19.760 2875.360 20.020 ;
      LAYER met2 ;
        RECT 2233.785 1700.410 2234.065 1704.000 ;
        RECT 2233.785 1700.270 2235.440 1700.410 ;
        RECT 2233.785 1700.000 2234.065 1700.270 ;
        RECT 2235.300 1689.530 2235.440 1700.270 ;
        RECT 2235.300 1689.390 2235.900 1689.530 ;
        RECT 2235.760 1687.490 2235.900 1689.390 ;
        RECT 2646.020 1688.110 2646.280 1688.430 ;
        RECT 2236.620 1687.770 2236.880 1688.090 ;
        RECT 2236.680 1687.490 2236.820 1687.770 ;
        RECT 2235.760 1687.350 2236.820 1687.490 ;
        RECT 2646.080 20.050 2646.220 1688.110 ;
        RECT 2646.020 19.730 2646.280 20.050 ;
        RECT 2875.100 19.730 2875.360 20.050 ;
        RECT 2875.160 2.400 2875.300 19.730 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2245.790 17.580 2246.110 17.640 ;
        RECT 2245.790 17.440 2280.520 17.580 ;
        RECT 2245.790 17.380 2246.110 17.440 ;
        RECT 2280.380 17.240 2280.520 17.440 ;
        RECT 2893.010 17.240 2893.330 17.300 ;
        RECT 2280.380 17.100 2893.330 17.240 ;
        RECT 2893.010 17.040 2893.330 17.100 ;
      LAYER via ;
        RECT 2245.820 17.380 2246.080 17.640 ;
        RECT 2893.040 17.040 2893.300 17.300 ;
      LAYER met2 ;
        RECT 2240.685 1700.000 2240.965 1704.000 ;
        RECT 2240.820 1688.965 2240.960 1700.000 ;
        RECT 2240.750 1688.595 2241.030 1688.965 ;
        RECT 2245.810 1688.595 2246.090 1688.965 ;
        RECT 2245.880 17.670 2246.020 1688.595 ;
        RECT 2245.820 17.350 2246.080 17.670 ;
        RECT 2893.040 17.010 2893.300 17.330 ;
        RECT 2893.100 2.400 2893.240 17.010 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 2240.750 1688.640 2241.030 1688.920 ;
        RECT 2245.810 1688.640 2246.090 1688.920 ;
      LAYER met3 ;
        RECT 2240.725 1688.930 2241.055 1688.945 ;
        RECT 2245.785 1688.930 2246.115 1688.945 ;
        RECT 2240.725 1688.630 2246.115 1688.930 ;
        RECT 2240.725 1688.615 2241.055 1688.630 ;
        RECT 2245.785 1688.615 2246.115 1688.630 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2652.890 19.620 2653.210 19.680 ;
        RECT 2910.950 19.620 2911.270 19.680 ;
        RECT 2652.890 19.480 2911.270 19.620 ;
        RECT 2652.890 19.420 2653.210 19.480 ;
        RECT 2910.950 19.420 2911.270 19.480 ;
      LAYER via ;
        RECT 2652.920 19.420 2653.180 19.680 ;
        RECT 2910.980 19.420 2911.240 19.680 ;
      LAYER met2 ;
        RECT 2247.585 1700.000 2247.865 1704.000 ;
        RECT 2247.720 1686.925 2247.860 1700.000 ;
        RECT 2247.650 1686.555 2247.930 1686.925 ;
        RECT 2652.910 1686.555 2653.190 1686.925 ;
        RECT 2652.980 19.710 2653.120 1686.555 ;
        RECT 2652.920 19.390 2653.180 19.710 ;
        RECT 2910.980 19.390 2911.240 19.710 ;
        RECT 2911.040 2.400 2911.180 19.390 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 2247.650 1686.600 2247.930 1686.880 ;
        RECT 2652.910 1686.600 2653.190 1686.880 ;
      LAYER met3 ;
        RECT 2247.625 1686.890 2247.955 1686.905 ;
        RECT 2652.885 1686.890 2653.215 1686.905 ;
        RECT 2247.625 1686.590 2653.215 1686.890 ;
        RECT 2247.625 1686.575 2247.955 1686.590 ;
        RECT 2652.885 1686.575 2653.215 1686.590 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 67.220 862.430 67.280 ;
        RECT 1471.150 67.220 1471.470 67.280 ;
        RECT 862.110 67.080 1471.470 67.220 ;
        RECT 862.110 67.020 862.430 67.080 ;
        RECT 1471.150 67.020 1471.470 67.080 ;
        RECT 858.890 2.960 859.210 3.020 ;
        RECT 862.110 2.960 862.430 3.020 ;
        RECT 858.890 2.820 862.430 2.960 ;
        RECT 858.890 2.760 859.210 2.820 ;
        RECT 862.110 2.760 862.430 2.820 ;
      LAYER via ;
        RECT 862.140 67.020 862.400 67.280 ;
        RECT 1471.180 67.020 1471.440 67.280 ;
        RECT 858.920 2.760 859.180 3.020 ;
        RECT 862.140 2.760 862.400 3.020 ;
      LAYER met2 ;
        RECT 1472.945 1700.410 1473.225 1704.000 ;
        RECT 1471.240 1700.270 1473.225 1700.410 ;
        RECT 1471.240 67.310 1471.380 1700.270 ;
        RECT 1472.945 1700.000 1473.225 1700.270 ;
        RECT 862.140 66.990 862.400 67.310 ;
        RECT 1471.180 66.990 1471.440 67.310 ;
        RECT 862.200 3.050 862.340 66.990 ;
        RECT 858.920 2.730 859.180 3.050 ;
        RECT 862.140 2.730 862.400 3.050 ;
        RECT 858.980 2.400 859.120 2.730 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 67.560 883.130 67.620 ;
        RECT 1478.050 67.560 1478.370 67.620 ;
        RECT 882.810 67.420 1478.370 67.560 ;
        RECT 882.810 67.360 883.130 67.420 ;
        RECT 1478.050 67.360 1478.370 67.420 ;
        RECT 876.830 34.580 877.150 34.640 ;
        RECT 882.810 34.580 883.130 34.640 ;
        RECT 876.830 34.440 883.130 34.580 ;
        RECT 876.830 34.380 877.150 34.440 ;
        RECT 882.810 34.380 883.130 34.440 ;
      LAYER via ;
        RECT 882.840 67.360 883.100 67.620 ;
        RECT 1478.080 67.360 1478.340 67.620 ;
        RECT 876.860 34.380 877.120 34.640 ;
        RECT 882.840 34.380 883.100 34.640 ;
      LAYER met2 ;
        RECT 1479.845 1700.410 1480.125 1704.000 ;
        RECT 1478.140 1700.270 1480.125 1700.410 ;
        RECT 1478.140 67.650 1478.280 1700.270 ;
        RECT 1479.845 1700.000 1480.125 1700.270 ;
        RECT 882.840 67.330 883.100 67.650 ;
        RECT 1478.080 67.330 1478.340 67.650 ;
        RECT 882.900 34.670 883.040 67.330 ;
        RECT 876.860 34.350 877.120 34.670 ;
        RECT 882.840 34.350 883.100 34.670 ;
        RECT 876.920 2.400 877.060 34.350 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 896.610 67.900 896.930 67.960 ;
        RECT 1484.950 67.900 1485.270 67.960 ;
        RECT 896.610 67.760 1485.270 67.900 ;
        RECT 896.610 67.700 896.930 67.760 ;
        RECT 1484.950 67.700 1485.270 67.760 ;
        RECT 894.770 2.960 895.090 3.020 ;
        RECT 896.610 2.960 896.930 3.020 ;
        RECT 894.770 2.820 896.930 2.960 ;
        RECT 894.770 2.760 895.090 2.820 ;
        RECT 896.610 2.760 896.930 2.820 ;
      LAYER via ;
        RECT 896.640 67.700 896.900 67.960 ;
        RECT 1484.980 67.700 1485.240 67.960 ;
        RECT 894.800 2.760 895.060 3.020 ;
        RECT 896.640 2.760 896.900 3.020 ;
      LAYER met2 ;
        RECT 1486.285 1700.410 1486.565 1704.000 ;
        RECT 1485.040 1700.270 1486.565 1700.410 ;
        RECT 1485.040 67.990 1485.180 1700.270 ;
        RECT 1486.285 1700.000 1486.565 1700.270 ;
        RECT 896.640 67.670 896.900 67.990 ;
        RECT 1484.980 67.670 1485.240 67.990 ;
        RECT 896.700 3.050 896.840 67.670 ;
        RECT 894.800 2.730 895.060 3.050 ;
        RECT 896.640 2.730 896.900 3.050 ;
        RECT 894.860 2.400 895.000 2.730 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 917.310 68.240 917.630 68.300 ;
        RECT 1491.390 68.240 1491.710 68.300 ;
        RECT 917.310 68.100 1491.710 68.240 ;
        RECT 917.310 68.040 917.630 68.100 ;
        RECT 1491.390 68.040 1491.710 68.100 ;
        RECT 912.710 2.960 913.030 3.020 ;
        RECT 917.310 2.960 917.630 3.020 ;
        RECT 912.710 2.820 917.630 2.960 ;
        RECT 912.710 2.760 913.030 2.820 ;
        RECT 917.310 2.760 917.630 2.820 ;
      LAYER via ;
        RECT 917.340 68.040 917.600 68.300 ;
        RECT 1491.420 68.040 1491.680 68.300 ;
        RECT 912.740 2.760 913.000 3.020 ;
        RECT 917.340 2.760 917.600 3.020 ;
      LAYER met2 ;
        RECT 1493.185 1700.410 1493.465 1704.000 ;
        RECT 1491.480 1700.270 1493.465 1700.410 ;
        RECT 1491.480 68.330 1491.620 1700.270 ;
        RECT 1493.185 1700.000 1493.465 1700.270 ;
        RECT 917.340 68.010 917.600 68.330 ;
        RECT 1491.420 68.010 1491.680 68.330 ;
        RECT 917.400 3.050 917.540 68.010 ;
        RECT 912.740 2.730 913.000 3.050 ;
        RECT 917.340 2.730 917.600 3.050 ;
        RECT 912.800 2.400 912.940 2.730 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 68.580 931.430 68.640 ;
        RECT 1498.290 68.580 1498.610 68.640 ;
        RECT 931.110 68.440 1498.610 68.580 ;
        RECT 931.110 68.380 931.430 68.440 ;
        RECT 1498.290 68.380 1498.610 68.440 ;
      LAYER via ;
        RECT 931.140 68.380 931.400 68.640 ;
        RECT 1498.320 68.380 1498.580 68.640 ;
      LAYER met2 ;
        RECT 1500.085 1700.410 1500.365 1704.000 ;
        RECT 1498.380 1700.270 1500.365 1700.410 ;
        RECT 1498.380 68.670 1498.520 1700.270 ;
        RECT 1500.085 1700.000 1500.365 1700.270 ;
        RECT 931.140 68.350 931.400 68.670 ;
        RECT 1498.320 68.350 1498.580 68.670 ;
        RECT 931.200 3.130 931.340 68.350 ;
        RECT 930.740 2.990 931.340 3.130 ;
        RECT 930.740 2.960 930.880 2.990 ;
        RECT 930.280 2.820 930.880 2.960 ;
        RECT 930.280 2.400 930.420 2.820 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 68.920 952.130 68.980 ;
        RECT 1505.190 68.920 1505.510 68.980 ;
        RECT 951.810 68.780 1505.510 68.920 ;
        RECT 951.810 68.720 952.130 68.780 ;
        RECT 1505.190 68.720 1505.510 68.780 ;
        RECT 948.130 2.960 948.450 3.020 ;
        RECT 951.810 2.960 952.130 3.020 ;
        RECT 948.130 2.820 952.130 2.960 ;
        RECT 948.130 2.760 948.450 2.820 ;
        RECT 951.810 2.760 952.130 2.820 ;
      LAYER via ;
        RECT 951.840 68.720 952.100 68.980 ;
        RECT 1505.220 68.720 1505.480 68.980 ;
        RECT 948.160 2.760 948.420 3.020 ;
        RECT 951.840 2.760 952.100 3.020 ;
      LAYER met2 ;
        RECT 1506.525 1700.410 1506.805 1704.000 ;
        RECT 1505.280 1700.270 1506.805 1700.410 ;
        RECT 1505.280 69.010 1505.420 1700.270 ;
        RECT 1506.525 1700.000 1506.805 1700.270 ;
        RECT 951.840 68.690 952.100 69.010 ;
        RECT 1505.220 68.690 1505.480 69.010 ;
        RECT 951.900 3.050 952.040 68.690 ;
        RECT 948.160 2.730 948.420 3.050 ;
        RECT 951.840 2.730 952.100 3.050 ;
        RECT 948.220 2.400 948.360 2.730 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 65.180 972.830 65.240 ;
        RECT 1512.090 65.180 1512.410 65.240 ;
        RECT 972.510 65.040 1512.410 65.180 ;
        RECT 972.510 64.980 972.830 65.040 ;
        RECT 1512.090 64.980 1512.410 65.040 ;
        RECT 966.070 34.580 966.390 34.640 ;
        RECT 972.510 34.580 972.830 34.640 ;
        RECT 966.070 34.440 972.830 34.580 ;
        RECT 966.070 34.380 966.390 34.440 ;
        RECT 972.510 34.380 972.830 34.440 ;
      LAYER via ;
        RECT 972.540 64.980 972.800 65.240 ;
        RECT 1512.120 64.980 1512.380 65.240 ;
        RECT 966.100 34.380 966.360 34.640 ;
        RECT 972.540 34.380 972.800 34.640 ;
      LAYER met2 ;
        RECT 1513.425 1700.410 1513.705 1704.000 ;
        RECT 1512.180 1700.270 1513.705 1700.410 ;
        RECT 1512.180 65.270 1512.320 1700.270 ;
        RECT 1513.425 1700.000 1513.705 1700.270 ;
        RECT 972.540 64.950 972.800 65.270 ;
        RECT 1512.120 64.950 1512.380 65.270 ;
        RECT 972.600 34.670 972.740 64.950 ;
        RECT 966.100 34.350 966.360 34.670 ;
        RECT 972.540 34.350 972.800 34.670 ;
        RECT 966.160 2.400 966.300 34.350 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 986.310 70.280 986.630 70.340 ;
        RECT 1519.450 70.280 1519.770 70.340 ;
        RECT 986.310 70.140 1519.770 70.280 ;
        RECT 986.310 70.080 986.630 70.140 ;
        RECT 1519.450 70.080 1519.770 70.140 ;
        RECT 984.010 2.960 984.330 3.020 ;
        RECT 986.310 2.960 986.630 3.020 ;
        RECT 984.010 2.820 986.630 2.960 ;
        RECT 984.010 2.760 984.330 2.820 ;
        RECT 986.310 2.760 986.630 2.820 ;
      LAYER via ;
        RECT 986.340 70.080 986.600 70.340 ;
        RECT 1519.480 70.080 1519.740 70.340 ;
        RECT 984.040 2.760 984.300 3.020 ;
        RECT 986.340 2.760 986.600 3.020 ;
      LAYER met2 ;
        RECT 1520.325 1700.410 1520.605 1704.000 ;
        RECT 1519.540 1700.270 1520.605 1700.410 ;
        RECT 1519.540 70.370 1519.680 1700.270 ;
        RECT 1520.325 1700.000 1520.605 1700.270 ;
        RECT 986.340 70.050 986.600 70.370 ;
        RECT 1519.480 70.050 1519.740 70.370 ;
        RECT 986.400 3.050 986.540 70.050 ;
        RECT 984.040 2.730 984.300 3.050 ;
        RECT 986.340 2.730 986.600 3.050 ;
        RECT 984.100 2.400 984.240 2.730 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1394.790 1678.140 1395.110 1678.200 ;
        RECT 1397.550 1678.140 1397.870 1678.200 ;
        RECT 1394.790 1678.000 1397.870 1678.140 ;
        RECT 1394.790 1677.940 1395.110 1678.000 ;
        RECT 1397.550 1677.940 1397.870 1678.000 ;
      LAYER via ;
        RECT 1394.820 1677.940 1395.080 1678.200 ;
        RECT 1397.580 1677.940 1397.840 1678.200 ;
      LAYER met2 ;
        RECT 1398.885 1700.410 1399.165 1704.000 ;
        RECT 1397.640 1700.270 1399.165 1700.410 ;
        RECT 1397.640 1678.230 1397.780 1700.270 ;
        RECT 1398.885 1700.000 1399.165 1700.270 ;
        RECT 1394.820 1677.910 1395.080 1678.230 ;
        RECT 1397.580 1677.910 1397.840 1678.230 ;
        RECT 1394.880 44.725 1395.020 1677.910 ;
        RECT 662.950 44.355 663.230 44.725 ;
        RECT 1394.810 44.355 1395.090 44.725 ;
        RECT 663.020 2.400 663.160 44.355 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 662.950 44.400 663.230 44.680 ;
        RECT 1394.810 44.400 1395.090 44.680 ;
      LAYER met3 ;
        RECT 662.925 44.690 663.255 44.705 ;
        RECT 1394.785 44.690 1395.115 44.705 ;
        RECT 662.925 44.390 1395.115 44.690 ;
        RECT 662.925 44.375 663.255 44.390 ;
        RECT 1394.785 44.375 1395.115 44.390 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1525.430 517.860 1525.750 518.120 ;
        RECT 1525.520 517.440 1525.660 517.860 ;
        RECT 1525.430 517.180 1525.750 517.440 ;
        RECT 1001.950 47.840 1002.270 47.900 ;
        RECT 1525.430 47.840 1525.750 47.900 ;
        RECT 1001.950 47.700 1525.750 47.840 ;
        RECT 1001.950 47.640 1002.270 47.700 ;
        RECT 1525.430 47.640 1525.750 47.700 ;
      LAYER via ;
        RECT 1525.460 517.860 1525.720 518.120 ;
        RECT 1525.460 517.180 1525.720 517.440 ;
        RECT 1001.980 47.640 1002.240 47.900 ;
        RECT 1525.460 47.640 1525.720 47.900 ;
      LAYER met2 ;
        RECT 1526.765 1700.410 1527.045 1704.000 ;
        RECT 1525.520 1700.270 1527.045 1700.410 ;
        RECT 1525.520 518.150 1525.660 1700.270 ;
        RECT 1526.765 1700.000 1527.045 1700.270 ;
        RECT 1525.460 517.830 1525.720 518.150 ;
        RECT 1525.460 517.150 1525.720 517.470 ;
        RECT 1525.520 47.930 1525.660 517.150 ;
        RECT 1001.980 47.610 1002.240 47.930 ;
        RECT 1525.460 47.610 1525.720 47.930 ;
        RECT 1002.040 2.400 1002.180 47.610 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1019.430 48.180 1019.750 48.240 ;
        RECT 1532.790 48.180 1533.110 48.240 ;
        RECT 1019.430 48.040 1533.110 48.180 ;
        RECT 1019.430 47.980 1019.750 48.040 ;
        RECT 1532.790 47.980 1533.110 48.040 ;
      LAYER via ;
        RECT 1019.460 47.980 1019.720 48.240 ;
        RECT 1532.820 47.980 1533.080 48.240 ;
      LAYER met2 ;
        RECT 1533.665 1700.410 1533.945 1704.000 ;
        RECT 1532.880 1700.270 1533.945 1700.410 ;
        RECT 1532.880 48.270 1533.020 1700.270 ;
        RECT 1533.665 1700.000 1533.945 1700.270 ;
        RECT 1019.460 47.950 1019.720 48.270 ;
        RECT 1532.820 47.950 1533.080 48.270 ;
        RECT 1019.520 2.400 1019.660 47.950 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 44.440 1037.690 44.500 ;
        RECT 1539.230 44.440 1539.550 44.500 ;
        RECT 1037.370 44.300 1539.550 44.440 ;
        RECT 1037.370 44.240 1037.690 44.300 ;
        RECT 1539.230 44.240 1539.550 44.300 ;
      LAYER via ;
        RECT 1037.400 44.240 1037.660 44.500 ;
        RECT 1539.260 44.240 1539.520 44.500 ;
      LAYER met2 ;
        RECT 1540.565 1700.410 1540.845 1704.000 ;
        RECT 1539.320 1700.270 1540.845 1700.410 ;
        RECT 1539.320 44.530 1539.460 1700.270 ;
        RECT 1540.565 1700.000 1540.845 1700.270 ;
        RECT 1037.400 44.210 1037.660 44.530 ;
        RECT 1539.260 44.210 1539.520 44.530 ;
        RECT 1037.460 2.400 1037.600 44.210 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1054.390 44.100 1054.710 44.160 ;
        RECT 1546.130 44.100 1546.450 44.160 ;
        RECT 1054.390 43.960 1546.450 44.100 ;
        RECT 1054.390 43.900 1054.710 43.960 ;
        RECT 1546.130 43.900 1546.450 43.960 ;
      LAYER via ;
        RECT 1054.420 43.900 1054.680 44.160 ;
        RECT 1546.160 43.900 1546.420 44.160 ;
      LAYER met2 ;
        RECT 1547.005 1700.410 1547.285 1704.000 ;
        RECT 1546.220 1700.270 1547.285 1700.410 ;
        RECT 1546.220 44.190 1546.360 1700.270 ;
        RECT 1547.005 1700.000 1547.285 1700.270 ;
        RECT 1054.420 43.870 1054.680 44.190 ;
        RECT 1546.160 43.870 1546.420 44.190 ;
        RECT 1054.480 28.970 1054.620 43.870 ;
        RECT 1054.480 28.830 1055.540 28.970 ;
        RECT 1055.400 2.400 1055.540 28.830 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1073.250 43.760 1073.570 43.820 ;
        RECT 1553.030 43.760 1553.350 43.820 ;
        RECT 1073.250 43.620 1553.350 43.760 ;
        RECT 1073.250 43.560 1073.570 43.620 ;
        RECT 1553.030 43.560 1553.350 43.620 ;
      LAYER via ;
        RECT 1073.280 43.560 1073.540 43.820 ;
        RECT 1553.060 43.560 1553.320 43.820 ;
      LAYER met2 ;
        RECT 1553.905 1700.410 1554.185 1704.000 ;
        RECT 1553.120 1700.270 1554.185 1700.410 ;
        RECT 1553.120 43.850 1553.260 1700.270 ;
        RECT 1553.905 1700.000 1554.185 1700.270 ;
        RECT 1073.280 43.530 1073.540 43.850 ;
        RECT 1553.060 43.530 1553.320 43.850 ;
        RECT 1073.340 2.400 1073.480 43.530 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.730 43.420 1091.050 43.480 ;
        RECT 1559.930 43.420 1560.250 43.480 ;
        RECT 1090.730 43.280 1560.250 43.420 ;
        RECT 1090.730 43.220 1091.050 43.280 ;
        RECT 1559.930 43.220 1560.250 43.280 ;
      LAYER via ;
        RECT 1090.760 43.220 1091.020 43.480 ;
        RECT 1559.960 43.220 1560.220 43.480 ;
      LAYER met2 ;
        RECT 1560.345 1700.410 1560.625 1704.000 ;
        RECT 1560.020 1700.270 1560.625 1700.410 ;
        RECT 1560.020 43.510 1560.160 1700.270 ;
        RECT 1560.345 1700.000 1560.625 1700.270 ;
        RECT 1090.760 43.190 1091.020 43.510 ;
        RECT 1559.960 43.190 1560.220 43.510 ;
        RECT 1090.820 2.400 1090.960 43.190 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1108.670 43.080 1108.990 43.140 ;
        RECT 1566.830 43.080 1567.150 43.140 ;
        RECT 1108.670 42.940 1567.150 43.080 ;
        RECT 1108.670 42.880 1108.990 42.940 ;
        RECT 1566.830 42.880 1567.150 42.940 ;
      LAYER via ;
        RECT 1108.700 42.880 1108.960 43.140 ;
        RECT 1566.860 42.880 1567.120 43.140 ;
      LAYER met2 ;
        RECT 1567.245 1700.000 1567.525 1704.000 ;
        RECT 1567.380 1690.210 1567.520 1700.000 ;
        RECT 1566.920 1690.070 1567.520 1690.210 ;
        RECT 1566.920 43.170 1567.060 1690.070 ;
        RECT 1108.700 42.850 1108.960 43.170 ;
        RECT 1566.860 42.850 1567.120 43.170 ;
        RECT 1108.760 2.400 1108.900 42.850 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.610 42.740 1126.930 42.800 ;
        RECT 1573.730 42.740 1574.050 42.800 ;
        RECT 1126.610 42.600 1574.050 42.740 ;
        RECT 1126.610 42.540 1126.930 42.600 ;
        RECT 1573.730 42.540 1574.050 42.600 ;
      LAYER via ;
        RECT 1126.640 42.540 1126.900 42.800 ;
        RECT 1573.760 42.540 1574.020 42.800 ;
      LAYER met2 ;
        RECT 1574.145 1700.410 1574.425 1704.000 ;
        RECT 1573.820 1700.270 1574.425 1700.410 ;
        RECT 1573.820 42.830 1573.960 1700.270 ;
        RECT 1574.145 1700.000 1574.425 1700.270 ;
        RECT 1126.640 42.510 1126.900 42.830 ;
        RECT 1573.760 42.510 1574.020 42.830 ;
        RECT 1126.700 2.400 1126.840 42.510 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1144.550 42.400 1144.870 42.460 ;
        RECT 1580.630 42.400 1580.950 42.460 ;
        RECT 1144.550 42.260 1580.950 42.400 ;
        RECT 1144.550 42.200 1144.870 42.260 ;
        RECT 1580.630 42.200 1580.950 42.260 ;
      LAYER via ;
        RECT 1144.580 42.200 1144.840 42.460 ;
        RECT 1580.660 42.200 1580.920 42.460 ;
      LAYER met2 ;
        RECT 1580.585 1700.000 1580.865 1704.000 ;
        RECT 1580.720 42.490 1580.860 1700.000 ;
        RECT 1144.580 42.170 1144.840 42.490 ;
        RECT 1580.660 42.170 1580.920 42.490 ;
        RECT 1144.640 2.400 1144.780 42.170 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 42.060 1162.810 42.120 ;
        RECT 1587.990 42.060 1588.310 42.120 ;
        RECT 1162.490 41.920 1588.310 42.060 ;
        RECT 1162.490 41.860 1162.810 41.920 ;
        RECT 1587.990 41.860 1588.310 41.920 ;
      LAYER via ;
        RECT 1162.520 41.860 1162.780 42.120 ;
        RECT 1588.020 41.860 1588.280 42.120 ;
      LAYER met2 ;
        RECT 1587.485 1700.000 1587.765 1704.000 ;
        RECT 1587.620 1666.410 1587.760 1700.000 ;
        RECT 1587.620 1666.270 1588.220 1666.410 ;
        RECT 1588.080 42.150 1588.220 1666.270 ;
        RECT 1162.520 41.830 1162.780 42.150 ;
        RECT 1588.020 41.830 1588.280 42.150 ;
        RECT 1162.580 2.400 1162.720 41.830 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1402.685 476.085 1402.855 524.195 ;
        RECT 1402.685 144.245 1402.855 222.615 ;
      LAYER mcon ;
        RECT 1402.685 524.025 1402.855 524.195 ;
        RECT 1402.685 222.445 1402.855 222.615 ;
      LAYER met1 ;
        RECT 1402.610 1594.160 1402.930 1594.220 ;
        RECT 1403.070 1594.160 1403.390 1594.220 ;
        RECT 1402.610 1594.020 1403.390 1594.160 ;
        RECT 1402.610 1593.960 1402.930 1594.020 ;
        RECT 1403.070 1593.960 1403.390 1594.020 ;
        RECT 1402.150 1511.200 1402.470 1511.260 ;
        RECT 1403.070 1511.200 1403.390 1511.260 ;
        RECT 1402.150 1511.060 1403.390 1511.200 ;
        RECT 1402.150 1511.000 1402.470 1511.060 ;
        RECT 1403.070 1511.000 1403.390 1511.060 ;
        RECT 1402.150 1414.640 1402.470 1414.700 ;
        RECT 1403.070 1414.640 1403.390 1414.700 ;
        RECT 1402.150 1414.500 1403.390 1414.640 ;
        RECT 1402.150 1414.440 1402.470 1414.500 ;
        RECT 1403.070 1414.440 1403.390 1414.500 ;
        RECT 1402.150 1318.080 1402.470 1318.140 ;
        RECT 1403.070 1318.080 1403.390 1318.140 ;
        RECT 1402.150 1317.940 1403.390 1318.080 ;
        RECT 1402.150 1317.880 1402.470 1317.940 ;
        RECT 1403.070 1317.880 1403.390 1317.940 ;
        RECT 1403.070 1173.580 1403.390 1173.640 ;
        RECT 1402.700 1173.440 1403.390 1173.580 ;
        RECT 1402.700 1172.960 1402.840 1173.440 ;
        RECT 1403.070 1173.380 1403.390 1173.440 ;
        RECT 1402.610 1172.700 1402.930 1172.960 ;
        RECT 1402.150 931.500 1402.470 931.560 ;
        RECT 1403.070 931.500 1403.390 931.560 ;
        RECT 1402.150 931.360 1403.390 931.500 ;
        RECT 1402.150 931.300 1402.470 931.360 ;
        RECT 1403.070 931.300 1403.390 931.360 ;
        RECT 1402.610 786.800 1402.930 787.060 ;
        RECT 1402.700 786.320 1402.840 786.800 ;
        RECT 1403.070 786.320 1403.390 786.380 ;
        RECT 1402.700 786.180 1403.390 786.320 ;
        RECT 1403.070 786.120 1403.390 786.180 ;
        RECT 1402.150 738.380 1402.470 738.440 ;
        RECT 1403.070 738.380 1403.390 738.440 ;
        RECT 1402.150 738.240 1403.390 738.380 ;
        RECT 1402.150 738.180 1402.470 738.240 ;
        RECT 1403.070 738.180 1403.390 738.240 ;
        RECT 1402.610 593.340 1402.930 593.600 ;
        RECT 1402.700 593.200 1402.840 593.340 ;
        RECT 1403.070 593.200 1403.390 593.260 ;
        RECT 1402.700 593.060 1403.390 593.200 ;
        RECT 1403.070 593.000 1403.390 593.060 ;
        RECT 1402.150 545.260 1402.470 545.320 ;
        RECT 1403.070 545.260 1403.390 545.320 ;
        RECT 1402.150 545.120 1403.390 545.260 ;
        RECT 1402.150 545.060 1402.470 545.120 ;
        RECT 1403.070 545.060 1403.390 545.120 ;
        RECT 1402.610 524.180 1402.930 524.240 ;
        RECT 1402.415 524.040 1402.930 524.180 ;
        RECT 1402.610 523.980 1402.930 524.040 ;
        RECT 1402.625 476.240 1402.915 476.285 ;
        RECT 1403.070 476.240 1403.390 476.300 ;
        RECT 1402.625 476.100 1403.390 476.240 ;
        RECT 1402.625 476.055 1402.915 476.100 ;
        RECT 1403.070 476.040 1403.390 476.100 ;
        RECT 1402.150 448.700 1402.470 448.760 ;
        RECT 1403.070 448.700 1403.390 448.760 ;
        RECT 1402.150 448.560 1403.390 448.700 ;
        RECT 1402.150 448.500 1402.470 448.560 ;
        RECT 1403.070 448.500 1403.390 448.560 ;
        RECT 1402.610 366.080 1402.930 366.140 ;
        RECT 1403.070 366.080 1403.390 366.140 ;
        RECT 1402.610 365.940 1403.390 366.080 ;
        RECT 1402.610 365.880 1402.930 365.940 ;
        RECT 1403.070 365.880 1403.390 365.940 ;
        RECT 1401.230 317.460 1401.550 317.520 ;
        RECT 1402.610 317.460 1402.930 317.520 ;
        RECT 1401.230 317.320 1402.930 317.460 ;
        RECT 1401.230 317.260 1401.550 317.320 ;
        RECT 1402.610 317.260 1402.930 317.320 ;
        RECT 1401.230 222.600 1401.550 222.660 ;
        RECT 1402.625 222.600 1402.915 222.645 ;
        RECT 1401.230 222.460 1402.915 222.600 ;
        RECT 1401.230 222.400 1401.550 222.460 ;
        RECT 1402.625 222.415 1402.915 222.460 ;
        RECT 1402.610 144.400 1402.930 144.460 ;
        RECT 1402.415 144.260 1402.930 144.400 ;
        RECT 1402.610 144.200 1402.930 144.260 ;
        RECT 1402.150 90.000 1402.470 90.060 ;
        RECT 1402.610 90.000 1402.930 90.060 ;
        RECT 1402.150 89.860 1402.930 90.000 ;
        RECT 1402.150 89.800 1402.470 89.860 ;
        RECT 1402.610 89.800 1402.930 89.860 ;
        RECT 680.410 46.140 680.730 46.200 ;
        RECT 1402.150 46.140 1402.470 46.200 ;
        RECT 680.410 46.000 1402.470 46.140 ;
        RECT 680.410 45.940 680.730 46.000 ;
        RECT 1402.150 45.940 1402.470 46.000 ;
      LAYER via ;
        RECT 1402.640 1593.960 1402.900 1594.220 ;
        RECT 1403.100 1593.960 1403.360 1594.220 ;
        RECT 1402.180 1511.000 1402.440 1511.260 ;
        RECT 1403.100 1511.000 1403.360 1511.260 ;
        RECT 1402.180 1414.440 1402.440 1414.700 ;
        RECT 1403.100 1414.440 1403.360 1414.700 ;
        RECT 1402.180 1317.880 1402.440 1318.140 ;
        RECT 1403.100 1317.880 1403.360 1318.140 ;
        RECT 1403.100 1173.380 1403.360 1173.640 ;
        RECT 1402.640 1172.700 1402.900 1172.960 ;
        RECT 1402.180 931.300 1402.440 931.560 ;
        RECT 1403.100 931.300 1403.360 931.560 ;
        RECT 1402.640 786.800 1402.900 787.060 ;
        RECT 1403.100 786.120 1403.360 786.380 ;
        RECT 1402.180 738.180 1402.440 738.440 ;
        RECT 1403.100 738.180 1403.360 738.440 ;
        RECT 1402.640 593.340 1402.900 593.600 ;
        RECT 1403.100 593.000 1403.360 593.260 ;
        RECT 1402.180 545.060 1402.440 545.320 ;
        RECT 1403.100 545.060 1403.360 545.320 ;
        RECT 1402.640 523.980 1402.900 524.240 ;
        RECT 1403.100 476.040 1403.360 476.300 ;
        RECT 1402.180 448.500 1402.440 448.760 ;
        RECT 1403.100 448.500 1403.360 448.760 ;
        RECT 1402.640 365.880 1402.900 366.140 ;
        RECT 1403.100 365.880 1403.360 366.140 ;
        RECT 1401.260 317.260 1401.520 317.520 ;
        RECT 1402.640 317.260 1402.900 317.520 ;
        RECT 1401.260 222.400 1401.520 222.660 ;
        RECT 1402.640 144.200 1402.900 144.460 ;
        RECT 1402.180 89.800 1402.440 90.060 ;
        RECT 1402.640 89.800 1402.900 90.060 ;
        RECT 680.440 45.940 680.700 46.200 ;
        RECT 1402.180 45.940 1402.440 46.200 ;
      LAYER met2 ;
        RECT 1405.785 1700.410 1406.065 1704.000 ;
        RECT 1404.540 1700.270 1406.065 1700.410 ;
        RECT 1404.540 1656.210 1404.680 1700.270 ;
        RECT 1405.785 1700.000 1406.065 1700.270 ;
        RECT 1403.160 1656.070 1404.680 1656.210 ;
        RECT 1403.160 1594.250 1403.300 1656.070 ;
        RECT 1402.640 1593.930 1402.900 1594.250 ;
        RECT 1403.100 1593.930 1403.360 1594.250 ;
        RECT 1402.700 1559.650 1402.840 1593.930 ;
        RECT 1402.700 1559.510 1403.300 1559.650 ;
        RECT 1403.160 1511.290 1403.300 1559.510 ;
        RECT 1402.180 1510.970 1402.440 1511.290 ;
        RECT 1403.100 1510.970 1403.360 1511.290 ;
        RECT 1402.240 1510.690 1402.380 1510.970 ;
        RECT 1402.240 1510.550 1402.840 1510.690 ;
        RECT 1402.700 1463.090 1402.840 1510.550 ;
        RECT 1402.700 1462.950 1403.300 1463.090 ;
        RECT 1403.160 1414.730 1403.300 1462.950 ;
        RECT 1402.180 1414.410 1402.440 1414.730 ;
        RECT 1403.100 1414.410 1403.360 1414.730 ;
        RECT 1402.240 1414.130 1402.380 1414.410 ;
        RECT 1402.240 1413.990 1402.840 1414.130 ;
        RECT 1402.700 1366.530 1402.840 1413.990 ;
        RECT 1402.700 1366.390 1403.300 1366.530 ;
        RECT 1403.160 1318.170 1403.300 1366.390 ;
        RECT 1402.180 1317.850 1402.440 1318.170 ;
        RECT 1403.100 1317.850 1403.360 1318.170 ;
        RECT 1402.240 1317.570 1402.380 1317.850 ;
        RECT 1402.240 1317.430 1402.840 1317.570 ;
        RECT 1402.700 1269.970 1402.840 1317.430 ;
        RECT 1402.700 1269.830 1403.300 1269.970 ;
        RECT 1403.160 1173.670 1403.300 1269.830 ;
        RECT 1403.100 1173.350 1403.360 1173.670 ;
        RECT 1402.640 1172.670 1402.900 1172.990 ;
        RECT 1402.700 1125.130 1402.840 1172.670 ;
        RECT 1402.240 1124.990 1402.840 1125.130 ;
        RECT 1402.240 1124.450 1402.380 1124.990 ;
        RECT 1402.240 1124.310 1402.840 1124.450 ;
        RECT 1402.700 1028.570 1402.840 1124.310 ;
        RECT 1402.240 1028.430 1402.840 1028.570 ;
        RECT 1402.240 1027.890 1402.380 1028.430 ;
        RECT 1402.240 1027.750 1402.840 1027.890 ;
        RECT 1402.700 932.010 1402.840 1027.750 ;
        RECT 1402.240 931.870 1402.840 932.010 ;
        RECT 1402.240 931.590 1402.380 931.870 ;
        RECT 1402.180 931.270 1402.440 931.590 ;
        RECT 1403.100 931.270 1403.360 931.590 ;
        RECT 1403.160 883.730 1403.300 931.270 ;
        RECT 1403.160 883.590 1403.760 883.730 ;
        RECT 1403.620 883.050 1403.760 883.590 ;
        RECT 1402.700 882.910 1403.760 883.050 ;
        RECT 1402.700 835.450 1402.840 882.910 ;
        RECT 1402.240 835.310 1402.840 835.450 ;
        RECT 1402.240 834.770 1402.380 835.310 ;
        RECT 1402.240 834.630 1402.840 834.770 ;
        RECT 1402.700 787.090 1402.840 834.630 ;
        RECT 1402.640 786.770 1402.900 787.090 ;
        RECT 1403.100 786.090 1403.360 786.410 ;
        RECT 1403.160 738.470 1403.300 786.090 ;
        RECT 1402.180 738.210 1402.440 738.470 ;
        RECT 1402.180 738.150 1402.840 738.210 ;
        RECT 1403.100 738.150 1403.360 738.470 ;
        RECT 1402.240 738.070 1402.840 738.150 ;
        RECT 1402.700 642.330 1402.840 738.070 ;
        RECT 1402.240 642.190 1402.840 642.330 ;
        RECT 1402.240 641.650 1402.380 642.190 ;
        RECT 1402.240 641.510 1402.840 641.650 ;
        RECT 1402.700 593.630 1402.840 641.510 ;
        RECT 1402.640 593.310 1402.900 593.630 ;
        RECT 1403.100 592.970 1403.360 593.290 ;
        RECT 1403.160 545.350 1403.300 592.970 ;
        RECT 1402.180 545.090 1402.440 545.350 ;
        RECT 1402.180 545.030 1402.840 545.090 ;
        RECT 1403.100 545.030 1403.360 545.350 ;
        RECT 1402.240 544.950 1402.840 545.030 ;
        RECT 1402.700 524.270 1402.840 544.950 ;
        RECT 1402.640 523.950 1402.900 524.270 ;
        RECT 1403.100 476.010 1403.360 476.330 ;
        RECT 1403.160 448.790 1403.300 476.010 ;
        RECT 1402.180 448.530 1402.440 448.790 ;
        RECT 1403.100 448.530 1403.360 448.790 ;
        RECT 1402.180 448.470 1403.360 448.530 ;
        RECT 1402.240 448.390 1403.300 448.470 ;
        RECT 1403.160 366.170 1403.300 448.390 ;
        RECT 1402.640 365.850 1402.900 366.170 ;
        RECT 1403.100 365.850 1403.360 366.170 ;
        RECT 1402.700 317.550 1402.840 365.850 ;
        RECT 1401.260 317.230 1401.520 317.550 ;
        RECT 1402.640 317.230 1402.900 317.550 ;
        RECT 1401.320 222.690 1401.460 317.230 ;
        RECT 1401.260 222.370 1401.520 222.690 ;
        RECT 1402.640 144.170 1402.900 144.490 ;
        RECT 1402.700 90.090 1402.840 144.170 ;
        RECT 1402.180 89.770 1402.440 90.090 ;
        RECT 1402.640 89.770 1402.900 90.090 ;
        RECT 1402.240 46.230 1402.380 89.770 ;
        RECT 680.440 45.910 680.700 46.230 ;
        RECT 1402.180 45.910 1402.440 46.230 ;
        RECT 680.500 2.400 680.640 45.910 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 44.780 1180.290 44.840 ;
        RECT 1594.890 44.780 1595.210 44.840 ;
        RECT 1179.970 44.640 1595.210 44.780 ;
        RECT 1179.970 44.580 1180.290 44.640 ;
        RECT 1594.890 44.580 1595.210 44.640 ;
      LAYER via ;
        RECT 1180.000 44.580 1180.260 44.840 ;
        RECT 1594.920 44.580 1595.180 44.840 ;
      LAYER met2 ;
        RECT 1594.385 1700.410 1594.665 1704.000 ;
        RECT 1594.385 1700.270 1595.120 1700.410 ;
        RECT 1594.385 1700.000 1594.665 1700.270 ;
        RECT 1594.980 44.870 1595.120 1700.270 ;
        RECT 1180.000 44.550 1180.260 44.870 ;
        RECT 1594.920 44.550 1595.180 44.870 ;
        RECT 1180.060 2.400 1180.200 44.550 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1197.910 45.120 1198.230 45.180 ;
        RECT 1601.790 45.120 1602.110 45.180 ;
        RECT 1197.910 44.980 1602.110 45.120 ;
        RECT 1197.910 44.920 1198.230 44.980 ;
        RECT 1601.790 44.920 1602.110 44.980 ;
      LAYER via ;
        RECT 1197.940 44.920 1198.200 45.180 ;
        RECT 1601.820 44.920 1602.080 45.180 ;
      LAYER met2 ;
        RECT 1600.825 1700.410 1601.105 1704.000 ;
        RECT 1600.825 1700.270 1602.020 1700.410 ;
        RECT 1600.825 1700.000 1601.105 1700.270 ;
        RECT 1601.880 45.210 1602.020 1700.270 ;
        RECT 1197.940 44.890 1198.200 45.210 ;
        RECT 1601.820 44.890 1602.080 45.210 ;
        RECT 1198.000 2.400 1198.140 44.890 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1215.850 41.720 1216.170 41.780 ;
        RECT 1608.690 41.720 1609.010 41.780 ;
        RECT 1215.850 41.580 1609.010 41.720 ;
        RECT 1215.850 41.520 1216.170 41.580 ;
        RECT 1608.690 41.520 1609.010 41.580 ;
      LAYER via ;
        RECT 1215.880 41.520 1216.140 41.780 ;
        RECT 1608.720 41.520 1608.980 41.780 ;
      LAYER met2 ;
        RECT 1607.725 1700.410 1608.005 1704.000 ;
        RECT 1607.725 1700.270 1608.920 1700.410 ;
        RECT 1607.725 1700.000 1608.005 1700.270 ;
        RECT 1608.780 41.810 1608.920 1700.270 ;
        RECT 1215.880 41.490 1216.140 41.810 ;
        RECT 1608.720 41.490 1608.980 41.810 ;
        RECT 1215.940 2.400 1216.080 41.490 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 45.460 1234.110 45.520 ;
        RECT 1615.590 45.460 1615.910 45.520 ;
        RECT 1233.790 45.320 1615.910 45.460 ;
        RECT 1233.790 45.260 1234.110 45.320 ;
        RECT 1615.590 45.260 1615.910 45.320 ;
      LAYER via ;
        RECT 1233.820 45.260 1234.080 45.520 ;
        RECT 1615.620 45.260 1615.880 45.520 ;
      LAYER met2 ;
        RECT 1614.625 1700.410 1614.905 1704.000 ;
        RECT 1614.625 1700.270 1615.820 1700.410 ;
        RECT 1614.625 1700.000 1614.905 1700.270 ;
        RECT 1615.680 45.550 1615.820 1700.270 ;
        RECT 1233.820 45.230 1234.080 45.550 ;
        RECT 1615.620 45.230 1615.880 45.550 ;
        RECT 1233.880 2.400 1234.020 45.230 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1616.050 1678.140 1616.370 1678.200 ;
        RECT 1619.270 1678.140 1619.590 1678.200 ;
        RECT 1616.050 1678.000 1619.590 1678.140 ;
        RECT 1616.050 1677.940 1616.370 1678.000 ;
        RECT 1619.270 1677.940 1619.590 1678.000 ;
        RECT 1251.730 45.800 1252.050 45.860 ;
        RECT 1616.050 45.800 1616.370 45.860 ;
        RECT 1251.730 45.660 1616.370 45.800 ;
        RECT 1251.730 45.600 1252.050 45.660 ;
        RECT 1616.050 45.600 1616.370 45.660 ;
      LAYER via ;
        RECT 1616.080 1677.940 1616.340 1678.200 ;
        RECT 1619.300 1677.940 1619.560 1678.200 ;
        RECT 1251.760 45.600 1252.020 45.860 ;
        RECT 1616.080 45.600 1616.340 45.860 ;
      LAYER met2 ;
        RECT 1621.065 1700.410 1621.345 1704.000 ;
        RECT 1619.360 1700.270 1621.345 1700.410 ;
        RECT 1619.360 1678.230 1619.500 1700.270 ;
        RECT 1621.065 1700.000 1621.345 1700.270 ;
        RECT 1616.080 1677.910 1616.340 1678.230 ;
        RECT 1619.300 1677.910 1619.560 1678.230 ;
        RECT 1616.140 45.890 1616.280 1677.910 ;
        RECT 1251.760 45.570 1252.020 45.890 ;
        RECT 1616.080 45.570 1616.340 45.890 ;
        RECT 1251.820 2.400 1251.960 45.570 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1622.030 1675.080 1622.350 1675.140 ;
        RECT 1626.630 1675.080 1626.950 1675.140 ;
        RECT 1622.030 1674.940 1626.950 1675.080 ;
        RECT 1622.030 1674.880 1622.350 1674.940 ;
        RECT 1626.630 1674.880 1626.950 1674.940 ;
        RECT 1269.210 30.840 1269.530 30.900 ;
        RECT 1622.030 30.840 1622.350 30.900 ;
        RECT 1269.210 30.700 1622.350 30.840 ;
        RECT 1269.210 30.640 1269.530 30.700 ;
        RECT 1622.030 30.640 1622.350 30.700 ;
      LAYER via ;
        RECT 1622.060 1674.880 1622.320 1675.140 ;
        RECT 1626.660 1674.880 1626.920 1675.140 ;
        RECT 1269.240 30.640 1269.500 30.900 ;
        RECT 1622.060 30.640 1622.320 30.900 ;
      LAYER met2 ;
        RECT 1627.965 1700.410 1628.245 1704.000 ;
        RECT 1626.720 1700.270 1628.245 1700.410 ;
        RECT 1626.720 1675.170 1626.860 1700.270 ;
        RECT 1627.965 1700.000 1628.245 1700.270 ;
        RECT 1622.060 1674.850 1622.320 1675.170 ;
        RECT 1626.660 1674.850 1626.920 1675.170 ;
        RECT 1622.120 30.930 1622.260 1674.850 ;
        RECT 1269.240 30.610 1269.500 30.930 ;
        RECT 1622.060 30.610 1622.320 30.930 ;
        RECT 1269.300 2.400 1269.440 30.610 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1628.930 1678.140 1629.250 1678.200 ;
        RECT 1633.070 1678.140 1633.390 1678.200 ;
        RECT 1628.930 1678.000 1633.390 1678.140 ;
        RECT 1628.930 1677.940 1629.250 1678.000 ;
        RECT 1633.070 1677.940 1633.390 1678.000 ;
        RECT 1287.150 31.180 1287.470 31.240 ;
        RECT 1628.930 31.180 1629.250 31.240 ;
        RECT 1287.150 31.040 1629.250 31.180 ;
        RECT 1287.150 30.980 1287.470 31.040 ;
        RECT 1628.930 30.980 1629.250 31.040 ;
      LAYER via ;
        RECT 1628.960 1677.940 1629.220 1678.200 ;
        RECT 1633.100 1677.940 1633.360 1678.200 ;
        RECT 1287.180 30.980 1287.440 31.240 ;
        RECT 1628.960 30.980 1629.220 31.240 ;
      LAYER met2 ;
        RECT 1634.405 1700.410 1634.685 1704.000 ;
        RECT 1633.160 1700.270 1634.685 1700.410 ;
        RECT 1633.160 1678.230 1633.300 1700.270 ;
        RECT 1634.405 1700.000 1634.685 1700.270 ;
        RECT 1628.960 1677.910 1629.220 1678.230 ;
        RECT 1633.100 1677.910 1633.360 1678.230 ;
        RECT 1629.020 31.270 1629.160 1677.910 ;
        RECT 1287.180 30.950 1287.440 31.270 ;
        RECT 1628.960 30.950 1629.220 31.270 ;
        RECT 1287.240 2.400 1287.380 30.950 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1635.830 1678.140 1636.150 1678.200 ;
        RECT 1639.510 1678.140 1639.830 1678.200 ;
        RECT 1635.830 1678.000 1639.830 1678.140 ;
        RECT 1635.830 1677.940 1636.150 1678.000 ;
        RECT 1639.510 1677.940 1639.830 1678.000 ;
        RECT 1305.090 31.520 1305.410 31.580 ;
        RECT 1635.830 31.520 1636.150 31.580 ;
        RECT 1305.090 31.380 1636.150 31.520 ;
        RECT 1305.090 31.320 1305.410 31.380 ;
        RECT 1635.830 31.320 1636.150 31.380 ;
      LAYER via ;
        RECT 1635.860 1677.940 1636.120 1678.200 ;
        RECT 1639.540 1677.940 1639.800 1678.200 ;
        RECT 1305.120 31.320 1305.380 31.580 ;
        RECT 1635.860 31.320 1636.120 31.580 ;
      LAYER met2 ;
        RECT 1641.305 1700.410 1641.585 1704.000 ;
        RECT 1639.600 1700.270 1641.585 1700.410 ;
        RECT 1639.600 1678.230 1639.740 1700.270 ;
        RECT 1641.305 1700.000 1641.585 1700.270 ;
        RECT 1635.860 1677.910 1636.120 1678.230 ;
        RECT 1639.540 1677.910 1639.800 1678.230 ;
        RECT 1635.920 31.610 1636.060 1677.910 ;
        RECT 1305.120 31.290 1305.380 31.610 ;
        RECT 1635.860 31.290 1636.120 31.610 ;
        RECT 1305.180 2.400 1305.320 31.290 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1383.750 1688.680 1384.070 1688.740 ;
        RECT 1648.250 1688.680 1648.570 1688.740 ;
        RECT 1383.750 1688.540 1648.570 1688.680 ;
        RECT 1383.750 1688.480 1384.070 1688.540 ;
        RECT 1648.250 1688.480 1648.570 1688.540 ;
        RECT 1323.030 18.600 1323.350 18.660 ;
        RECT 1381.910 18.600 1382.230 18.660 ;
        RECT 1323.030 18.460 1382.230 18.600 ;
        RECT 1323.030 18.400 1323.350 18.460 ;
        RECT 1381.910 18.400 1382.230 18.460 ;
      LAYER via ;
        RECT 1383.780 1688.480 1384.040 1688.740 ;
        RECT 1648.280 1688.480 1648.540 1688.740 ;
        RECT 1323.060 18.400 1323.320 18.660 ;
        RECT 1381.940 18.400 1382.200 18.660 ;
      LAYER met2 ;
        RECT 1648.205 1700.000 1648.485 1704.000 ;
        RECT 1648.340 1688.770 1648.480 1700.000 ;
        RECT 1383.780 1688.450 1384.040 1688.770 ;
        RECT 1648.280 1688.450 1648.540 1688.770 ;
        RECT 1383.840 19.450 1383.980 1688.450 ;
        RECT 1382.000 19.310 1383.980 19.450 ;
        RECT 1382.000 18.690 1382.140 19.310 ;
        RECT 1323.060 18.370 1323.320 18.690 ;
        RECT 1381.940 18.370 1382.200 18.690 ;
        RECT 1323.120 2.400 1323.260 18.370 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1630.845 1686.655 1631.015 1686.995 ;
        RECT 1632.225 1686.655 1632.395 1688.015 ;
        RECT 1630.845 1686.485 1632.395 1686.655 ;
      LAYER mcon ;
        RECT 1632.225 1687.845 1632.395 1688.015 ;
        RECT 1630.845 1686.825 1631.015 1686.995 ;
      LAYER met1 ;
        RECT 1632.165 1688.000 1632.455 1688.045 ;
        RECT 1651.930 1688.000 1652.250 1688.060 ;
        RECT 1632.165 1687.860 1652.250 1688.000 ;
        RECT 1632.165 1687.815 1632.455 1687.860 ;
        RECT 1651.930 1687.800 1652.250 1687.860 ;
        RECT 1345.110 1686.980 1345.430 1687.040 ;
        RECT 1630.785 1686.980 1631.075 1687.025 ;
        RECT 1345.110 1686.840 1631.075 1686.980 ;
        RECT 1345.110 1686.780 1345.430 1686.840 ;
        RECT 1630.785 1686.795 1631.075 1686.840 ;
        RECT 1340.510 20.640 1340.830 20.700 ;
        RECT 1345.110 20.640 1345.430 20.700 ;
        RECT 1340.510 20.500 1345.430 20.640 ;
        RECT 1340.510 20.440 1340.830 20.500 ;
        RECT 1345.110 20.440 1345.430 20.500 ;
      LAYER via ;
        RECT 1651.960 1687.800 1652.220 1688.060 ;
        RECT 1345.140 1686.780 1345.400 1687.040 ;
        RECT 1340.540 20.440 1340.800 20.700 ;
        RECT 1345.140 20.440 1345.400 20.700 ;
      LAYER met2 ;
        RECT 1654.645 1700.410 1654.925 1704.000 ;
        RECT 1653.400 1700.270 1654.925 1700.410 ;
        RECT 1653.400 1688.850 1653.540 1700.270 ;
        RECT 1654.645 1700.000 1654.925 1700.270 ;
        RECT 1652.020 1688.710 1653.540 1688.850 ;
        RECT 1652.020 1688.090 1652.160 1688.710 ;
        RECT 1651.960 1687.770 1652.220 1688.090 ;
        RECT 1345.140 1686.750 1345.400 1687.070 ;
        RECT 1345.200 20.730 1345.340 1686.750 ;
        RECT 1340.540 20.410 1340.800 20.730 ;
        RECT 1345.140 20.410 1345.400 20.730 ;
        RECT 1340.600 2.400 1340.740 20.410 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1408.590 1678.140 1408.910 1678.200 ;
        RECT 1410.890 1678.140 1411.210 1678.200 ;
        RECT 1408.590 1678.000 1411.210 1678.140 ;
        RECT 1408.590 1677.940 1408.910 1678.000 ;
        RECT 1410.890 1677.940 1411.210 1678.000 ;
        RECT 698.350 46.480 698.670 46.540 ;
        RECT 1408.590 46.480 1408.910 46.540 ;
        RECT 698.350 46.340 1408.910 46.480 ;
        RECT 698.350 46.280 698.670 46.340 ;
        RECT 1408.590 46.280 1408.910 46.340 ;
      LAYER via ;
        RECT 1408.620 1677.940 1408.880 1678.200 ;
        RECT 1410.920 1677.940 1411.180 1678.200 ;
        RECT 698.380 46.280 698.640 46.540 ;
        RECT 1408.620 46.280 1408.880 46.540 ;
      LAYER met2 ;
        RECT 1412.225 1700.410 1412.505 1704.000 ;
        RECT 1410.980 1700.270 1412.505 1700.410 ;
        RECT 1410.980 1678.230 1411.120 1700.270 ;
        RECT 1412.225 1700.000 1412.505 1700.270 ;
        RECT 1408.620 1677.910 1408.880 1678.230 ;
        RECT 1410.920 1677.910 1411.180 1678.230 ;
        RECT 1408.680 46.570 1408.820 1677.910 ;
        RECT 698.380 46.250 698.640 46.570 ;
        RECT 1408.620 46.250 1408.880 46.570 ;
        RECT 698.440 2.400 698.580 46.250 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.450 14.860 1358.770 14.920 ;
        RECT 1369.490 14.860 1369.810 14.920 ;
        RECT 1358.450 14.720 1369.810 14.860 ;
        RECT 1358.450 14.660 1358.770 14.720 ;
        RECT 1369.490 14.660 1369.810 14.720 ;
      LAYER via ;
        RECT 1358.480 14.660 1358.740 14.920 ;
        RECT 1369.520 14.660 1369.780 14.920 ;
      LAYER met2 ;
        RECT 1661.545 1700.000 1661.825 1704.000 ;
        RECT 1661.680 1686.925 1661.820 1700.000 ;
        RECT 1369.510 1686.555 1369.790 1686.925 ;
        RECT 1661.610 1686.555 1661.890 1686.925 ;
        RECT 1369.580 14.950 1369.720 1686.555 ;
        RECT 1358.480 14.630 1358.740 14.950 ;
        RECT 1369.520 14.630 1369.780 14.950 ;
        RECT 1358.540 2.400 1358.680 14.630 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
      LAYER via2 ;
        RECT 1369.510 1686.600 1369.790 1686.880 ;
        RECT 1661.610 1686.600 1661.890 1686.880 ;
      LAYER met3 ;
        RECT 1369.485 1686.890 1369.815 1686.905 ;
        RECT 1661.585 1686.890 1661.915 1686.905 ;
        RECT 1369.485 1686.590 1661.915 1686.890 ;
        RECT 1369.485 1686.575 1369.815 1686.590 ;
        RECT 1661.585 1686.575 1661.915 1686.590 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.490 1688.340 1668.810 1688.400 ;
        RECT 1631.780 1688.200 1668.810 1688.340 ;
        RECT 1383.290 1688.000 1383.610 1688.060 ;
        RECT 1631.780 1688.000 1631.920 1688.200 ;
        RECT 1668.490 1688.140 1668.810 1688.200 ;
        RECT 1383.290 1687.860 1631.920 1688.000 ;
        RECT 1383.290 1687.800 1383.610 1687.860 ;
        RECT 1376.390 20.640 1376.710 20.700 ;
        RECT 1383.290 20.640 1383.610 20.700 ;
        RECT 1376.390 20.500 1383.610 20.640 ;
        RECT 1376.390 20.440 1376.710 20.500 ;
        RECT 1383.290 20.440 1383.610 20.500 ;
      LAYER via ;
        RECT 1383.320 1687.800 1383.580 1688.060 ;
        RECT 1668.520 1688.140 1668.780 1688.400 ;
        RECT 1376.420 20.440 1376.680 20.700 ;
        RECT 1383.320 20.440 1383.580 20.700 ;
      LAYER met2 ;
        RECT 1668.445 1700.000 1668.725 1704.000 ;
        RECT 1668.580 1688.430 1668.720 1700.000 ;
        RECT 1668.520 1688.110 1668.780 1688.430 ;
        RECT 1383.320 1687.770 1383.580 1688.090 ;
        RECT 1383.380 20.730 1383.520 1687.770 ;
        RECT 1376.420 20.410 1376.680 20.730 ;
        RECT 1383.320 20.410 1383.580 20.730 ;
        RECT 1376.480 2.400 1376.620 20.410 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1438.565 1686.485 1438.735 1688.355 ;
        RECT 1631.305 1686.825 1631.475 1688.355 ;
      LAYER mcon ;
        RECT 1438.565 1688.185 1438.735 1688.355 ;
        RECT 1631.305 1688.185 1631.475 1688.355 ;
      LAYER met1 ;
        RECT 1438.505 1688.340 1438.795 1688.385 ;
        RECT 1631.245 1688.340 1631.535 1688.385 ;
        RECT 1438.505 1688.200 1631.535 1688.340 ;
        RECT 1438.505 1688.155 1438.795 1688.200 ;
        RECT 1631.245 1688.155 1631.535 1688.200 ;
        RECT 1631.245 1686.980 1631.535 1687.025 ;
        RECT 1672.630 1686.980 1672.950 1687.040 ;
        RECT 1631.245 1686.840 1672.950 1686.980 ;
        RECT 1631.245 1686.795 1631.535 1686.840 ;
        RECT 1672.630 1686.780 1672.950 1686.840 ;
        RECT 1399.850 1686.640 1400.170 1686.700 ;
        RECT 1438.505 1686.640 1438.795 1686.685 ;
        RECT 1399.850 1686.500 1438.795 1686.640 ;
        RECT 1399.850 1686.440 1400.170 1686.500 ;
        RECT 1438.505 1686.455 1438.795 1686.500 ;
        RECT 1394.330 20.640 1394.650 20.700 ;
        RECT 1399.850 20.640 1400.170 20.700 ;
        RECT 1394.330 20.500 1400.170 20.640 ;
        RECT 1394.330 20.440 1394.650 20.500 ;
        RECT 1399.850 20.440 1400.170 20.500 ;
      LAYER via ;
        RECT 1672.660 1686.780 1672.920 1687.040 ;
        RECT 1399.880 1686.440 1400.140 1686.700 ;
        RECT 1394.360 20.440 1394.620 20.700 ;
        RECT 1399.880 20.440 1400.140 20.700 ;
      LAYER met2 ;
        RECT 1674.885 1700.410 1675.165 1704.000 ;
        RECT 1673.180 1700.270 1675.165 1700.410 ;
        RECT 1673.180 1688.850 1673.320 1700.270 ;
        RECT 1674.885 1700.000 1675.165 1700.270 ;
        RECT 1672.720 1688.710 1673.320 1688.850 ;
        RECT 1672.720 1687.070 1672.860 1688.710 ;
        RECT 1672.660 1686.750 1672.920 1687.070 ;
        RECT 1399.880 1686.410 1400.140 1686.730 ;
        RECT 1399.940 20.730 1400.080 1686.410 ;
        RECT 1394.360 20.410 1394.620 20.730 ;
        RECT 1399.880 20.410 1400.140 20.730 ;
        RECT 1394.420 2.400 1394.560 20.410 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1454.665 16.745 1454.835 17.595 ;
        RECT 1631.765 16.745 1631.935 17.595 ;
      LAYER mcon ;
        RECT 1454.665 17.425 1454.835 17.595 ;
        RECT 1631.765 17.425 1631.935 17.595 ;
      LAYER met1 ;
        RECT 1674.010 1686.980 1674.330 1687.040 ;
        RECT 1681.830 1686.980 1682.150 1687.040 ;
        RECT 1674.010 1686.840 1682.150 1686.980 ;
        RECT 1674.010 1686.780 1674.330 1686.840 ;
        RECT 1681.830 1686.780 1682.150 1686.840 ;
        RECT 1454.605 17.580 1454.895 17.625 ;
        RECT 1631.705 17.580 1631.995 17.625 ;
        RECT 1674.010 17.580 1674.330 17.640 ;
        RECT 1454.605 17.440 1631.995 17.580 ;
        RECT 1454.605 17.395 1454.895 17.440 ;
        RECT 1631.705 17.395 1631.995 17.440 ;
        RECT 1656.620 17.440 1674.330 17.580 ;
        RECT 1454.605 16.900 1454.895 16.945 ;
        RECT 1439.040 16.760 1454.895 16.900 ;
        RECT 1412.270 15.880 1412.590 15.940 ;
        RECT 1439.040 15.880 1439.180 16.760 ;
        RECT 1454.605 16.715 1454.895 16.760 ;
        RECT 1631.705 16.900 1631.995 16.945 ;
        RECT 1656.620 16.900 1656.760 17.440 ;
        RECT 1674.010 17.380 1674.330 17.440 ;
        RECT 1631.705 16.760 1656.760 16.900 ;
        RECT 1631.705 16.715 1631.995 16.760 ;
        RECT 1412.270 15.740 1439.180 15.880 ;
        RECT 1412.270 15.680 1412.590 15.740 ;
      LAYER via ;
        RECT 1674.040 1686.780 1674.300 1687.040 ;
        RECT 1681.860 1686.780 1682.120 1687.040 ;
        RECT 1412.300 15.680 1412.560 15.940 ;
        RECT 1674.040 17.380 1674.300 17.640 ;
      LAYER met2 ;
        RECT 1681.785 1700.000 1682.065 1704.000 ;
        RECT 1681.920 1687.070 1682.060 1700.000 ;
        RECT 1674.040 1686.750 1674.300 1687.070 ;
        RECT 1681.860 1686.750 1682.120 1687.070 ;
        RECT 1674.100 17.670 1674.240 1686.750 ;
        RECT 1674.040 17.350 1674.300 17.670 ;
        RECT 1412.300 15.650 1412.560 15.970 ;
        RECT 1412.360 2.400 1412.500 15.650 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1684.665 241.485 1684.835 289.595 ;
        RECT 1632.225 16.065 1632.395 18.615 ;
      LAYER mcon ;
        RECT 1684.665 289.425 1684.835 289.595 ;
        RECT 1632.225 18.445 1632.395 18.615 ;
      LAYER met1 ;
        RECT 1684.590 303.520 1684.910 303.580 ;
        RECT 1685.510 303.520 1685.830 303.580 ;
        RECT 1684.590 303.380 1685.830 303.520 ;
        RECT 1684.590 303.320 1684.910 303.380 ;
        RECT 1685.510 303.320 1685.830 303.380 ;
        RECT 1684.605 289.580 1684.895 289.625 ;
        RECT 1685.510 289.580 1685.830 289.640 ;
        RECT 1684.605 289.440 1685.830 289.580 ;
        RECT 1684.605 289.395 1684.895 289.440 ;
        RECT 1685.510 289.380 1685.830 289.440 ;
        RECT 1684.590 241.640 1684.910 241.700 ;
        RECT 1684.395 241.500 1684.910 241.640 ;
        RECT 1684.590 241.440 1684.910 241.500 ;
        RECT 1429.750 18.600 1430.070 18.660 ;
        RECT 1632.165 18.600 1632.455 18.645 ;
        RECT 1429.750 18.460 1632.455 18.600 ;
        RECT 1429.750 18.400 1430.070 18.460 ;
        RECT 1632.165 18.415 1632.455 18.460 ;
        RECT 1632.165 16.220 1632.455 16.265 ;
        RECT 1684.590 16.220 1684.910 16.280 ;
        RECT 1632.165 16.080 1684.910 16.220 ;
        RECT 1632.165 16.035 1632.455 16.080 ;
        RECT 1684.590 16.020 1684.910 16.080 ;
      LAYER via ;
        RECT 1684.620 303.320 1684.880 303.580 ;
        RECT 1685.540 303.320 1685.800 303.580 ;
        RECT 1685.540 289.380 1685.800 289.640 ;
        RECT 1684.620 241.440 1684.880 241.700 ;
        RECT 1429.780 18.400 1430.040 18.660 ;
        RECT 1684.620 16.020 1684.880 16.280 ;
      LAYER met2 ;
        RECT 1688.685 1701.090 1688.965 1704.000 ;
        RECT 1686.980 1700.950 1688.965 1701.090 ;
        RECT 1686.980 1688.170 1687.120 1700.950 ;
        RECT 1688.685 1700.000 1688.965 1700.950 ;
        RECT 1684.680 1688.030 1687.120 1688.170 ;
        RECT 1684.680 303.610 1684.820 1688.030 ;
        RECT 1684.620 303.290 1684.880 303.610 ;
        RECT 1685.540 303.290 1685.800 303.610 ;
        RECT 1685.600 289.670 1685.740 303.290 ;
        RECT 1685.540 289.350 1685.800 289.670 ;
        RECT 1684.620 241.410 1684.880 241.730 ;
        RECT 1684.680 241.245 1684.820 241.410 ;
        RECT 1684.610 240.875 1684.890 241.245 ;
        RECT 1685.070 240.195 1685.350 240.565 ;
        RECT 1685.140 110.570 1685.280 240.195 ;
        RECT 1684.680 110.430 1685.280 110.570 ;
        RECT 1429.780 18.370 1430.040 18.690 ;
        RECT 1429.840 2.400 1429.980 18.370 ;
        RECT 1684.680 16.310 1684.820 110.430 ;
        RECT 1684.620 15.990 1684.880 16.310 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
      LAYER via2 ;
        RECT 1684.610 240.920 1684.890 241.200 ;
        RECT 1685.070 240.240 1685.350 240.520 ;
      LAYER met3 ;
        RECT 1684.585 241.210 1684.915 241.225 ;
        RECT 1683.910 240.910 1684.915 241.210 ;
        RECT 1683.910 240.530 1684.210 240.910 ;
        RECT 1684.585 240.895 1684.915 240.910 ;
        RECT 1685.045 240.530 1685.375 240.545 ;
        RECT 1683.910 240.230 1685.375 240.530 ;
        RECT 1685.045 240.215 1685.375 240.230 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1683.285 1684.445 1683.455 1685.295 ;
      LAYER mcon ;
        RECT 1683.285 1685.125 1683.455 1685.295 ;
      LAYER met1 ;
        RECT 1683.225 1685.280 1683.515 1685.325 ;
        RECT 1695.170 1685.280 1695.490 1685.340 ;
        RECT 1683.225 1685.140 1695.490 1685.280 ;
        RECT 1683.225 1685.095 1683.515 1685.140 ;
        RECT 1695.170 1685.080 1695.490 1685.140 ;
        RECT 1583.850 1684.600 1584.170 1684.660 ;
        RECT 1683.225 1684.600 1683.515 1684.645 ;
        RECT 1583.850 1684.460 1683.515 1684.600 ;
        RECT 1583.850 1684.400 1584.170 1684.460 ;
        RECT 1683.225 1684.415 1683.515 1684.460 ;
        RECT 1447.690 15.880 1448.010 15.940 ;
        RECT 1582.930 15.880 1583.250 15.940 ;
        RECT 1447.690 15.740 1583.250 15.880 ;
        RECT 1447.690 15.680 1448.010 15.740 ;
        RECT 1582.930 15.680 1583.250 15.740 ;
      LAYER via ;
        RECT 1695.200 1685.080 1695.460 1685.340 ;
        RECT 1583.880 1684.400 1584.140 1684.660 ;
        RECT 1447.720 15.680 1447.980 15.940 ;
        RECT 1582.960 15.680 1583.220 15.940 ;
      LAYER met2 ;
        RECT 1695.125 1700.000 1695.405 1704.000 ;
        RECT 1695.260 1685.370 1695.400 1700.000 ;
        RECT 1695.200 1685.050 1695.460 1685.370 ;
        RECT 1583.880 1684.370 1584.140 1684.690 ;
        RECT 1583.940 1666.410 1584.080 1684.370 ;
        RECT 1583.480 1666.270 1584.080 1666.410 ;
        RECT 1583.480 24.890 1583.620 1666.270 ;
        RECT 1583.020 24.750 1583.620 24.890 ;
        RECT 1583.020 15.970 1583.160 24.750 ;
        RECT 1447.720 15.650 1447.980 15.970 ;
        RECT 1582.960 15.650 1583.220 15.970 ;
        RECT 1447.780 2.400 1447.920 15.650 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1465.630 19.620 1465.950 19.680 ;
        RECT 1698.390 19.620 1698.710 19.680 ;
        RECT 1465.630 19.480 1698.710 19.620 ;
        RECT 1465.630 19.420 1465.950 19.480 ;
        RECT 1698.390 19.420 1698.710 19.480 ;
      LAYER via ;
        RECT 1465.660 19.420 1465.920 19.680 ;
        RECT 1698.420 19.420 1698.680 19.680 ;
      LAYER met2 ;
        RECT 1702.025 1700.410 1702.305 1704.000 ;
        RECT 1700.780 1700.270 1702.305 1700.410 ;
        RECT 1700.780 1688.680 1700.920 1700.270 ;
        RECT 1702.025 1700.000 1702.305 1700.270 ;
        RECT 1698.480 1688.540 1700.920 1688.680 ;
        RECT 1698.480 19.710 1698.620 1688.540 ;
        RECT 1465.660 19.390 1465.920 19.710 ;
        RECT 1698.420 19.390 1698.680 19.710 ;
        RECT 1465.720 2.400 1465.860 19.390 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1517.225 1685.805 1517.395 1690.395 ;
      LAYER mcon ;
        RECT 1517.225 1690.225 1517.395 1690.395 ;
      LAYER met1 ;
        RECT 1517.165 1690.380 1517.455 1690.425 ;
        RECT 1708.970 1690.380 1709.290 1690.440 ;
        RECT 1517.165 1690.240 1709.290 1690.380 ;
        RECT 1517.165 1690.195 1517.455 1690.240 ;
        RECT 1708.970 1690.180 1709.290 1690.240 ;
        RECT 1489.550 1685.960 1489.870 1686.020 ;
        RECT 1517.165 1685.960 1517.455 1686.005 ;
        RECT 1489.550 1685.820 1517.455 1685.960 ;
        RECT 1489.550 1685.760 1489.870 1685.820 ;
        RECT 1517.165 1685.775 1517.455 1685.820 ;
        RECT 1483.570 20.640 1483.890 20.700 ;
        RECT 1489.550 20.640 1489.870 20.700 ;
        RECT 1483.570 20.500 1489.870 20.640 ;
        RECT 1483.570 20.440 1483.890 20.500 ;
        RECT 1489.550 20.440 1489.870 20.500 ;
      LAYER via ;
        RECT 1709.000 1690.180 1709.260 1690.440 ;
        RECT 1489.580 1685.760 1489.840 1686.020 ;
        RECT 1483.600 20.440 1483.860 20.700 ;
        RECT 1489.580 20.440 1489.840 20.700 ;
      LAYER met2 ;
        RECT 1708.925 1700.000 1709.205 1704.000 ;
        RECT 1709.060 1690.470 1709.200 1700.000 ;
        RECT 1709.000 1690.150 1709.260 1690.470 ;
        RECT 1489.580 1685.730 1489.840 1686.050 ;
        RECT 1489.640 20.730 1489.780 1685.730 ;
        RECT 1483.600 20.410 1483.860 20.730 ;
        RECT 1489.580 20.410 1489.840 20.730 ;
        RECT 1483.660 2.400 1483.800 20.410 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1715.410 1685.620 1715.730 1685.680 ;
        RECT 1631.780 1685.480 1715.730 1685.620 ;
        RECT 1597.650 1684.940 1597.970 1685.000 ;
        RECT 1631.780 1684.940 1631.920 1685.480 ;
        RECT 1715.410 1685.420 1715.730 1685.480 ;
        RECT 1597.650 1684.800 1631.920 1684.940 ;
        RECT 1597.650 1684.740 1597.970 1684.800 ;
        RECT 1597.190 15.540 1597.510 15.600 ;
        RECT 1566.460 15.400 1597.510 15.540 ;
        RECT 1501.510 15.200 1501.830 15.260 ;
        RECT 1566.460 15.200 1566.600 15.400 ;
        RECT 1597.190 15.340 1597.510 15.400 ;
        RECT 1501.510 15.060 1566.600 15.200 ;
        RECT 1501.510 15.000 1501.830 15.060 ;
      LAYER via ;
        RECT 1597.680 1684.740 1597.940 1685.000 ;
        RECT 1715.440 1685.420 1715.700 1685.680 ;
        RECT 1501.540 15.000 1501.800 15.260 ;
        RECT 1597.220 15.340 1597.480 15.600 ;
      LAYER met2 ;
        RECT 1715.365 1700.000 1715.645 1704.000 ;
        RECT 1715.500 1685.710 1715.640 1700.000 ;
        RECT 1715.440 1685.390 1715.700 1685.710 ;
        RECT 1597.680 1684.710 1597.940 1685.030 ;
        RECT 1597.740 1670.490 1597.880 1684.710 ;
        RECT 1597.280 1670.350 1597.880 1670.490 ;
        RECT 1597.280 15.630 1597.420 1670.350 ;
        RECT 1597.220 15.310 1597.480 15.630 ;
        RECT 1501.540 14.970 1501.800 15.290 ;
        RECT 1501.600 2.400 1501.740 14.970 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1632.225 1683.765 1632.395 1685.295 ;
        RECT 1682.825 1685.125 1682.995 1690.055 ;
      LAYER mcon ;
        RECT 1682.825 1689.885 1682.995 1690.055 ;
        RECT 1632.225 1685.125 1632.395 1685.295 ;
      LAYER met1 ;
        RECT 1682.765 1690.040 1683.055 1690.085 ;
        RECT 1722.310 1690.040 1722.630 1690.100 ;
        RECT 1682.765 1689.900 1722.630 1690.040 ;
        RECT 1682.765 1689.855 1683.055 1689.900 ;
        RECT 1722.310 1689.840 1722.630 1689.900 ;
        RECT 1632.165 1685.280 1632.455 1685.325 ;
        RECT 1682.765 1685.280 1683.055 1685.325 ;
        RECT 1632.165 1685.140 1683.055 1685.280 ;
        RECT 1632.165 1685.095 1632.455 1685.140 ;
        RECT 1682.765 1685.095 1683.055 1685.140 ;
        RECT 1611.450 1683.920 1611.770 1683.980 ;
        RECT 1632.165 1683.920 1632.455 1683.965 ;
        RECT 1611.450 1683.780 1632.455 1683.920 ;
        RECT 1611.450 1683.720 1611.770 1683.780 ;
        RECT 1632.165 1683.735 1632.455 1683.780 ;
        RECT 1518.990 14.860 1519.310 14.920 ;
        RECT 1610.990 14.860 1611.310 14.920 ;
        RECT 1518.990 14.720 1611.310 14.860 ;
        RECT 1518.990 14.660 1519.310 14.720 ;
        RECT 1610.990 14.660 1611.310 14.720 ;
      LAYER via ;
        RECT 1722.340 1689.840 1722.600 1690.100 ;
        RECT 1611.480 1683.720 1611.740 1683.980 ;
        RECT 1519.020 14.660 1519.280 14.920 ;
        RECT 1611.020 14.660 1611.280 14.920 ;
      LAYER met2 ;
        RECT 1722.265 1700.000 1722.545 1704.000 ;
        RECT 1722.400 1690.130 1722.540 1700.000 ;
        RECT 1722.340 1689.810 1722.600 1690.130 ;
        RECT 1611.480 1683.690 1611.740 1684.010 ;
        RECT 1611.540 1670.490 1611.680 1683.690 ;
        RECT 1611.080 1670.350 1611.680 1670.490 ;
        RECT 1611.080 14.950 1611.220 1670.350 ;
        RECT 1519.020 14.630 1519.280 14.950 ;
        RECT 1611.020 14.630 1611.280 14.950 ;
        RECT 1519.080 2.400 1519.220 14.630 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1415.030 1678.140 1415.350 1678.200 ;
        RECT 1417.790 1678.140 1418.110 1678.200 ;
        RECT 1415.030 1678.000 1418.110 1678.140 ;
        RECT 1415.030 1677.940 1415.350 1678.000 ;
        RECT 1417.790 1677.940 1418.110 1678.000 ;
        RECT 716.290 46.820 716.610 46.880 ;
        RECT 1415.030 46.820 1415.350 46.880 ;
        RECT 716.290 46.680 1415.350 46.820 ;
        RECT 716.290 46.620 716.610 46.680 ;
        RECT 1415.030 46.620 1415.350 46.680 ;
      LAYER via ;
        RECT 1415.060 1677.940 1415.320 1678.200 ;
        RECT 1417.820 1677.940 1418.080 1678.200 ;
        RECT 716.320 46.620 716.580 46.880 ;
        RECT 1415.060 46.620 1415.320 46.880 ;
      LAYER met2 ;
        RECT 1419.125 1700.410 1419.405 1704.000 ;
        RECT 1417.880 1700.270 1419.405 1700.410 ;
        RECT 1417.880 1678.230 1418.020 1700.270 ;
        RECT 1419.125 1700.000 1419.405 1700.270 ;
        RECT 1415.060 1677.910 1415.320 1678.230 ;
        RECT 1417.820 1677.910 1418.080 1678.230 ;
        RECT 1415.120 46.910 1415.260 1677.910 ;
        RECT 716.320 46.590 716.580 46.910 ;
        RECT 1415.060 46.590 1415.320 46.910 ;
        RECT 716.380 2.400 716.520 46.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1726.065 1545.725 1726.235 1593.835 ;
        RECT 1726.065 1401.225 1726.235 1448.995 ;
        RECT 1726.065 1304.665 1726.235 1352.435 ;
        RECT 1726.065 1207.425 1726.235 1255.875 ;
        RECT 1725.145 963.645 1725.315 1007.335 ;
        RECT 1726.065 724.625 1726.235 814.215 ;
        RECT 1726.065 572.645 1726.235 620.755 ;
        RECT 1726.065 493.425 1726.235 524.195 ;
        RECT 1726.065 379.525 1726.235 469.115 ;
        RECT 1726.065 282.965 1726.235 331.075 ;
        RECT 1726.065 144.925 1726.235 234.515 ;
        RECT 1726.065 48.365 1726.235 137.955 ;
      LAYER mcon ;
        RECT 1726.065 1593.665 1726.235 1593.835 ;
        RECT 1726.065 1448.825 1726.235 1448.995 ;
        RECT 1726.065 1352.265 1726.235 1352.435 ;
        RECT 1726.065 1255.705 1726.235 1255.875 ;
        RECT 1725.145 1007.165 1725.315 1007.335 ;
        RECT 1726.065 814.045 1726.235 814.215 ;
        RECT 1726.065 620.585 1726.235 620.755 ;
        RECT 1726.065 524.025 1726.235 524.195 ;
        RECT 1726.065 468.945 1726.235 469.115 ;
        RECT 1726.065 330.905 1726.235 331.075 ;
        RECT 1726.065 234.345 1726.235 234.515 ;
        RECT 1726.065 137.785 1726.235 137.955 ;
      LAYER met1 ;
        RECT 1725.990 1695.480 1726.310 1695.540 ;
        RECT 1728.750 1695.480 1729.070 1695.540 ;
        RECT 1725.990 1695.340 1729.070 1695.480 ;
        RECT 1725.990 1695.280 1726.310 1695.340 ;
        RECT 1728.750 1695.280 1729.070 1695.340 ;
        RECT 1725.990 1593.820 1726.310 1593.880 ;
        RECT 1725.795 1593.680 1726.310 1593.820 ;
        RECT 1725.990 1593.620 1726.310 1593.680 ;
        RECT 1726.005 1545.880 1726.295 1545.925 ;
        RECT 1726.450 1545.880 1726.770 1545.940 ;
        RECT 1726.005 1545.740 1726.770 1545.880 ;
        RECT 1726.005 1545.695 1726.295 1545.740 ;
        RECT 1726.450 1545.680 1726.770 1545.740 ;
        RECT 1725.990 1448.980 1726.310 1449.040 ;
        RECT 1725.795 1448.840 1726.310 1448.980 ;
        RECT 1725.990 1448.780 1726.310 1448.840 ;
        RECT 1725.990 1401.380 1726.310 1401.440 ;
        RECT 1725.795 1401.240 1726.310 1401.380 ;
        RECT 1725.990 1401.180 1726.310 1401.240 ;
        RECT 1725.990 1352.420 1726.310 1352.480 ;
        RECT 1725.795 1352.280 1726.310 1352.420 ;
        RECT 1725.990 1352.220 1726.310 1352.280 ;
        RECT 1725.990 1304.820 1726.310 1304.880 ;
        RECT 1725.795 1304.680 1726.310 1304.820 ;
        RECT 1725.990 1304.620 1726.310 1304.680 ;
        RECT 1725.990 1255.860 1726.310 1255.920 ;
        RECT 1725.795 1255.720 1726.310 1255.860 ;
        RECT 1725.990 1255.660 1726.310 1255.720 ;
        RECT 1725.990 1207.580 1726.310 1207.640 ;
        RECT 1725.795 1207.440 1726.310 1207.580 ;
        RECT 1725.990 1207.380 1726.310 1207.440 ;
        RECT 1726.910 1159.440 1727.230 1159.700 ;
        RECT 1726.450 1159.300 1726.770 1159.360 ;
        RECT 1727.000 1159.300 1727.140 1159.440 ;
        RECT 1726.450 1159.160 1727.140 1159.300 ;
        RECT 1726.450 1159.100 1726.770 1159.160 ;
        RECT 1725.990 1111.020 1726.310 1111.080 ;
        RECT 1726.450 1111.020 1726.770 1111.080 ;
        RECT 1725.990 1110.880 1726.770 1111.020 ;
        RECT 1725.990 1110.820 1726.310 1110.880 ;
        RECT 1726.450 1110.820 1726.770 1110.880 ;
        RECT 1726.910 1062.880 1727.230 1063.140 ;
        RECT 1726.450 1062.740 1726.770 1062.800 ;
        RECT 1727.000 1062.740 1727.140 1062.880 ;
        RECT 1726.450 1062.600 1727.140 1062.740 ;
        RECT 1726.450 1062.540 1726.770 1062.600 ;
        RECT 1725.085 1007.320 1725.375 1007.365 ;
        RECT 1725.990 1007.320 1726.310 1007.380 ;
        RECT 1725.085 1007.180 1726.310 1007.320 ;
        RECT 1725.085 1007.135 1725.375 1007.180 ;
        RECT 1725.990 1007.120 1726.310 1007.180 ;
        RECT 1725.070 963.800 1725.390 963.860 ;
        RECT 1724.875 963.660 1725.390 963.800 ;
        RECT 1725.070 963.600 1725.390 963.660 ;
        RECT 1725.070 953.260 1725.390 953.320 ;
        RECT 1726.450 953.260 1726.770 953.320 ;
        RECT 1725.070 953.120 1726.770 953.260 ;
        RECT 1725.070 953.060 1725.390 953.120 ;
        RECT 1726.450 953.060 1726.770 953.120 ;
        RECT 1725.070 855.340 1725.390 855.400 ;
        RECT 1725.990 855.340 1726.310 855.400 ;
        RECT 1725.070 855.200 1726.310 855.340 ;
        RECT 1725.070 855.140 1725.390 855.200 ;
        RECT 1725.990 855.140 1726.310 855.200 ;
        RECT 1725.990 814.200 1726.310 814.260 ;
        RECT 1725.795 814.060 1726.310 814.200 ;
        RECT 1725.990 814.000 1726.310 814.060 ;
        RECT 1726.005 724.780 1726.295 724.825 ;
        RECT 1726.450 724.780 1726.770 724.840 ;
        RECT 1726.005 724.640 1726.770 724.780 ;
        RECT 1726.005 724.595 1726.295 724.640 ;
        RECT 1726.450 724.580 1726.770 724.640 ;
        RECT 1725.990 717.640 1726.310 717.700 ;
        RECT 1726.910 717.640 1727.230 717.700 ;
        RECT 1725.990 717.500 1727.230 717.640 ;
        RECT 1725.990 717.440 1726.310 717.500 ;
        RECT 1726.910 717.440 1727.230 717.500 ;
        RECT 1725.990 628.220 1726.310 628.280 ;
        RECT 1726.910 628.220 1727.230 628.280 ;
        RECT 1725.990 628.080 1727.230 628.220 ;
        RECT 1725.990 628.020 1726.310 628.080 ;
        RECT 1726.910 628.020 1727.230 628.080 ;
        RECT 1725.990 620.740 1726.310 620.800 ;
        RECT 1725.795 620.600 1726.310 620.740 ;
        RECT 1725.990 620.540 1726.310 620.600 ;
        RECT 1725.990 572.800 1726.310 572.860 ;
        RECT 1725.795 572.660 1726.310 572.800 ;
        RECT 1725.990 572.600 1726.310 572.660 ;
        RECT 1725.990 524.180 1726.310 524.240 ;
        RECT 1725.795 524.040 1726.310 524.180 ;
        RECT 1725.990 523.980 1726.310 524.040 ;
        RECT 1726.005 493.580 1726.295 493.625 ;
        RECT 1726.910 493.580 1727.230 493.640 ;
        RECT 1726.005 493.440 1727.230 493.580 ;
        RECT 1726.005 493.395 1726.295 493.440 ;
        RECT 1726.910 493.380 1727.230 493.440 ;
        RECT 1726.005 469.100 1726.295 469.145 ;
        RECT 1726.910 469.100 1727.230 469.160 ;
        RECT 1726.005 468.960 1727.230 469.100 ;
        RECT 1726.005 468.915 1726.295 468.960 ;
        RECT 1726.910 468.900 1727.230 468.960 ;
        RECT 1725.990 379.680 1726.310 379.740 ;
        RECT 1725.795 379.540 1726.310 379.680 ;
        RECT 1725.990 379.480 1726.310 379.540 ;
        RECT 1725.990 331.060 1726.310 331.120 ;
        RECT 1725.795 330.920 1726.310 331.060 ;
        RECT 1725.990 330.860 1726.310 330.920 ;
        RECT 1725.990 283.120 1726.310 283.180 ;
        RECT 1725.795 282.980 1726.310 283.120 ;
        RECT 1725.990 282.920 1726.310 282.980 ;
        RECT 1725.990 234.500 1726.310 234.560 ;
        RECT 1725.795 234.360 1726.310 234.500 ;
        RECT 1725.990 234.300 1726.310 234.360 ;
        RECT 1726.005 145.080 1726.295 145.125 ;
        RECT 1726.450 145.080 1726.770 145.140 ;
        RECT 1726.005 144.940 1726.770 145.080 ;
        RECT 1726.005 144.895 1726.295 144.940 ;
        RECT 1726.450 144.880 1726.770 144.940 ;
        RECT 1726.005 137.940 1726.295 137.985 ;
        RECT 1726.450 137.940 1726.770 138.000 ;
        RECT 1726.005 137.800 1726.770 137.940 ;
        RECT 1726.005 137.755 1726.295 137.800 ;
        RECT 1726.450 137.740 1726.770 137.800 ;
        RECT 1725.990 48.520 1726.310 48.580 ;
        RECT 1725.795 48.380 1726.310 48.520 ;
        RECT 1725.990 48.320 1726.310 48.380 ;
        RECT 1721.020 20.840 1725.300 20.980 ;
        RECT 1536.930 20.640 1537.250 20.700 ;
        RECT 1721.020 20.640 1721.160 20.840 ;
        RECT 1536.930 20.500 1721.160 20.640 ;
        RECT 1725.160 20.640 1725.300 20.840 ;
        RECT 1725.990 20.640 1726.310 20.700 ;
        RECT 1725.160 20.500 1726.310 20.640 ;
        RECT 1536.930 20.440 1537.250 20.500 ;
        RECT 1725.990 20.440 1726.310 20.500 ;
      LAYER via ;
        RECT 1726.020 1695.280 1726.280 1695.540 ;
        RECT 1728.780 1695.280 1729.040 1695.540 ;
        RECT 1726.020 1593.620 1726.280 1593.880 ;
        RECT 1726.480 1545.680 1726.740 1545.940 ;
        RECT 1726.020 1448.780 1726.280 1449.040 ;
        RECT 1726.020 1401.180 1726.280 1401.440 ;
        RECT 1726.020 1352.220 1726.280 1352.480 ;
        RECT 1726.020 1304.620 1726.280 1304.880 ;
        RECT 1726.020 1255.660 1726.280 1255.920 ;
        RECT 1726.020 1207.380 1726.280 1207.640 ;
        RECT 1726.940 1159.440 1727.200 1159.700 ;
        RECT 1726.480 1159.100 1726.740 1159.360 ;
        RECT 1726.020 1110.820 1726.280 1111.080 ;
        RECT 1726.480 1110.820 1726.740 1111.080 ;
        RECT 1726.940 1062.880 1727.200 1063.140 ;
        RECT 1726.480 1062.540 1726.740 1062.800 ;
        RECT 1726.020 1007.120 1726.280 1007.380 ;
        RECT 1725.100 963.600 1725.360 963.860 ;
        RECT 1725.100 953.060 1725.360 953.320 ;
        RECT 1726.480 953.060 1726.740 953.320 ;
        RECT 1725.100 855.140 1725.360 855.400 ;
        RECT 1726.020 855.140 1726.280 855.400 ;
        RECT 1726.020 814.000 1726.280 814.260 ;
        RECT 1726.480 724.580 1726.740 724.840 ;
        RECT 1726.020 717.440 1726.280 717.700 ;
        RECT 1726.940 717.440 1727.200 717.700 ;
        RECT 1726.020 628.020 1726.280 628.280 ;
        RECT 1726.940 628.020 1727.200 628.280 ;
        RECT 1726.020 620.540 1726.280 620.800 ;
        RECT 1726.020 572.600 1726.280 572.860 ;
        RECT 1726.020 523.980 1726.280 524.240 ;
        RECT 1726.940 493.380 1727.200 493.640 ;
        RECT 1726.940 468.900 1727.200 469.160 ;
        RECT 1726.020 379.480 1726.280 379.740 ;
        RECT 1726.020 330.860 1726.280 331.120 ;
        RECT 1726.020 282.920 1726.280 283.180 ;
        RECT 1726.020 234.300 1726.280 234.560 ;
        RECT 1726.480 144.880 1726.740 145.140 ;
        RECT 1726.480 137.740 1726.740 138.000 ;
        RECT 1726.020 48.320 1726.280 48.580 ;
        RECT 1536.960 20.440 1537.220 20.700 ;
        RECT 1726.020 20.440 1726.280 20.700 ;
      LAYER met2 ;
        RECT 1728.705 1700.000 1728.985 1704.000 ;
        RECT 1728.840 1695.570 1728.980 1700.000 ;
        RECT 1726.020 1695.250 1726.280 1695.570 ;
        RECT 1728.780 1695.250 1729.040 1695.570 ;
        RECT 1726.080 1645.330 1726.220 1695.250 ;
        RECT 1726.080 1645.190 1726.680 1645.330 ;
        RECT 1726.540 1642.610 1726.680 1645.190 ;
        RECT 1726.080 1642.470 1726.680 1642.610 ;
        RECT 1726.080 1593.910 1726.220 1642.470 ;
        RECT 1726.020 1593.590 1726.280 1593.910 ;
        RECT 1726.480 1545.880 1726.740 1545.970 ;
        RECT 1726.080 1545.740 1726.740 1545.880 ;
        RECT 1726.080 1449.070 1726.220 1545.740 ;
        RECT 1726.480 1545.650 1726.740 1545.740 ;
        RECT 1726.020 1448.750 1726.280 1449.070 ;
        RECT 1726.020 1401.150 1726.280 1401.470 ;
        RECT 1726.080 1400.700 1726.220 1401.150 ;
        RECT 1726.080 1400.560 1726.680 1400.700 ;
        RECT 1726.540 1352.930 1726.680 1400.560 ;
        RECT 1726.080 1352.790 1726.680 1352.930 ;
        RECT 1726.080 1352.510 1726.220 1352.790 ;
        RECT 1726.020 1352.190 1726.280 1352.510 ;
        RECT 1726.020 1304.590 1726.280 1304.910 ;
        RECT 1726.080 1304.140 1726.220 1304.590 ;
        RECT 1726.080 1304.000 1726.680 1304.140 ;
        RECT 1726.540 1257.165 1726.680 1304.000 ;
        RECT 1726.470 1256.795 1726.750 1257.165 ;
        RECT 1726.010 1256.115 1726.290 1256.485 ;
        RECT 1726.080 1255.950 1726.220 1256.115 ;
        RECT 1726.020 1255.630 1726.280 1255.950 ;
        RECT 1726.080 1207.670 1726.220 1207.825 ;
        RECT 1726.020 1207.410 1726.280 1207.670 ;
        RECT 1726.020 1207.350 1727.140 1207.410 ;
        RECT 1726.080 1207.270 1727.140 1207.350 ;
        RECT 1727.000 1159.730 1727.140 1207.270 ;
        RECT 1726.940 1159.410 1727.200 1159.730 ;
        RECT 1726.480 1159.070 1726.740 1159.390 ;
        RECT 1726.080 1111.110 1726.220 1111.265 ;
        RECT 1726.540 1111.110 1726.680 1159.070 ;
        RECT 1726.020 1110.850 1726.280 1111.110 ;
        RECT 1726.480 1110.850 1726.740 1111.110 ;
        RECT 1726.020 1110.790 1727.140 1110.850 ;
        RECT 1726.080 1110.710 1727.140 1110.790 ;
        RECT 1727.000 1063.170 1727.140 1110.710 ;
        RECT 1726.940 1062.850 1727.200 1063.170 ;
        RECT 1726.480 1062.510 1726.740 1062.830 ;
        RECT 1726.540 1014.460 1726.680 1062.510 ;
        RECT 1726.080 1014.320 1726.680 1014.460 ;
        RECT 1726.080 1007.410 1726.220 1014.320 ;
        RECT 1726.020 1007.090 1726.280 1007.410 ;
        RECT 1725.100 963.570 1725.360 963.890 ;
        RECT 1725.160 953.350 1725.300 963.570 ;
        RECT 1725.100 953.030 1725.360 953.350 ;
        RECT 1726.480 953.030 1726.740 953.350 ;
        RECT 1726.540 862.765 1726.680 953.030 ;
        RECT 1725.090 862.395 1725.370 862.765 ;
        RECT 1726.470 862.395 1726.750 862.765 ;
        RECT 1725.160 855.430 1725.300 862.395 ;
        RECT 1725.100 855.110 1725.360 855.430 ;
        RECT 1726.020 855.110 1726.280 855.430 ;
        RECT 1726.080 814.290 1726.220 855.110 ;
        RECT 1726.020 813.970 1726.280 814.290 ;
        RECT 1726.480 724.610 1726.740 724.870 ;
        RECT 1726.080 724.550 1726.740 724.610 ;
        RECT 1726.080 724.470 1726.680 724.550 ;
        RECT 1726.080 717.730 1726.220 724.470 ;
        RECT 1726.020 717.410 1726.280 717.730 ;
        RECT 1726.940 717.410 1727.200 717.730 ;
        RECT 1727.000 628.310 1727.140 717.410 ;
        RECT 1726.020 627.990 1726.280 628.310 ;
        RECT 1726.940 627.990 1727.200 628.310 ;
        RECT 1726.080 620.830 1726.220 627.990 ;
        RECT 1726.020 620.510 1726.280 620.830 ;
        RECT 1726.020 572.570 1726.280 572.890 ;
        RECT 1726.080 524.270 1726.220 572.570 ;
        RECT 1726.020 523.950 1726.280 524.270 ;
        RECT 1726.940 493.350 1727.200 493.670 ;
        RECT 1727.000 469.190 1727.140 493.350 ;
        RECT 1726.940 468.870 1727.200 469.190 ;
        RECT 1726.020 379.450 1726.280 379.770 ;
        RECT 1726.080 331.150 1726.220 379.450 ;
        RECT 1726.020 330.830 1726.280 331.150 ;
        RECT 1726.020 282.890 1726.280 283.210 ;
        RECT 1726.080 234.590 1726.220 282.890 ;
        RECT 1726.020 234.270 1726.280 234.590 ;
        RECT 1726.480 144.850 1726.740 145.170 ;
        RECT 1726.540 138.030 1726.680 144.850 ;
        RECT 1726.480 137.710 1726.740 138.030 ;
        RECT 1726.020 48.290 1726.280 48.610 ;
        RECT 1726.080 20.730 1726.220 48.290 ;
        RECT 1536.960 20.410 1537.220 20.730 ;
        RECT 1726.020 20.410 1726.280 20.730 ;
        RECT 1537.020 2.400 1537.160 20.410 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
      LAYER via2 ;
        RECT 1726.470 1256.840 1726.750 1257.120 ;
        RECT 1726.010 1256.160 1726.290 1256.440 ;
        RECT 1725.090 862.440 1725.370 862.720 ;
        RECT 1726.470 862.440 1726.750 862.720 ;
      LAYER met3 ;
        RECT 1726.445 1257.130 1726.775 1257.145 ;
        RECT 1725.310 1256.830 1726.775 1257.130 ;
        RECT 1725.310 1256.450 1725.610 1256.830 ;
        RECT 1726.445 1256.815 1726.775 1256.830 ;
        RECT 1725.985 1256.450 1726.315 1256.465 ;
        RECT 1725.310 1256.150 1726.315 1256.450 ;
        RECT 1725.985 1256.135 1726.315 1256.150 ;
        RECT 1725.065 862.730 1725.395 862.745 ;
        RECT 1726.445 862.730 1726.775 862.745 ;
        RECT 1725.065 862.430 1726.775 862.730 ;
        RECT 1725.065 862.415 1725.395 862.430 ;
        RECT 1726.445 862.415 1726.775 862.430 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1709.045 1684.445 1709.215 1686.655 ;
      LAYER mcon ;
        RECT 1709.045 1686.485 1709.215 1686.655 ;
      LAYER met1 ;
        RECT 1708.985 1686.640 1709.275 1686.685 ;
        RECT 1735.650 1686.640 1735.970 1686.700 ;
        RECT 1708.985 1686.500 1735.970 1686.640 ;
        RECT 1708.985 1686.455 1709.275 1686.500 ;
        RECT 1735.650 1686.440 1735.970 1686.500 ;
        RECT 1708.985 1684.600 1709.275 1684.645 ;
        RECT 1683.760 1684.460 1709.275 1684.600 ;
        RECT 1631.690 1684.260 1632.010 1684.320 ;
        RECT 1683.760 1684.260 1683.900 1684.460 ;
        RECT 1708.985 1684.415 1709.275 1684.460 ;
        RECT 1631.690 1684.120 1683.900 1684.260 ;
        RECT 1631.690 1684.060 1632.010 1684.120 ;
        RECT 1630.770 14.860 1631.090 14.920 ;
        RECT 1613.840 14.720 1631.090 14.860 ;
        RECT 1554.870 14.520 1555.190 14.580 ;
        RECT 1613.840 14.520 1613.980 14.720 ;
        RECT 1630.770 14.660 1631.090 14.720 ;
        RECT 1554.870 14.380 1613.980 14.520 ;
        RECT 1554.870 14.320 1555.190 14.380 ;
      LAYER via ;
        RECT 1735.680 1686.440 1735.940 1686.700 ;
        RECT 1631.720 1684.060 1631.980 1684.320 ;
        RECT 1554.900 14.320 1555.160 14.580 ;
        RECT 1630.800 14.660 1631.060 14.920 ;
      LAYER met2 ;
        RECT 1735.605 1700.000 1735.885 1704.000 ;
        RECT 1735.740 1686.730 1735.880 1700.000 ;
        RECT 1735.680 1686.410 1735.940 1686.730 ;
        RECT 1631.720 1684.030 1631.980 1684.350 ;
        RECT 1631.780 23.700 1631.920 1684.030 ;
        RECT 1630.860 23.560 1631.920 23.700 ;
        RECT 1630.860 14.950 1631.000 23.560 ;
        RECT 1630.800 14.630 1631.060 14.950 ;
        RECT 1554.900 14.290 1555.160 14.610 ;
        RECT 1554.960 2.400 1555.100 14.290 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1739.865 1642.285 1740.035 1690.395 ;
        RECT 1739.865 1594.005 1740.035 1641.775 ;
        RECT 1739.865 1497.785 1740.035 1545.215 ;
        RECT 1739.865 1304.665 1740.035 1352.435 ;
        RECT 1739.865 1207.425 1740.035 1255.875 ;
        RECT 1739.865 580.125 1740.035 627.895 ;
        RECT 1739.865 483.565 1740.035 531.335 ;
        RECT 1739.865 324.445 1740.035 372.555 ;
        RECT 1739.405 228.225 1739.575 275.995 ;
        RECT 1656.145 17.085 1657.235 17.255 ;
      LAYER mcon ;
        RECT 1739.865 1690.225 1740.035 1690.395 ;
        RECT 1739.865 1641.605 1740.035 1641.775 ;
        RECT 1739.865 1545.045 1740.035 1545.215 ;
        RECT 1739.865 1352.265 1740.035 1352.435 ;
        RECT 1739.865 1255.705 1740.035 1255.875 ;
        RECT 1739.865 627.725 1740.035 627.895 ;
        RECT 1739.865 531.165 1740.035 531.335 ;
        RECT 1739.865 372.385 1740.035 372.555 ;
        RECT 1739.405 275.825 1739.575 275.995 ;
        RECT 1657.065 17.085 1657.235 17.255 ;
      LAYER met1 ;
        RECT 1739.805 1690.380 1740.095 1690.425 ;
        RECT 1741.170 1690.380 1741.490 1690.440 ;
        RECT 1739.805 1690.240 1741.490 1690.380 ;
        RECT 1739.805 1690.195 1740.095 1690.240 ;
        RECT 1741.170 1690.180 1741.490 1690.240 ;
        RECT 1739.790 1642.440 1740.110 1642.500 ;
        RECT 1739.595 1642.300 1740.110 1642.440 ;
        RECT 1739.790 1642.240 1740.110 1642.300 ;
        RECT 1739.790 1641.760 1740.110 1641.820 ;
        RECT 1739.595 1641.620 1740.110 1641.760 ;
        RECT 1739.790 1641.560 1740.110 1641.620 ;
        RECT 1739.790 1594.160 1740.110 1594.220 ;
        RECT 1739.595 1594.020 1740.110 1594.160 ;
        RECT 1739.790 1593.960 1740.110 1594.020 ;
        RECT 1739.790 1546.360 1740.110 1546.620 ;
        RECT 1739.880 1545.940 1740.020 1546.360 ;
        RECT 1739.790 1545.680 1740.110 1545.940 ;
        RECT 1739.790 1545.200 1740.110 1545.260 ;
        RECT 1739.595 1545.060 1740.110 1545.200 ;
        RECT 1739.790 1545.000 1740.110 1545.060 ;
        RECT 1739.790 1497.940 1740.110 1498.000 ;
        RECT 1739.595 1497.800 1740.110 1497.940 ;
        RECT 1739.790 1497.740 1740.110 1497.800 ;
        RECT 1739.790 1497.260 1740.110 1497.320 ;
        RECT 1740.250 1497.260 1740.570 1497.320 ;
        RECT 1739.790 1497.120 1740.570 1497.260 ;
        RECT 1739.790 1497.060 1740.110 1497.120 ;
        RECT 1740.250 1497.060 1740.570 1497.120 ;
        RECT 1738.870 1448.980 1739.190 1449.040 ;
        RECT 1739.790 1448.980 1740.110 1449.040 ;
        RECT 1738.870 1448.840 1740.110 1448.980 ;
        RECT 1738.870 1448.780 1739.190 1448.840 ;
        RECT 1739.790 1448.780 1740.110 1448.840 ;
        RECT 1739.790 1400.700 1740.110 1400.760 ;
        RECT 1740.250 1400.700 1740.570 1400.760 ;
        RECT 1739.790 1400.560 1740.570 1400.700 ;
        RECT 1739.790 1400.500 1740.110 1400.560 ;
        RECT 1740.250 1400.500 1740.570 1400.560 ;
        RECT 1739.790 1352.420 1740.110 1352.480 ;
        RECT 1739.595 1352.280 1740.110 1352.420 ;
        RECT 1739.790 1352.220 1740.110 1352.280 ;
        RECT 1739.790 1304.820 1740.110 1304.880 ;
        RECT 1739.595 1304.680 1740.110 1304.820 ;
        RECT 1739.790 1304.620 1740.110 1304.680 ;
        RECT 1739.790 1304.140 1740.110 1304.200 ;
        RECT 1739.790 1304.000 1740.480 1304.140 ;
        RECT 1739.790 1303.940 1740.110 1304.000 ;
        RECT 1740.340 1303.860 1740.480 1304.000 ;
        RECT 1740.250 1303.600 1740.570 1303.860 ;
        RECT 1739.790 1255.860 1740.110 1255.920 ;
        RECT 1739.595 1255.720 1740.110 1255.860 ;
        RECT 1739.790 1255.660 1740.110 1255.720 ;
        RECT 1739.790 1207.580 1740.110 1207.640 ;
        RECT 1739.595 1207.440 1740.110 1207.580 ;
        RECT 1739.790 1207.380 1740.110 1207.440 ;
        RECT 1739.790 1111.020 1740.110 1111.080 ;
        RECT 1740.710 1111.020 1741.030 1111.080 ;
        RECT 1739.790 1110.880 1741.030 1111.020 ;
        RECT 1739.790 1110.820 1740.110 1110.880 ;
        RECT 1740.710 1110.820 1741.030 1110.880 ;
        RECT 1739.790 1014.460 1740.110 1014.520 ;
        RECT 1740.710 1014.460 1741.030 1014.520 ;
        RECT 1739.790 1014.320 1741.030 1014.460 ;
        RECT 1739.790 1014.260 1740.110 1014.320 ;
        RECT 1740.710 1014.260 1741.030 1014.320 ;
        RECT 1739.790 917.900 1740.110 917.960 ;
        RECT 1740.710 917.900 1741.030 917.960 ;
        RECT 1739.790 917.760 1741.030 917.900 ;
        RECT 1739.790 917.700 1740.110 917.760 ;
        RECT 1740.710 917.700 1741.030 917.760 ;
        RECT 1739.790 772.720 1740.110 772.780 ;
        RECT 1740.710 772.720 1741.030 772.780 ;
        RECT 1739.790 772.580 1741.030 772.720 ;
        RECT 1739.790 772.520 1740.110 772.580 ;
        RECT 1740.710 772.520 1741.030 772.580 ;
        RECT 1739.790 676.160 1740.110 676.220 ;
        RECT 1740.710 676.160 1741.030 676.220 ;
        RECT 1739.790 676.020 1741.030 676.160 ;
        RECT 1739.790 675.960 1740.110 676.020 ;
        RECT 1740.710 675.960 1741.030 676.020 ;
        RECT 1739.790 627.880 1740.110 627.940 ;
        RECT 1739.595 627.740 1740.110 627.880 ;
        RECT 1739.790 627.680 1740.110 627.740 ;
        RECT 1739.790 580.280 1740.110 580.340 ;
        RECT 1739.595 580.140 1740.110 580.280 ;
        RECT 1739.790 580.080 1740.110 580.140 ;
        RECT 1739.790 579.600 1740.110 579.660 ;
        RECT 1740.710 579.600 1741.030 579.660 ;
        RECT 1739.790 579.460 1741.030 579.600 ;
        RECT 1739.790 579.400 1740.110 579.460 ;
        RECT 1740.710 579.400 1741.030 579.460 ;
        RECT 1739.790 531.320 1740.110 531.380 ;
        RECT 1739.595 531.180 1740.110 531.320 ;
        RECT 1739.790 531.120 1740.110 531.180 ;
        RECT 1739.790 483.720 1740.110 483.780 ;
        RECT 1739.595 483.580 1740.110 483.720 ;
        RECT 1739.790 483.520 1740.110 483.580 ;
        RECT 1739.790 483.040 1740.110 483.100 ;
        RECT 1740.250 483.040 1740.570 483.100 ;
        RECT 1739.790 482.900 1740.570 483.040 ;
        RECT 1739.790 482.840 1740.110 482.900 ;
        RECT 1740.250 482.840 1740.570 482.900 ;
        RECT 1739.805 372.540 1740.095 372.585 ;
        RECT 1740.250 372.540 1740.570 372.600 ;
        RECT 1739.805 372.400 1740.570 372.540 ;
        RECT 1739.805 372.355 1740.095 372.400 ;
        RECT 1740.250 372.340 1740.570 372.400 ;
        RECT 1739.790 324.600 1740.110 324.660 ;
        RECT 1739.595 324.460 1740.110 324.600 ;
        RECT 1739.790 324.400 1740.110 324.460 ;
        RECT 1739.345 275.980 1739.635 276.025 ;
        RECT 1739.790 275.980 1740.110 276.040 ;
        RECT 1739.345 275.840 1740.110 275.980 ;
        RECT 1739.345 275.795 1739.635 275.840 ;
        RECT 1739.790 275.780 1740.110 275.840 ;
        RECT 1739.345 228.380 1739.635 228.425 ;
        RECT 1739.790 228.380 1740.110 228.440 ;
        RECT 1739.345 228.240 1740.110 228.380 ;
        RECT 1739.345 228.195 1739.635 228.240 ;
        RECT 1739.790 228.180 1740.110 228.240 ;
        RECT 1740.250 34.580 1740.570 34.640 ;
        RECT 1741.170 34.580 1741.490 34.640 ;
        RECT 1740.250 34.440 1741.490 34.580 ;
        RECT 1740.250 34.380 1740.570 34.440 ;
        RECT 1741.170 34.380 1741.490 34.440 ;
        RECT 1572.810 17.240 1573.130 17.300 ;
        RECT 1656.085 17.240 1656.375 17.285 ;
        RECT 1572.810 17.100 1656.375 17.240 ;
        RECT 1572.810 17.040 1573.130 17.100 ;
        RECT 1656.085 17.055 1656.375 17.100 ;
        RECT 1657.005 17.240 1657.295 17.285 ;
        RECT 1740.250 17.240 1740.570 17.300 ;
        RECT 1657.005 17.100 1740.570 17.240 ;
        RECT 1657.005 17.055 1657.295 17.100 ;
        RECT 1740.250 17.040 1740.570 17.100 ;
      LAYER via ;
        RECT 1741.200 1690.180 1741.460 1690.440 ;
        RECT 1739.820 1642.240 1740.080 1642.500 ;
        RECT 1739.820 1641.560 1740.080 1641.820 ;
        RECT 1739.820 1593.960 1740.080 1594.220 ;
        RECT 1739.820 1546.360 1740.080 1546.620 ;
        RECT 1739.820 1545.680 1740.080 1545.940 ;
        RECT 1739.820 1545.000 1740.080 1545.260 ;
        RECT 1739.820 1497.740 1740.080 1498.000 ;
        RECT 1739.820 1497.060 1740.080 1497.320 ;
        RECT 1740.280 1497.060 1740.540 1497.320 ;
        RECT 1738.900 1448.780 1739.160 1449.040 ;
        RECT 1739.820 1448.780 1740.080 1449.040 ;
        RECT 1739.820 1400.500 1740.080 1400.760 ;
        RECT 1740.280 1400.500 1740.540 1400.760 ;
        RECT 1739.820 1352.220 1740.080 1352.480 ;
        RECT 1739.820 1304.620 1740.080 1304.880 ;
        RECT 1739.820 1303.940 1740.080 1304.200 ;
        RECT 1740.280 1303.600 1740.540 1303.860 ;
        RECT 1739.820 1255.660 1740.080 1255.920 ;
        RECT 1739.820 1207.380 1740.080 1207.640 ;
        RECT 1739.820 1110.820 1740.080 1111.080 ;
        RECT 1740.740 1110.820 1741.000 1111.080 ;
        RECT 1739.820 1014.260 1740.080 1014.520 ;
        RECT 1740.740 1014.260 1741.000 1014.520 ;
        RECT 1739.820 917.700 1740.080 917.960 ;
        RECT 1740.740 917.700 1741.000 917.960 ;
        RECT 1739.820 772.520 1740.080 772.780 ;
        RECT 1740.740 772.520 1741.000 772.780 ;
        RECT 1739.820 675.960 1740.080 676.220 ;
        RECT 1740.740 675.960 1741.000 676.220 ;
        RECT 1739.820 627.680 1740.080 627.940 ;
        RECT 1739.820 580.080 1740.080 580.340 ;
        RECT 1739.820 579.400 1740.080 579.660 ;
        RECT 1740.740 579.400 1741.000 579.660 ;
        RECT 1739.820 531.120 1740.080 531.380 ;
        RECT 1739.820 483.520 1740.080 483.780 ;
        RECT 1739.820 482.840 1740.080 483.100 ;
        RECT 1740.280 482.840 1740.540 483.100 ;
        RECT 1740.280 372.340 1740.540 372.600 ;
        RECT 1739.820 324.400 1740.080 324.660 ;
        RECT 1739.820 275.780 1740.080 276.040 ;
        RECT 1739.820 228.180 1740.080 228.440 ;
        RECT 1740.280 34.380 1740.540 34.640 ;
        RECT 1741.200 34.380 1741.460 34.640 ;
        RECT 1572.840 17.040 1573.100 17.300 ;
        RECT 1740.280 17.040 1740.540 17.300 ;
      LAYER met2 ;
        RECT 1742.505 1700.410 1742.785 1704.000 ;
        RECT 1741.260 1700.270 1742.785 1700.410 ;
        RECT 1741.260 1690.470 1741.400 1700.270 ;
        RECT 1742.505 1700.000 1742.785 1700.270 ;
        RECT 1741.200 1690.150 1741.460 1690.470 ;
        RECT 1739.820 1642.210 1740.080 1642.530 ;
        RECT 1739.880 1641.850 1740.020 1642.210 ;
        RECT 1739.820 1641.530 1740.080 1641.850 ;
        RECT 1739.820 1593.930 1740.080 1594.250 ;
        RECT 1739.880 1546.650 1740.020 1593.930 ;
        RECT 1739.820 1546.330 1740.080 1546.650 ;
        RECT 1739.820 1545.650 1740.080 1545.970 ;
        RECT 1739.880 1545.290 1740.020 1545.650 ;
        RECT 1739.820 1544.970 1740.080 1545.290 ;
        RECT 1739.820 1497.710 1740.080 1498.030 ;
        RECT 1739.880 1497.350 1740.020 1497.710 ;
        RECT 1739.820 1497.030 1740.080 1497.350 ;
        RECT 1740.280 1497.030 1740.540 1497.350 ;
        RECT 1740.340 1449.490 1740.480 1497.030 ;
        RECT 1739.880 1449.350 1740.480 1449.490 ;
        RECT 1739.880 1449.070 1740.020 1449.350 ;
        RECT 1738.900 1448.750 1739.160 1449.070 ;
        RECT 1739.820 1448.750 1740.080 1449.070 ;
        RECT 1738.960 1401.325 1739.100 1448.750 ;
        RECT 1738.890 1400.955 1739.170 1401.325 ;
        RECT 1739.810 1400.955 1740.090 1401.325 ;
        RECT 1739.880 1400.790 1740.020 1400.955 ;
        RECT 1739.820 1400.470 1740.080 1400.790 ;
        RECT 1740.280 1400.470 1740.540 1400.790 ;
        RECT 1740.340 1352.930 1740.480 1400.470 ;
        RECT 1739.880 1352.790 1740.480 1352.930 ;
        RECT 1739.880 1352.510 1740.020 1352.790 ;
        RECT 1739.820 1352.190 1740.080 1352.510 ;
        RECT 1739.820 1304.590 1740.080 1304.910 ;
        RECT 1739.880 1304.230 1740.020 1304.590 ;
        RECT 1739.820 1303.910 1740.080 1304.230 ;
        RECT 1740.280 1303.570 1740.540 1303.890 ;
        RECT 1740.340 1256.370 1740.480 1303.570 ;
        RECT 1739.880 1256.230 1740.480 1256.370 ;
        RECT 1739.880 1255.950 1740.020 1256.230 ;
        RECT 1739.820 1255.630 1740.080 1255.950 ;
        RECT 1739.820 1207.350 1740.080 1207.670 ;
        RECT 1739.880 1159.245 1740.020 1207.350 ;
        RECT 1739.810 1158.875 1740.090 1159.245 ;
        RECT 1740.730 1158.875 1741.010 1159.245 ;
        RECT 1740.800 1111.110 1740.940 1158.875 ;
        RECT 1739.820 1110.790 1740.080 1111.110 ;
        RECT 1740.740 1110.790 1741.000 1111.110 ;
        RECT 1739.880 1062.685 1740.020 1110.790 ;
        RECT 1739.810 1062.315 1740.090 1062.685 ;
        RECT 1740.730 1062.315 1741.010 1062.685 ;
        RECT 1740.800 1014.550 1740.940 1062.315 ;
        RECT 1739.820 1014.230 1740.080 1014.550 ;
        RECT 1740.740 1014.230 1741.000 1014.550 ;
        RECT 1739.880 966.125 1740.020 1014.230 ;
        RECT 1739.810 965.755 1740.090 966.125 ;
        RECT 1740.730 965.755 1741.010 966.125 ;
        RECT 1740.800 917.990 1740.940 965.755 ;
        RECT 1739.820 917.670 1740.080 917.990 ;
        RECT 1740.740 917.670 1741.000 917.990 ;
        RECT 1739.880 869.565 1740.020 917.670 ;
        RECT 1739.810 869.195 1740.090 869.565 ;
        RECT 1740.730 869.195 1741.010 869.565 ;
        RECT 1740.800 821.285 1740.940 869.195 ;
        RECT 1739.810 820.915 1740.090 821.285 ;
        RECT 1740.730 820.915 1741.010 821.285 ;
        RECT 1739.880 772.810 1740.020 820.915 ;
        RECT 1739.820 772.490 1740.080 772.810 ;
        RECT 1740.740 772.490 1741.000 772.810 ;
        RECT 1740.800 724.725 1740.940 772.490 ;
        RECT 1739.810 724.355 1740.090 724.725 ;
        RECT 1740.730 724.355 1741.010 724.725 ;
        RECT 1739.880 676.250 1740.020 724.355 ;
        RECT 1739.820 675.930 1740.080 676.250 ;
        RECT 1740.740 675.930 1741.000 676.250 ;
        RECT 1740.800 628.165 1740.940 675.930 ;
        RECT 1739.810 627.795 1740.090 628.165 ;
        RECT 1740.730 627.795 1741.010 628.165 ;
        RECT 1739.820 627.650 1740.080 627.795 ;
        RECT 1739.820 580.050 1740.080 580.370 ;
        RECT 1739.880 579.690 1740.020 580.050 ;
        RECT 1739.820 579.370 1740.080 579.690 ;
        RECT 1740.740 579.370 1741.000 579.690 ;
        RECT 1740.800 531.605 1740.940 579.370 ;
        RECT 1739.810 531.235 1740.090 531.605 ;
        RECT 1740.730 531.235 1741.010 531.605 ;
        RECT 1739.820 531.090 1740.080 531.235 ;
        RECT 1739.820 483.490 1740.080 483.810 ;
        RECT 1739.880 483.130 1740.020 483.490 ;
        RECT 1739.820 482.810 1740.080 483.130 ;
        RECT 1740.280 482.810 1740.540 483.130 ;
        RECT 1740.340 448.530 1740.480 482.810 ;
        RECT 1739.880 448.390 1740.480 448.530 ;
        RECT 1739.880 434.930 1740.020 448.390 ;
        RECT 1739.880 434.790 1740.480 434.930 ;
        RECT 1740.340 400.930 1740.480 434.790 ;
        RECT 1740.340 400.790 1740.940 400.930 ;
        RECT 1740.800 373.050 1740.940 400.790 ;
        RECT 1740.340 372.910 1740.940 373.050 ;
        RECT 1740.340 372.630 1740.480 372.910 ;
        RECT 1740.280 372.310 1740.540 372.630 ;
        RECT 1739.820 324.370 1740.080 324.690 ;
        RECT 1739.880 276.070 1740.020 324.370 ;
        RECT 1739.820 275.750 1740.080 276.070 ;
        RECT 1739.820 228.150 1740.080 228.470 ;
        RECT 1739.880 227.645 1740.020 228.150 ;
        RECT 1739.810 227.275 1740.090 227.645 ;
        RECT 1740.270 226.595 1740.550 226.965 ;
        RECT 1740.340 131.085 1740.480 226.595 ;
        RECT 1740.270 130.715 1740.550 131.085 ;
        RECT 1741.190 130.715 1741.470 131.085 ;
        RECT 1741.260 124.285 1741.400 130.715 ;
        RECT 1740.270 123.915 1740.550 124.285 ;
        RECT 1741.190 123.915 1741.470 124.285 ;
        RECT 1740.340 81.330 1740.480 123.915 ;
        RECT 1740.340 81.190 1741.400 81.330 ;
        RECT 1741.260 34.670 1741.400 81.190 ;
        RECT 1740.280 34.350 1740.540 34.670 ;
        RECT 1741.200 34.350 1741.460 34.670 ;
        RECT 1740.340 17.330 1740.480 34.350 ;
        RECT 1572.840 17.010 1573.100 17.330 ;
        RECT 1740.280 17.010 1740.540 17.330 ;
        RECT 1572.900 2.400 1573.040 17.010 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 1738.890 1401.000 1739.170 1401.280 ;
        RECT 1739.810 1401.000 1740.090 1401.280 ;
        RECT 1739.810 1158.920 1740.090 1159.200 ;
        RECT 1740.730 1158.920 1741.010 1159.200 ;
        RECT 1739.810 1062.360 1740.090 1062.640 ;
        RECT 1740.730 1062.360 1741.010 1062.640 ;
        RECT 1739.810 965.800 1740.090 966.080 ;
        RECT 1740.730 965.800 1741.010 966.080 ;
        RECT 1739.810 869.240 1740.090 869.520 ;
        RECT 1740.730 869.240 1741.010 869.520 ;
        RECT 1739.810 820.960 1740.090 821.240 ;
        RECT 1740.730 820.960 1741.010 821.240 ;
        RECT 1739.810 724.400 1740.090 724.680 ;
        RECT 1740.730 724.400 1741.010 724.680 ;
        RECT 1739.810 627.840 1740.090 628.120 ;
        RECT 1740.730 627.840 1741.010 628.120 ;
        RECT 1739.810 531.280 1740.090 531.560 ;
        RECT 1740.730 531.280 1741.010 531.560 ;
        RECT 1739.810 227.320 1740.090 227.600 ;
        RECT 1740.270 226.640 1740.550 226.920 ;
        RECT 1740.270 130.760 1740.550 131.040 ;
        RECT 1741.190 130.760 1741.470 131.040 ;
        RECT 1740.270 123.960 1740.550 124.240 ;
        RECT 1741.190 123.960 1741.470 124.240 ;
      LAYER met3 ;
        RECT 1738.865 1401.290 1739.195 1401.305 ;
        RECT 1739.785 1401.290 1740.115 1401.305 ;
        RECT 1738.865 1400.990 1740.115 1401.290 ;
        RECT 1738.865 1400.975 1739.195 1400.990 ;
        RECT 1739.785 1400.975 1740.115 1400.990 ;
        RECT 1739.785 1159.210 1740.115 1159.225 ;
        RECT 1740.705 1159.210 1741.035 1159.225 ;
        RECT 1739.785 1158.910 1741.035 1159.210 ;
        RECT 1739.785 1158.895 1740.115 1158.910 ;
        RECT 1740.705 1158.895 1741.035 1158.910 ;
        RECT 1739.785 1062.650 1740.115 1062.665 ;
        RECT 1740.705 1062.650 1741.035 1062.665 ;
        RECT 1739.785 1062.350 1741.035 1062.650 ;
        RECT 1739.785 1062.335 1740.115 1062.350 ;
        RECT 1740.705 1062.335 1741.035 1062.350 ;
        RECT 1739.785 966.090 1740.115 966.105 ;
        RECT 1740.705 966.090 1741.035 966.105 ;
        RECT 1739.785 965.790 1741.035 966.090 ;
        RECT 1739.785 965.775 1740.115 965.790 ;
        RECT 1740.705 965.775 1741.035 965.790 ;
        RECT 1739.785 869.530 1740.115 869.545 ;
        RECT 1740.705 869.530 1741.035 869.545 ;
        RECT 1739.785 869.230 1741.035 869.530 ;
        RECT 1739.785 869.215 1740.115 869.230 ;
        RECT 1740.705 869.215 1741.035 869.230 ;
        RECT 1739.785 821.250 1740.115 821.265 ;
        RECT 1740.705 821.250 1741.035 821.265 ;
        RECT 1739.785 820.950 1741.035 821.250 ;
        RECT 1739.785 820.935 1740.115 820.950 ;
        RECT 1740.705 820.935 1741.035 820.950 ;
        RECT 1739.785 724.690 1740.115 724.705 ;
        RECT 1740.705 724.690 1741.035 724.705 ;
        RECT 1739.785 724.390 1741.035 724.690 ;
        RECT 1739.785 724.375 1740.115 724.390 ;
        RECT 1740.705 724.375 1741.035 724.390 ;
        RECT 1739.785 628.130 1740.115 628.145 ;
        RECT 1740.705 628.130 1741.035 628.145 ;
        RECT 1739.785 627.830 1741.035 628.130 ;
        RECT 1739.785 627.815 1740.115 627.830 ;
        RECT 1740.705 627.815 1741.035 627.830 ;
        RECT 1739.785 531.570 1740.115 531.585 ;
        RECT 1740.705 531.570 1741.035 531.585 ;
        RECT 1739.785 531.270 1741.035 531.570 ;
        RECT 1739.785 531.255 1740.115 531.270 ;
        RECT 1740.705 531.255 1741.035 531.270 ;
        RECT 1739.785 227.610 1740.115 227.625 ;
        RECT 1739.110 227.310 1740.115 227.610 ;
        RECT 1739.110 226.930 1739.410 227.310 ;
        RECT 1739.785 227.295 1740.115 227.310 ;
        RECT 1740.245 226.930 1740.575 226.945 ;
        RECT 1739.110 226.630 1740.575 226.930 ;
        RECT 1740.245 226.615 1740.575 226.630 ;
        RECT 1740.245 131.050 1740.575 131.065 ;
        RECT 1741.165 131.050 1741.495 131.065 ;
        RECT 1740.245 130.750 1741.495 131.050 ;
        RECT 1740.245 130.735 1740.575 130.750 ;
        RECT 1741.165 130.735 1741.495 130.750 ;
        RECT 1740.245 124.250 1740.575 124.265 ;
        RECT 1741.165 124.250 1741.495 124.265 ;
        RECT 1740.245 123.950 1741.495 124.250 ;
        RECT 1740.245 123.935 1740.575 123.950 ;
        RECT 1741.165 123.935 1741.495 123.950 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1708.585 1684.785 1708.755 1689.375 ;
        RECT 1633.145 14.195 1633.315 14.535 ;
        RECT 1631.765 14.025 1633.315 14.195 ;
      LAYER mcon ;
        RECT 1708.585 1689.205 1708.755 1689.375 ;
        RECT 1633.145 14.365 1633.315 14.535 ;
      LAYER met1 ;
        RECT 1708.525 1689.360 1708.815 1689.405 ;
        RECT 1747.150 1689.360 1747.470 1689.420 ;
        RECT 1708.525 1689.220 1747.470 1689.360 ;
        RECT 1708.525 1689.175 1708.815 1689.220 ;
        RECT 1747.150 1689.160 1747.470 1689.220 ;
        RECT 1638.590 1684.940 1638.910 1685.000 ;
        RECT 1708.525 1684.940 1708.815 1684.985 ;
        RECT 1638.590 1684.800 1708.815 1684.940 ;
        RECT 1638.590 1684.740 1638.910 1684.800 ;
        RECT 1708.525 1684.755 1708.815 1684.800 ;
        RECT 1633.085 14.520 1633.375 14.565 ;
        RECT 1638.590 14.520 1638.910 14.580 ;
        RECT 1633.085 14.380 1638.910 14.520 ;
        RECT 1633.085 14.335 1633.375 14.380 ;
        RECT 1638.590 14.320 1638.910 14.380 ;
        RECT 1590.290 14.180 1590.610 14.240 ;
        RECT 1631.705 14.180 1631.995 14.225 ;
        RECT 1590.290 14.040 1631.995 14.180 ;
        RECT 1590.290 13.980 1590.610 14.040 ;
        RECT 1631.705 13.995 1631.995 14.040 ;
      LAYER via ;
        RECT 1747.180 1689.160 1747.440 1689.420 ;
        RECT 1638.620 1684.740 1638.880 1685.000 ;
        RECT 1638.620 14.320 1638.880 14.580 ;
        RECT 1590.320 13.980 1590.580 14.240 ;
      LAYER met2 ;
        RECT 1748.945 1700.410 1749.225 1704.000 ;
        RECT 1747.240 1700.270 1749.225 1700.410 ;
        RECT 1747.240 1689.450 1747.380 1700.270 ;
        RECT 1748.945 1700.000 1749.225 1700.270 ;
        RECT 1747.180 1689.130 1747.440 1689.450 ;
        RECT 1638.620 1684.710 1638.880 1685.030 ;
        RECT 1638.680 14.610 1638.820 1684.710 ;
        RECT 1638.620 14.290 1638.880 14.610 ;
        RECT 1590.320 13.950 1590.580 14.270 ;
        RECT 1590.380 2.400 1590.520 13.950 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1652.925 17.425 1653.095 18.955 ;
      LAYER mcon ;
        RECT 1652.925 18.785 1653.095 18.955 ;
      LAYER met1 ;
        RECT 1652.865 18.940 1653.155 18.985 ;
        RECT 1754.050 18.940 1754.370 19.000 ;
        RECT 1652.865 18.800 1754.370 18.940 ;
        RECT 1652.865 18.755 1653.155 18.800 ;
        RECT 1754.050 18.740 1754.370 18.800 ;
        RECT 1632.150 17.580 1632.470 17.640 ;
        RECT 1652.865 17.580 1653.155 17.625 ;
        RECT 1632.150 17.440 1653.155 17.580 ;
        RECT 1632.150 17.380 1632.470 17.440 ;
        RECT 1652.865 17.395 1653.155 17.440 ;
        RECT 1608.230 16.900 1608.550 16.960 ;
        RECT 1631.230 16.900 1631.550 16.960 ;
        RECT 1608.230 16.760 1631.550 16.900 ;
        RECT 1608.230 16.700 1608.550 16.760 ;
        RECT 1631.230 16.700 1631.550 16.760 ;
      LAYER via ;
        RECT 1754.080 18.740 1754.340 19.000 ;
        RECT 1632.180 17.380 1632.440 17.640 ;
        RECT 1608.260 16.700 1608.520 16.960 ;
        RECT 1631.260 16.700 1631.520 16.960 ;
      LAYER met2 ;
        RECT 1755.845 1700.410 1756.125 1704.000 ;
        RECT 1754.140 1700.270 1756.125 1700.410 ;
        RECT 1754.140 19.030 1754.280 1700.270 ;
        RECT 1755.845 1700.000 1756.125 1700.270 ;
        RECT 1754.080 18.710 1754.340 19.030 ;
        RECT 1632.180 17.410 1632.440 17.670 ;
        RECT 1631.320 17.350 1632.440 17.410 ;
        RECT 1631.320 17.270 1632.380 17.350 ;
        RECT 1631.320 16.990 1631.460 17.270 ;
        RECT 1608.260 16.670 1608.520 16.990 ;
        RECT 1631.260 16.670 1631.520 16.990 ;
        RECT 1608.320 2.400 1608.460 16.670 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1728.365 1686.825 1728.535 1688.695 ;
      LAYER mcon ;
        RECT 1728.365 1688.525 1728.535 1688.695 ;
      LAYER met1 ;
        RECT 1728.305 1688.680 1728.595 1688.725 ;
        RECT 1700.780 1688.540 1728.595 1688.680 ;
        RECT 1652.390 1688.000 1652.710 1688.060 ;
        RECT 1700.780 1688.000 1700.920 1688.540 ;
        RECT 1728.305 1688.495 1728.595 1688.540 ;
        RECT 1652.390 1687.860 1700.920 1688.000 ;
        RECT 1652.390 1687.800 1652.710 1687.860 ;
        RECT 1728.305 1686.980 1728.595 1687.025 ;
        RECT 1760.950 1686.980 1761.270 1687.040 ;
        RECT 1728.305 1686.840 1761.270 1686.980 ;
        RECT 1728.305 1686.795 1728.595 1686.840 ;
        RECT 1760.950 1686.780 1761.270 1686.840 ;
        RECT 1626.170 18.940 1626.490 19.000 ;
        RECT 1652.390 18.940 1652.710 19.000 ;
        RECT 1626.170 18.800 1652.710 18.940 ;
        RECT 1626.170 18.740 1626.490 18.800 ;
        RECT 1652.390 18.740 1652.710 18.800 ;
      LAYER via ;
        RECT 1652.420 1687.800 1652.680 1688.060 ;
        RECT 1760.980 1686.780 1761.240 1687.040 ;
        RECT 1626.200 18.740 1626.460 19.000 ;
        RECT 1652.420 18.740 1652.680 19.000 ;
      LAYER met2 ;
        RECT 1762.745 1700.410 1763.025 1704.000 ;
        RECT 1761.040 1700.270 1763.025 1700.410 ;
        RECT 1652.420 1687.770 1652.680 1688.090 ;
        RECT 1652.480 19.030 1652.620 1687.770 ;
        RECT 1761.040 1687.070 1761.180 1700.270 ;
        RECT 1762.745 1700.000 1763.025 1700.270 ;
        RECT 1760.980 1686.750 1761.240 1687.070 ;
        RECT 1626.200 18.710 1626.460 19.030 ;
        RECT 1652.420 18.710 1652.680 19.030 ;
        RECT 1626.260 2.400 1626.400 18.710 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1727.905 1685.125 1728.075 1687.675 ;
      LAYER mcon ;
        RECT 1727.905 1687.505 1728.075 1687.675 ;
      LAYER met1 ;
        RECT 1673.090 1687.660 1673.410 1687.720 ;
        RECT 1727.845 1687.660 1728.135 1687.705 ;
        RECT 1673.090 1687.520 1728.135 1687.660 ;
        RECT 1673.090 1687.460 1673.410 1687.520 ;
        RECT 1727.845 1687.475 1728.135 1687.520 ;
        RECT 1727.845 1685.280 1728.135 1685.325 ;
        RECT 1769.230 1685.280 1769.550 1685.340 ;
        RECT 1727.845 1685.140 1769.550 1685.280 ;
        RECT 1727.845 1685.095 1728.135 1685.140 ;
        RECT 1769.230 1685.080 1769.550 1685.140 ;
        RECT 1644.110 18.600 1644.430 18.660 ;
        RECT 1673.090 18.600 1673.410 18.660 ;
        RECT 1644.110 18.460 1673.410 18.600 ;
        RECT 1644.110 18.400 1644.430 18.460 ;
        RECT 1673.090 18.400 1673.410 18.460 ;
      LAYER via ;
        RECT 1673.120 1687.460 1673.380 1687.720 ;
        RECT 1769.260 1685.080 1769.520 1685.340 ;
        RECT 1644.140 18.400 1644.400 18.660 ;
        RECT 1673.120 18.400 1673.380 18.660 ;
      LAYER met2 ;
        RECT 1769.185 1700.000 1769.465 1704.000 ;
        RECT 1673.120 1687.430 1673.380 1687.750 ;
        RECT 1673.180 18.690 1673.320 1687.430 ;
        RECT 1769.320 1685.370 1769.460 1700.000 ;
        RECT 1769.260 1685.050 1769.520 1685.370 ;
        RECT 1644.140 18.370 1644.400 18.690 ;
        RECT 1673.120 18.370 1673.380 18.690 ;
        RECT 1644.200 2.400 1644.340 18.370 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.050 16.900 1662.370 16.960 ;
        RECT 1774.290 16.900 1774.610 16.960 ;
        RECT 1662.050 16.760 1774.610 16.900 ;
        RECT 1662.050 16.700 1662.370 16.760 ;
        RECT 1774.290 16.700 1774.610 16.760 ;
      LAYER via ;
        RECT 1662.080 16.700 1662.340 16.960 ;
        RECT 1774.320 16.700 1774.580 16.960 ;
      LAYER met2 ;
        RECT 1776.085 1700.410 1776.365 1704.000 ;
        RECT 1774.380 1700.270 1776.365 1700.410 ;
        RECT 1774.380 16.990 1774.520 1700.270 ;
        RECT 1776.085 1700.000 1776.365 1700.270 ;
        RECT 1662.080 16.670 1662.340 16.990 ;
        RECT 1774.320 16.670 1774.580 16.990 ;
        RECT 1662.140 2.400 1662.280 16.670 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1679.530 14.180 1679.850 14.240 ;
        RECT 1782.570 14.180 1782.890 14.240 ;
        RECT 1679.530 14.040 1782.890 14.180 ;
        RECT 1679.530 13.980 1679.850 14.040 ;
        RECT 1782.570 13.980 1782.890 14.040 ;
      LAYER via ;
        RECT 1679.560 13.980 1679.820 14.240 ;
        RECT 1782.600 13.980 1782.860 14.240 ;
      LAYER met2 ;
        RECT 1782.985 1700.410 1783.265 1704.000 ;
        RECT 1782.660 1700.270 1783.265 1700.410 ;
        RECT 1782.660 14.270 1782.800 1700.270 ;
        RECT 1782.985 1700.000 1783.265 1700.270 ;
        RECT 1679.560 13.950 1679.820 14.270 ;
        RECT 1782.600 13.950 1782.860 14.270 ;
        RECT 1679.620 2.400 1679.760 13.950 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.470 18.600 1697.790 18.660 ;
        RECT 1788.090 18.600 1788.410 18.660 ;
        RECT 1697.470 18.460 1788.410 18.600 ;
        RECT 1697.470 18.400 1697.790 18.460 ;
        RECT 1788.090 18.400 1788.410 18.460 ;
      LAYER via ;
        RECT 1697.500 18.400 1697.760 18.660 ;
        RECT 1788.120 18.400 1788.380 18.660 ;
      LAYER met2 ;
        RECT 1789.425 1700.410 1789.705 1704.000 ;
        RECT 1788.180 1700.270 1789.705 1700.410 ;
        RECT 1788.180 18.690 1788.320 1700.270 ;
        RECT 1789.425 1700.000 1789.705 1700.270 ;
        RECT 1697.500 18.370 1697.760 18.690 ;
        RECT 1788.120 18.370 1788.380 18.690 ;
        RECT 1697.560 2.400 1697.700 18.370 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.930 1665.900 1422.250 1665.960 ;
        RECT 1424.230 1665.900 1424.550 1665.960 ;
        RECT 1421.930 1665.760 1424.550 1665.900 ;
        RECT 1421.930 1665.700 1422.250 1665.760 ;
        RECT 1424.230 1665.700 1424.550 1665.760 ;
        RECT 734.230 47.160 734.550 47.220 ;
        RECT 1421.930 47.160 1422.250 47.220 ;
        RECT 734.230 47.020 1422.250 47.160 ;
        RECT 734.230 46.960 734.550 47.020 ;
        RECT 1421.930 46.960 1422.250 47.020 ;
      LAYER via ;
        RECT 1421.960 1665.700 1422.220 1665.960 ;
        RECT 1424.260 1665.700 1424.520 1665.960 ;
        RECT 734.260 46.960 734.520 47.220 ;
        RECT 1421.960 46.960 1422.220 47.220 ;
      LAYER met2 ;
        RECT 1426.025 1700.410 1426.305 1704.000 ;
        RECT 1424.320 1700.270 1426.305 1700.410 ;
        RECT 1424.320 1665.990 1424.460 1700.270 ;
        RECT 1426.025 1700.000 1426.305 1700.270 ;
        RECT 1421.960 1665.670 1422.220 1665.990 ;
        RECT 1424.260 1665.670 1424.520 1665.990 ;
        RECT 1422.020 47.250 1422.160 1665.670 ;
        RECT 734.260 46.930 734.520 47.250 ;
        RECT 1421.960 46.930 1422.220 47.250 ;
        RECT 734.320 2.400 734.460 46.930 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1749.525 19.125 1749.695 20.655 ;
      LAYER mcon ;
        RECT 1749.525 20.485 1749.695 20.655 ;
      LAYER met1 ;
        RECT 1776.590 1689.360 1776.910 1689.420 ;
        RECT 1796.370 1689.360 1796.690 1689.420 ;
        RECT 1776.590 1689.220 1796.690 1689.360 ;
        RECT 1776.590 1689.160 1776.910 1689.220 ;
        RECT 1796.370 1689.160 1796.690 1689.220 ;
        RECT 1749.465 20.640 1749.755 20.685 ;
        RECT 1776.590 20.640 1776.910 20.700 ;
        RECT 1749.465 20.500 1776.910 20.640 ;
        RECT 1749.465 20.455 1749.755 20.500 ;
        RECT 1776.590 20.440 1776.910 20.500 ;
        RECT 1715.410 19.620 1715.730 19.680 ;
        RECT 1715.410 19.480 1721.620 19.620 ;
        RECT 1715.410 19.420 1715.730 19.480 ;
        RECT 1721.480 19.280 1721.620 19.480 ;
        RECT 1749.465 19.280 1749.755 19.325 ;
        RECT 1721.480 19.140 1749.755 19.280 ;
        RECT 1749.465 19.095 1749.755 19.140 ;
      LAYER via ;
        RECT 1776.620 1689.160 1776.880 1689.420 ;
        RECT 1796.400 1689.160 1796.660 1689.420 ;
        RECT 1776.620 20.440 1776.880 20.700 ;
        RECT 1715.440 19.420 1715.700 19.680 ;
      LAYER met2 ;
        RECT 1796.325 1700.000 1796.605 1704.000 ;
        RECT 1796.460 1689.450 1796.600 1700.000 ;
        RECT 1776.620 1689.130 1776.880 1689.450 ;
        RECT 1796.400 1689.130 1796.660 1689.450 ;
        RECT 1776.680 20.730 1776.820 1689.130 ;
        RECT 1776.620 20.410 1776.880 20.730 ;
        RECT 1715.440 19.390 1715.700 19.710 ;
        RECT 1715.500 2.400 1715.640 19.390 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1783.490 1688.680 1783.810 1688.740 ;
        RECT 1802.810 1688.680 1803.130 1688.740 ;
        RECT 1783.490 1688.540 1803.130 1688.680 ;
        RECT 1783.490 1688.480 1783.810 1688.540 ;
        RECT 1802.810 1688.480 1803.130 1688.540 ;
        RECT 1733.350 20.300 1733.670 20.360 ;
        RECT 1783.490 20.300 1783.810 20.360 ;
        RECT 1733.350 20.160 1783.810 20.300 ;
        RECT 1733.350 20.100 1733.670 20.160 ;
        RECT 1783.490 20.100 1783.810 20.160 ;
      LAYER via ;
        RECT 1783.520 1688.480 1783.780 1688.740 ;
        RECT 1802.840 1688.480 1803.100 1688.740 ;
        RECT 1733.380 20.100 1733.640 20.360 ;
        RECT 1783.520 20.100 1783.780 20.360 ;
      LAYER met2 ;
        RECT 1802.765 1700.000 1803.045 1704.000 ;
        RECT 1802.900 1688.770 1803.040 1700.000 ;
        RECT 1783.520 1688.450 1783.780 1688.770 ;
        RECT 1802.840 1688.450 1803.100 1688.770 ;
        RECT 1783.580 20.390 1783.720 1688.450 ;
        RECT 1733.380 20.070 1733.640 20.390 ;
        RECT 1783.520 20.070 1783.780 20.390 ;
        RECT 1733.440 2.400 1733.580 20.070 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1808.790 17.580 1809.110 17.640 ;
        RECT 1790.940 17.440 1809.110 17.580 ;
        RECT 1751.290 17.240 1751.610 17.300 ;
        RECT 1790.940 17.240 1791.080 17.440 ;
        RECT 1808.790 17.380 1809.110 17.440 ;
        RECT 1751.290 17.100 1791.080 17.240 ;
        RECT 1751.290 17.040 1751.610 17.100 ;
      LAYER via ;
        RECT 1751.320 17.040 1751.580 17.300 ;
        RECT 1808.820 17.380 1809.080 17.640 ;
      LAYER met2 ;
        RECT 1809.665 1700.410 1809.945 1704.000 ;
        RECT 1808.880 1700.270 1809.945 1700.410 ;
        RECT 1808.880 17.670 1809.020 1700.270 ;
        RECT 1809.665 1700.000 1809.945 1700.270 ;
        RECT 1808.820 17.350 1809.080 17.670 ;
        RECT 1751.320 17.010 1751.580 17.330 ;
        RECT 1751.380 2.400 1751.520 17.010 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1790.390 1688.000 1790.710 1688.060 ;
        RECT 1816.610 1688.000 1816.930 1688.060 ;
        RECT 1790.390 1687.860 1816.930 1688.000 ;
        RECT 1790.390 1687.800 1790.710 1687.860 ;
        RECT 1816.610 1687.800 1816.930 1687.860 ;
        RECT 1768.770 17.920 1769.090 17.980 ;
        RECT 1790.390 17.920 1790.710 17.980 ;
        RECT 1768.770 17.780 1790.710 17.920 ;
        RECT 1768.770 17.720 1769.090 17.780 ;
        RECT 1790.390 17.720 1790.710 17.780 ;
      LAYER via ;
        RECT 1790.420 1687.800 1790.680 1688.060 ;
        RECT 1816.640 1687.800 1816.900 1688.060 ;
        RECT 1768.800 17.720 1769.060 17.980 ;
        RECT 1790.420 17.720 1790.680 17.980 ;
      LAYER met2 ;
        RECT 1816.565 1700.000 1816.845 1704.000 ;
        RECT 1816.700 1688.090 1816.840 1700.000 ;
        RECT 1790.420 1687.770 1790.680 1688.090 ;
        RECT 1816.640 1687.770 1816.900 1688.090 ;
        RECT 1790.480 18.010 1790.620 1687.770 ;
        RECT 1768.800 17.690 1769.060 18.010 ;
        RECT 1790.420 17.690 1790.680 18.010 ;
        RECT 1768.860 2.400 1769.000 17.690 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1797.290 1685.280 1797.610 1685.340 ;
        RECT 1823.050 1685.280 1823.370 1685.340 ;
        RECT 1797.290 1685.140 1823.370 1685.280 ;
        RECT 1797.290 1685.080 1797.610 1685.140 ;
        RECT 1823.050 1685.080 1823.370 1685.140 ;
        RECT 1786.710 15.540 1787.030 15.600 ;
        RECT 1797.290 15.540 1797.610 15.600 ;
        RECT 1786.710 15.400 1797.610 15.540 ;
        RECT 1786.710 15.340 1787.030 15.400 ;
        RECT 1797.290 15.340 1797.610 15.400 ;
      LAYER via ;
        RECT 1797.320 1685.080 1797.580 1685.340 ;
        RECT 1823.080 1685.080 1823.340 1685.340 ;
        RECT 1786.740 15.340 1787.000 15.600 ;
        RECT 1797.320 15.340 1797.580 15.600 ;
      LAYER met2 ;
        RECT 1823.005 1700.000 1823.285 1704.000 ;
        RECT 1823.140 1685.370 1823.280 1700.000 ;
        RECT 1797.320 1685.050 1797.580 1685.370 ;
        RECT 1823.080 1685.050 1823.340 1685.370 ;
        RECT 1797.380 15.630 1797.520 1685.050 ;
        RECT 1786.740 15.310 1787.000 15.630 ;
        RECT 1797.320 15.310 1797.580 15.630 ;
        RECT 1786.800 2.400 1786.940 15.310 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1811.090 1684.260 1811.410 1684.320 ;
        RECT 1829.950 1684.260 1830.270 1684.320 ;
        RECT 1811.090 1684.120 1830.270 1684.260 ;
        RECT 1811.090 1684.060 1811.410 1684.120 ;
        RECT 1829.950 1684.060 1830.270 1684.120 ;
        RECT 1804.650 19.960 1804.970 20.020 ;
        RECT 1811.090 19.960 1811.410 20.020 ;
        RECT 1804.650 19.820 1811.410 19.960 ;
        RECT 1804.650 19.760 1804.970 19.820 ;
        RECT 1811.090 19.760 1811.410 19.820 ;
      LAYER via ;
        RECT 1811.120 1684.060 1811.380 1684.320 ;
        RECT 1829.980 1684.060 1830.240 1684.320 ;
        RECT 1804.680 19.760 1804.940 20.020 ;
        RECT 1811.120 19.760 1811.380 20.020 ;
      LAYER met2 ;
        RECT 1829.905 1700.000 1830.185 1704.000 ;
        RECT 1830.040 1684.350 1830.180 1700.000 ;
        RECT 1811.120 1684.030 1811.380 1684.350 ;
        RECT 1829.980 1684.030 1830.240 1684.350 ;
        RECT 1811.180 20.050 1811.320 1684.030 ;
        RECT 1804.680 19.730 1804.940 20.050 ;
        RECT 1811.120 19.730 1811.380 20.050 ;
        RECT 1804.740 2.400 1804.880 19.730 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1831.790 1684.600 1832.110 1684.660 ;
        RECT 1836.850 1684.600 1837.170 1684.660 ;
        RECT 1831.790 1684.460 1837.170 1684.600 ;
        RECT 1831.790 1684.400 1832.110 1684.460 ;
        RECT 1836.850 1684.400 1837.170 1684.460 ;
        RECT 1822.590 20.640 1822.910 20.700 ;
        RECT 1831.790 20.640 1832.110 20.700 ;
        RECT 1822.590 20.500 1832.110 20.640 ;
        RECT 1822.590 20.440 1822.910 20.500 ;
        RECT 1831.790 20.440 1832.110 20.500 ;
      LAYER via ;
        RECT 1831.820 1684.400 1832.080 1684.660 ;
        RECT 1836.880 1684.400 1837.140 1684.660 ;
        RECT 1822.620 20.440 1822.880 20.700 ;
        RECT 1831.820 20.440 1832.080 20.700 ;
      LAYER met2 ;
        RECT 1836.805 1700.000 1837.085 1704.000 ;
        RECT 1836.940 1684.690 1837.080 1700.000 ;
        RECT 1831.820 1684.370 1832.080 1684.690 ;
        RECT 1836.880 1684.370 1837.140 1684.690 ;
        RECT 1831.880 20.730 1832.020 1684.370 ;
        RECT 1822.620 20.410 1822.880 20.730 ;
        RECT 1831.820 20.410 1832.080 20.730 ;
        RECT 1822.680 2.400 1822.820 20.410 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1840.070 20.640 1840.390 20.700 ;
        RECT 1842.370 20.640 1842.690 20.700 ;
        RECT 1840.070 20.500 1842.690 20.640 ;
        RECT 1840.070 20.440 1840.390 20.500 ;
        RECT 1842.370 20.440 1842.690 20.500 ;
      LAYER via ;
        RECT 1840.100 20.440 1840.360 20.700 ;
        RECT 1842.400 20.440 1842.660 20.700 ;
      LAYER met2 ;
        RECT 1843.245 1700.410 1843.525 1704.000 ;
        RECT 1842.460 1700.270 1843.525 1700.410 ;
        RECT 1842.460 20.730 1842.600 1700.270 ;
        RECT 1843.245 1700.000 1843.525 1700.270 ;
        RECT 1840.100 20.410 1840.360 20.730 ;
        RECT 1842.400 20.410 1842.660 20.730 ;
        RECT 1840.160 2.400 1840.300 20.410 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1850.190 1689.360 1850.510 1689.420 ;
        RECT 1855.250 1689.360 1855.570 1689.420 ;
        RECT 1850.190 1689.220 1855.570 1689.360 ;
        RECT 1850.190 1689.160 1850.510 1689.220 ;
        RECT 1855.250 1689.160 1855.570 1689.220 ;
        RECT 1855.250 17.580 1855.570 17.640 ;
        RECT 1858.010 17.580 1858.330 17.640 ;
        RECT 1855.250 17.440 1858.330 17.580 ;
        RECT 1855.250 17.380 1855.570 17.440 ;
        RECT 1858.010 17.380 1858.330 17.440 ;
      LAYER via ;
        RECT 1850.220 1689.160 1850.480 1689.420 ;
        RECT 1855.280 1689.160 1855.540 1689.420 ;
        RECT 1855.280 17.380 1855.540 17.640 ;
        RECT 1858.040 17.380 1858.300 17.640 ;
      LAYER met2 ;
        RECT 1850.145 1700.000 1850.425 1704.000 ;
        RECT 1850.280 1689.450 1850.420 1700.000 ;
        RECT 1850.220 1689.130 1850.480 1689.450 ;
        RECT 1855.280 1689.130 1855.540 1689.450 ;
        RECT 1855.340 17.670 1855.480 1689.130 ;
        RECT 1855.280 17.350 1855.540 17.670 ;
        RECT 1858.040 17.350 1858.300 17.670 ;
        RECT 1858.100 2.400 1858.240 17.350 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1857.090 1687.660 1857.410 1687.720 ;
        RECT 1870.430 1687.660 1870.750 1687.720 ;
        RECT 1857.090 1687.520 1870.750 1687.660 ;
        RECT 1857.090 1687.460 1857.410 1687.520 ;
        RECT 1870.430 1687.460 1870.750 1687.520 ;
      LAYER via ;
        RECT 1857.120 1687.460 1857.380 1687.720 ;
        RECT 1870.460 1687.460 1870.720 1687.720 ;
      LAYER met2 ;
        RECT 1857.045 1700.000 1857.325 1704.000 ;
        RECT 1857.180 1687.750 1857.320 1700.000 ;
        RECT 1857.120 1687.430 1857.380 1687.750 ;
        RECT 1870.460 1687.430 1870.720 1687.750 ;
        RECT 1870.520 16.730 1870.660 1687.430 ;
        RECT 1870.520 16.590 1876.180 16.730 ;
        RECT 1876.040 2.400 1876.180 16.590 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1428.830 1678.140 1429.150 1678.200 ;
        RECT 1430.670 1678.140 1430.990 1678.200 ;
        RECT 1428.830 1678.000 1430.990 1678.140 ;
        RECT 1428.830 1677.940 1429.150 1678.000 ;
        RECT 1430.670 1677.940 1430.990 1678.000 ;
        RECT 752.170 47.500 752.490 47.560 ;
        RECT 1428.830 47.500 1429.150 47.560 ;
        RECT 752.170 47.360 1429.150 47.500 ;
        RECT 752.170 47.300 752.490 47.360 ;
        RECT 1428.830 47.300 1429.150 47.360 ;
      LAYER via ;
        RECT 1428.860 1677.940 1429.120 1678.200 ;
        RECT 1430.700 1677.940 1430.960 1678.200 ;
        RECT 752.200 47.300 752.460 47.560 ;
        RECT 1428.860 47.300 1429.120 47.560 ;
      LAYER met2 ;
        RECT 1432.465 1700.410 1432.745 1704.000 ;
        RECT 1430.760 1700.270 1432.745 1700.410 ;
        RECT 1430.760 1678.230 1430.900 1700.270 ;
        RECT 1432.465 1700.000 1432.745 1700.270 ;
        RECT 1428.860 1677.910 1429.120 1678.230 ;
        RECT 1430.700 1677.910 1430.960 1678.230 ;
        RECT 1428.920 47.590 1429.060 1677.910 ;
        RECT 752.200 47.270 752.460 47.590 ;
        RECT 1428.860 47.270 1429.120 47.590 ;
        RECT 752.260 2.400 752.400 47.270 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1863.530 1688.340 1863.850 1688.400 ;
        RECT 1869.510 1688.340 1869.830 1688.400 ;
        RECT 1863.530 1688.200 1869.830 1688.340 ;
        RECT 1863.530 1688.140 1863.850 1688.200 ;
        RECT 1869.510 1688.140 1869.830 1688.200 ;
        RECT 1869.510 17.240 1869.830 17.300 ;
        RECT 1893.890 17.240 1894.210 17.300 ;
        RECT 1869.510 17.100 1894.210 17.240 ;
        RECT 1869.510 17.040 1869.830 17.100 ;
        RECT 1893.890 17.040 1894.210 17.100 ;
      LAYER via ;
        RECT 1863.560 1688.140 1863.820 1688.400 ;
        RECT 1869.540 1688.140 1869.800 1688.400 ;
        RECT 1869.540 17.040 1869.800 17.300 ;
        RECT 1893.920 17.040 1894.180 17.300 ;
      LAYER met2 ;
        RECT 1863.485 1700.000 1863.765 1704.000 ;
        RECT 1863.620 1688.430 1863.760 1700.000 ;
        RECT 1863.560 1688.110 1863.820 1688.430 ;
        RECT 1869.540 1688.110 1869.800 1688.430 ;
        RECT 1869.600 17.330 1869.740 1688.110 ;
        RECT 1869.540 17.010 1869.800 17.330 ;
        RECT 1893.920 17.010 1894.180 17.330 ;
        RECT 1893.980 2.400 1894.120 17.010 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1870.430 1688.680 1870.750 1688.740 ;
        RECT 1876.410 1688.680 1876.730 1688.740 ;
        RECT 1870.430 1688.540 1876.730 1688.680 ;
        RECT 1870.430 1688.480 1870.750 1688.540 ;
        RECT 1876.410 1688.480 1876.730 1688.540 ;
        RECT 1876.410 16.560 1876.730 16.620 ;
        RECT 1911.830 16.560 1912.150 16.620 ;
        RECT 1876.410 16.420 1912.150 16.560 ;
        RECT 1876.410 16.360 1876.730 16.420 ;
        RECT 1911.830 16.360 1912.150 16.420 ;
      LAYER via ;
        RECT 1870.460 1688.480 1870.720 1688.740 ;
        RECT 1876.440 1688.480 1876.700 1688.740 ;
        RECT 1876.440 16.360 1876.700 16.620 ;
        RECT 1911.860 16.360 1912.120 16.620 ;
      LAYER met2 ;
        RECT 1870.385 1700.000 1870.665 1704.000 ;
        RECT 1870.520 1688.770 1870.660 1700.000 ;
        RECT 1870.460 1688.450 1870.720 1688.770 ;
        RECT 1876.440 1688.450 1876.700 1688.770 ;
        RECT 1876.500 16.650 1876.640 1688.450 ;
        RECT 1876.440 16.330 1876.700 16.650 ;
        RECT 1911.860 16.330 1912.120 16.650 ;
        RECT 1911.920 2.400 1912.060 16.330 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1876.870 1688.000 1877.190 1688.060 ;
        RECT 1883.310 1688.000 1883.630 1688.060 ;
        RECT 1876.870 1687.860 1883.630 1688.000 ;
        RECT 1876.870 1687.800 1877.190 1687.860 ;
        RECT 1883.310 1687.800 1883.630 1687.860 ;
        RECT 1883.310 18.600 1883.630 18.660 ;
        RECT 1929.310 18.600 1929.630 18.660 ;
        RECT 1883.310 18.460 1929.630 18.600 ;
        RECT 1883.310 18.400 1883.630 18.460 ;
        RECT 1929.310 18.400 1929.630 18.460 ;
      LAYER via ;
        RECT 1876.900 1687.800 1877.160 1688.060 ;
        RECT 1883.340 1687.800 1883.600 1688.060 ;
        RECT 1883.340 18.400 1883.600 18.660 ;
        RECT 1929.340 18.400 1929.600 18.660 ;
      LAYER met2 ;
        RECT 1876.825 1700.000 1877.105 1704.000 ;
        RECT 1876.960 1688.090 1877.100 1700.000 ;
        RECT 1876.900 1687.770 1877.160 1688.090 ;
        RECT 1883.340 1687.770 1883.600 1688.090 ;
        RECT 1883.400 18.690 1883.540 1687.770 ;
        RECT 1883.340 18.370 1883.600 18.690 ;
        RECT 1929.340 18.370 1929.600 18.690 ;
        RECT 1929.400 2.400 1929.540 18.370 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1883.770 1687.320 1884.090 1687.380 ;
        RECT 1890.210 1687.320 1890.530 1687.380 ;
        RECT 1883.770 1687.180 1890.530 1687.320 ;
        RECT 1883.770 1687.120 1884.090 1687.180 ;
        RECT 1890.210 1687.120 1890.530 1687.180 ;
        RECT 1890.210 17.920 1890.530 17.980 ;
        RECT 1947.250 17.920 1947.570 17.980 ;
        RECT 1890.210 17.780 1947.570 17.920 ;
        RECT 1890.210 17.720 1890.530 17.780 ;
        RECT 1947.250 17.720 1947.570 17.780 ;
      LAYER via ;
        RECT 1883.800 1687.120 1884.060 1687.380 ;
        RECT 1890.240 1687.120 1890.500 1687.380 ;
        RECT 1890.240 17.720 1890.500 17.980 ;
        RECT 1947.280 17.720 1947.540 17.980 ;
      LAYER met2 ;
        RECT 1883.725 1700.000 1884.005 1704.000 ;
        RECT 1883.860 1687.410 1884.000 1700.000 ;
        RECT 1883.800 1687.090 1884.060 1687.410 ;
        RECT 1890.240 1687.090 1890.500 1687.410 ;
        RECT 1890.300 18.010 1890.440 1687.090 ;
        RECT 1890.240 17.690 1890.500 18.010 ;
        RECT 1947.280 17.690 1947.540 18.010 ;
        RECT 1947.340 2.400 1947.480 17.690 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1908.700 1687.860 1925.860 1688.000 ;
        RECT 1890.670 1687.660 1890.990 1687.720 ;
        RECT 1908.700 1687.660 1908.840 1687.860 ;
        RECT 1890.670 1687.520 1908.840 1687.660 ;
        RECT 1925.720 1687.660 1925.860 1687.860 ;
        RECT 1935.290 1687.660 1935.610 1687.720 ;
        RECT 1925.720 1687.520 1935.610 1687.660 ;
        RECT 1890.670 1687.460 1890.990 1687.520 ;
        RECT 1935.290 1687.460 1935.610 1687.520 ;
        RECT 1935.290 19.280 1935.610 19.340 ;
        RECT 1965.190 19.280 1965.510 19.340 ;
        RECT 1935.290 19.140 1965.510 19.280 ;
        RECT 1935.290 19.080 1935.610 19.140 ;
        RECT 1965.190 19.080 1965.510 19.140 ;
      LAYER via ;
        RECT 1890.700 1687.460 1890.960 1687.720 ;
        RECT 1935.320 1687.460 1935.580 1687.720 ;
        RECT 1935.320 19.080 1935.580 19.340 ;
        RECT 1965.220 19.080 1965.480 19.340 ;
      LAYER met2 ;
        RECT 1890.625 1700.000 1890.905 1704.000 ;
        RECT 1890.760 1687.750 1890.900 1700.000 ;
        RECT 1890.700 1687.430 1890.960 1687.750 ;
        RECT 1935.320 1687.430 1935.580 1687.750 ;
        RECT 1935.380 19.370 1935.520 1687.430 ;
        RECT 1935.320 19.050 1935.580 19.370 ;
        RECT 1965.220 19.050 1965.480 19.370 ;
        RECT 1965.280 2.400 1965.420 19.050 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1929.845 1686.145 1930.015 1689.375 ;
      LAYER mcon ;
        RECT 1929.845 1689.205 1930.015 1689.375 ;
      LAYER met1 ;
        RECT 1897.110 1689.700 1897.430 1689.760 ;
        RECT 1897.110 1689.560 1916.200 1689.700 ;
        RECT 1897.110 1689.500 1897.430 1689.560 ;
        RECT 1916.060 1689.360 1916.200 1689.560 ;
        RECT 1929.785 1689.360 1930.075 1689.405 ;
        RECT 1916.060 1689.220 1930.075 1689.360 ;
        RECT 1929.785 1689.175 1930.075 1689.220 ;
        RECT 1929.785 1686.300 1930.075 1686.345 ;
        RECT 1962.890 1686.300 1963.210 1686.360 ;
        RECT 1929.785 1686.160 1963.210 1686.300 ;
        RECT 1929.785 1686.115 1930.075 1686.160 ;
        RECT 1962.890 1686.100 1963.210 1686.160 ;
        RECT 1962.890 14.520 1963.210 14.580 ;
        RECT 1983.130 14.520 1983.450 14.580 ;
        RECT 1962.890 14.380 1983.450 14.520 ;
        RECT 1962.890 14.320 1963.210 14.380 ;
        RECT 1983.130 14.320 1983.450 14.380 ;
      LAYER via ;
        RECT 1897.140 1689.500 1897.400 1689.760 ;
        RECT 1962.920 1686.100 1963.180 1686.360 ;
        RECT 1962.920 14.320 1963.180 14.580 ;
        RECT 1983.160 14.320 1983.420 14.580 ;
      LAYER met2 ;
        RECT 1897.065 1700.000 1897.345 1704.000 ;
        RECT 1897.200 1689.790 1897.340 1700.000 ;
        RECT 1897.140 1689.470 1897.400 1689.790 ;
        RECT 1962.920 1686.070 1963.180 1686.390 ;
        RECT 1962.980 14.610 1963.120 1686.070 ;
        RECT 1962.920 14.290 1963.180 14.610 ;
        RECT 1983.160 14.290 1983.420 14.610 ;
        RECT 1983.220 2.400 1983.360 14.290 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1919.265 1685.805 1919.435 1688.695 ;
        RECT 1942.725 1685.805 1942.895 1689.375 ;
      LAYER mcon ;
        RECT 1942.725 1689.205 1942.895 1689.375 ;
        RECT 1919.265 1688.525 1919.435 1688.695 ;
      LAYER met1 ;
        RECT 1904.010 1689.160 1904.330 1689.420 ;
        RECT 1942.665 1689.360 1942.955 1689.405 ;
        RECT 1976.690 1689.360 1977.010 1689.420 ;
        RECT 1942.665 1689.220 1977.010 1689.360 ;
        RECT 1942.665 1689.175 1942.955 1689.220 ;
        RECT 1976.690 1689.160 1977.010 1689.220 ;
        RECT 1904.100 1689.020 1904.240 1689.160 ;
        RECT 1904.100 1688.880 1911.600 1689.020 ;
        RECT 1911.460 1688.680 1911.600 1688.880 ;
        RECT 1919.205 1688.680 1919.495 1688.725 ;
        RECT 1911.460 1688.540 1919.495 1688.680 ;
        RECT 1919.205 1688.495 1919.495 1688.540 ;
        RECT 1919.205 1685.960 1919.495 1686.005 ;
        RECT 1942.665 1685.960 1942.955 1686.005 ;
        RECT 1919.205 1685.820 1942.955 1685.960 ;
        RECT 1919.205 1685.775 1919.495 1685.820 ;
        RECT 1942.665 1685.775 1942.955 1685.820 ;
        RECT 1976.690 17.240 1977.010 17.300 ;
        RECT 2001.070 17.240 2001.390 17.300 ;
        RECT 1976.690 17.100 2001.390 17.240 ;
        RECT 1976.690 17.040 1977.010 17.100 ;
        RECT 2001.070 17.040 2001.390 17.100 ;
      LAYER via ;
        RECT 1904.040 1689.160 1904.300 1689.420 ;
        RECT 1976.720 1689.160 1976.980 1689.420 ;
        RECT 1976.720 17.040 1976.980 17.300 ;
        RECT 2001.100 17.040 2001.360 17.300 ;
      LAYER met2 ;
        RECT 1903.965 1700.000 1904.245 1704.000 ;
        RECT 1904.100 1689.450 1904.240 1700.000 ;
        RECT 1904.040 1689.130 1904.300 1689.450 ;
        RECT 1976.720 1689.130 1976.980 1689.450 ;
        RECT 1976.780 17.330 1976.920 1689.130 ;
        RECT 1976.720 17.010 1976.980 17.330 ;
        RECT 2001.100 17.010 2001.360 17.330 ;
        RECT 2001.160 2.400 2001.300 17.010 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1910.450 15.880 1910.770 15.940 ;
        RECT 2018.550 15.880 2018.870 15.940 ;
        RECT 1910.450 15.740 2018.870 15.880 ;
        RECT 1910.450 15.680 1910.770 15.740 ;
        RECT 2018.550 15.680 2018.870 15.740 ;
      LAYER via ;
        RECT 1910.480 15.680 1910.740 15.940 ;
        RECT 2018.580 15.680 2018.840 15.940 ;
      LAYER met2 ;
        RECT 1910.865 1700.410 1911.145 1704.000 ;
        RECT 1910.540 1700.270 1911.145 1700.410 ;
        RECT 1910.540 15.970 1910.680 1700.270 ;
        RECT 1910.865 1700.000 1911.145 1700.270 ;
        RECT 1910.480 15.650 1910.740 15.970 ;
        RECT 2018.580 15.650 2018.840 15.970 ;
        RECT 2018.640 2.400 2018.780 15.650 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 16.560 1918.130 16.620 ;
        RECT 2036.490 16.560 2036.810 16.620 ;
        RECT 1917.810 16.420 2036.810 16.560 ;
        RECT 1917.810 16.360 1918.130 16.420 ;
        RECT 2036.490 16.360 2036.810 16.420 ;
      LAYER via ;
        RECT 1917.840 16.360 1918.100 16.620 ;
        RECT 2036.520 16.360 2036.780 16.620 ;
      LAYER met2 ;
        RECT 1917.305 1700.410 1917.585 1704.000 ;
        RECT 1917.305 1700.270 1918.040 1700.410 ;
        RECT 1917.305 1700.000 1917.585 1700.270 ;
        RECT 1917.900 16.650 1918.040 1700.270 ;
        RECT 1917.840 16.330 1918.100 16.650 ;
        RECT 2036.520 16.330 2036.780 16.650 ;
        RECT 2036.580 2.400 2036.720 16.330 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1952.845 1688.525 1953.015 1690.395 ;
      LAYER mcon ;
        RECT 1952.845 1690.225 1953.015 1690.395 ;
      LAYER met1 ;
        RECT 1924.250 1690.380 1924.570 1690.440 ;
        RECT 1952.785 1690.380 1953.075 1690.425 ;
        RECT 1924.250 1690.240 1953.075 1690.380 ;
        RECT 1924.250 1690.180 1924.570 1690.240 ;
        RECT 1952.785 1690.195 1953.075 1690.240 ;
        RECT 1997.390 1689.700 1997.710 1689.760 ;
        RECT 1979.540 1689.560 1997.710 1689.700 ;
        RECT 1952.785 1688.680 1953.075 1688.725 ;
        RECT 1979.540 1688.680 1979.680 1689.560 ;
        RECT 1997.390 1689.500 1997.710 1689.560 ;
        RECT 1952.785 1688.540 1979.680 1688.680 ;
        RECT 1952.785 1688.495 1953.075 1688.540 ;
        RECT 1997.390 14.520 1997.710 14.580 ;
        RECT 2054.430 14.520 2054.750 14.580 ;
        RECT 1997.390 14.380 2054.750 14.520 ;
        RECT 1997.390 14.320 1997.710 14.380 ;
        RECT 2054.430 14.320 2054.750 14.380 ;
      LAYER via ;
        RECT 1924.280 1690.180 1924.540 1690.440 ;
        RECT 1997.420 1689.500 1997.680 1689.760 ;
        RECT 1997.420 14.320 1997.680 14.580 ;
        RECT 2054.460 14.320 2054.720 14.580 ;
      LAYER met2 ;
        RECT 1924.205 1700.000 1924.485 1704.000 ;
        RECT 1924.340 1690.470 1924.480 1700.000 ;
        RECT 1924.280 1690.150 1924.540 1690.470 ;
        RECT 1997.420 1689.470 1997.680 1689.790 ;
        RECT 1997.480 14.610 1997.620 1689.470 ;
        RECT 1997.420 14.290 1997.680 14.610 ;
        RECT 2054.460 14.290 2054.720 14.610 ;
        RECT 2054.520 2.400 2054.660 14.290 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 772.410 49.880 772.730 49.940 ;
        RECT 1435.730 49.880 1436.050 49.940 ;
        RECT 772.410 49.740 1436.050 49.880 ;
        RECT 772.410 49.680 772.730 49.740 ;
        RECT 1435.730 49.680 1436.050 49.740 ;
        RECT 769.650 2.960 769.970 3.020 ;
        RECT 772.410 2.960 772.730 3.020 ;
        RECT 769.650 2.820 772.730 2.960 ;
        RECT 769.650 2.760 769.970 2.820 ;
        RECT 772.410 2.760 772.730 2.820 ;
      LAYER via ;
        RECT 772.440 49.680 772.700 49.940 ;
        RECT 1435.760 49.680 1436.020 49.940 ;
        RECT 769.680 2.760 769.940 3.020 ;
        RECT 772.440 2.760 772.700 3.020 ;
      LAYER met2 ;
        RECT 1439.365 1700.410 1439.645 1704.000 ;
        RECT 1437.660 1700.270 1439.645 1700.410 ;
        RECT 1437.660 1677.970 1437.800 1700.270 ;
        RECT 1439.365 1700.000 1439.645 1700.270 ;
        RECT 1435.820 1677.830 1437.800 1677.970 ;
        RECT 1435.820 49.970 1435.960 1677.830 ;
        RECT 772.440 49.650 772.700 49.970 ;
        RECT 1435.760 49.650 1436.020 49.970 ;
        RECT 772.500 3.050 772.640 49.650 ;
        RECT 769.680 2.730 769.940 3.050 ;
        RECT 772.440 2.730 772.700 3.050 ;
        RECT 769.740 2.400 769.880 2.730 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1970.325 18.105 1970.495 20.315 ;
      LAYER mcon ;
        RECT 1970.325 20.145 1970.495 20.315 ;
      LAYER met1 ;
        RECT 1970.265 20.300 1970.555 20.345 ;
        RECT 2072.370 20.300 2072.690 20.360 ;
        RECT 1970.265 20.160 2072.690 20.300 ;
        RECT 1970.265 20.115 1970.555 20.160 ;
        RECT 2072.370 20.100 2072.690 20.160 ;
        RECT 1931.610 18.600 1931.930 18.660 ;
        RECT 1931.610 18.460 1935.980 18.600 ;
        RECT 1931.610 18.400 1931.930 18.460 ;
        RECT 1935.840 18.260 1935.980 18.460 ;
        RECT 1970.265 18.260 1970.555 18.305 ;
        RECT 1935.840 18.120 1970.555 18.260 ;
        RECT 1970.265 18.075 1970.555 18.120 ;
      LAYER via ;
        RECT 2072.400 20.100 2072.660 20.360 ;
        RECT 1931.640 18.400 1931.900 18.660 ;
      LAYER met2 ;
        RECT 1931.105 1700.410 1931.385 1704.000 ;
        RECT 1931.105 1700.270 1931.840 1700.410 ;
        RECT 1931.105 1700.000 1931.385 1700.270 ;
        RECT 1931.700 18.690 1931.840 1700.270 ;
        RECT 2072.400 20.070 2072.660 20.390 ;
        RECT 1931.640 18.370 1931.900 18.690 ;
        RECT 2072.460 2.400 2072.600 20.070 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1938.510 20.640 1938.830 20.700 ;
        RECT 2089.850 20.640 2090.170 20.700 ;
        RECT 1938.510 20.500 2090.170 20.640 ;
        RECT 1938.510 20.440 1938.830 20.500 ;
        RECT 2089.850 20.440 2090.170 20.500 ;
      LAYER via ;
        RECT 1938.540 20.440 1938.800 20.700 ;
        RECT 2089.880 20.440 2090.140 20.700 ;
      LAYER met2 ;
        RECT 1937.545 1700.410 1937.825 1704.000 ;
        RECT 1937.545 1700.270 1938.740 1700.410 ;
        RECT 1937.545 1700.000 1937.825 1700.270 ;
        RECT 1938.600 20.730 1938.740 1700.270 ;
        RECT 1938.540 20.410 1938.800 20.730 ;
        RECT 2089.880 20.410 2090.140 20.730 ;
        RECT 2089.940 2.400 2090.080 20.410 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1945.410 19.960 1945.730 20.020 ;
        RECT 1945.410 19.820 1969.560 19.960 ;
        RECT 1945.410 19.760 1945.730 19.820 ;
        RECT 1969.420 19.280 1969.560 19.820 ;
        RECT 2107.790 19.280 2108.110 19.340 ;
        RECT 1969.420 19.140 2108.110 19.280 ;
        RECT 2107.790 19.080 2108.110 19.140 ;
      LAYER via ;
        RECT 1945.440 19.760 1945.700 20.020 ;
        RECT 2107.820 19.080 2108.080 19.340 ;
      LAYER met2 ;
        RECT 1944.445 1700.410 1944.725 1704.000 ;
        RECT 1944.445 1700.270 1945.640 1700.410 ;
        RECT 1944.445 1700.000 1944.725 1700.270 ;
        RECT 1945.500 20.050 1945.640 1700.270 ;
        RECT 1945.440 19.730 1945.700 20.050 ;
        RECT 2107.820 19.050 2108.080 19.370 ;
        RECT 2107.880 2.400 2108.020 19.050 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1984.585 1687.165 1984.755 1690.055 ;
      LAYER mcon ;
        RECT 1984.585 1689.885 1984.755 1690.055 ;
      LAYER met1 ;
        RECT 1951.390 1690.040 1951.710 1690.100 ;
        RECT 1984.525 1690.040 1984.815 1690.085 ;
        RECT 1951.390 1689.900 1984.815 1690.040 ;
        RECT 1951.390 1689.840 1951.710 1689.900 ;
        RECT 1984.525 1689.855 1984.815 1689.900 ;
        RECT 1984.525 1687.320 1984.815 1687.365 ;
        RECT 2011.190 1687.320 2011.510 1687.380 ;
        RECT 1984.525 1687.180 2011.510 1687.320 ;
        RECT 1984.525 1687.135 1984.815 1687.180 ;
        RECT 2011.190 1687.120 2011.510 1687.180 ;
        RECT 2013.030 15.200 2013.350 15.260 ;
        RECT 2125.730 15.200 2126.050 15.260 ;
        RECT 2013.030 15.060 2126.050 15.200 ;
        RECT 2013.030 15.000 2013.350 15.060 ;
        RECT 2125.730 15.000 2126.050 15.060 ;
      LAYER via ;
        RECT 1951.420 1689.840 1951.680 1690.100 ;
        RECT 2011.220 1687.120 2011.480 1687.380 ;
        RECT 2013.060 15.000 2013.320 15.260 ;
        RECT 2125.760 15.000 2126.020 15.260 ;
      LAYER met2 ;
        RECT 1951.345 1700.000 1951.625 1704.000 ;
        RECT 1951.480 1690.130 1951.620 1700.000 ;
        RECT 1951.420 1689.810 1951.680 1690.130 ;
        RECT 2011.220 1687.090 2011.480 1687.410 ;
        RECT 2011.280 24.890 2011.420 1687.090 ;
        RECT 2011.280 24.750 2013.260 24.890 ;
        RECT 2013.120 15.290 2013.260 24.750 ;
        RECT 2013.060 14.970 2013.320 15.290 ;
        RECT 2125.760 14.970 2126.020 15.290 ;
        RECT 2125.820 2.400 2125.960 14.970 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1972.165 17.425 1972.335 18.615 ;
      LAYER mcon ;
        RECT 1972.165 18.445 1972.335 18.615 ;
      LAYER met1 ;
        RECT 1972.105 18.600 1972.395 18.645 ;
        RECT 2143.670 18.600 2143.990 18.660 ;
        RECT 1972.105 18.460 2143.990 18.600 ;
        RECT 1972.105 18.415 1972.395 18.460 ;
        RECT 2143.670 18.400 2143.990 18.460 ;
        RECT 1958.750 17.920 1959.070 17.980 ;
        RECT 1958.750 17.780 1959.900 17.920 ;
        RECT 1958.750 17.720 1959.070 17.780 ;
        RECT 1959.760 17.580 1959.900 17.780 ;
        RECT 1972.105 17.580 1972.395 17.625 ;
        RECT 1959.760 17.440 1972.395 17.580 ;
        RECT 1972.105 17.395 1972.395 17.440 ;
      LAYER via ;
        RECT 2143.700 18.400 2143.960 18.660 ;
        RECT 1958.780 17.720 1959.040 17.980 ;
      LAYER met2 ;
        RECT 1957.785 1700.410 1958.065 1704.000 ;
        RECT 1957.785 1700.270 1959.440 1700.410 ;
        RECT 1957.785 1700.000 1958.065 1700.270 ;
        RECT 1959.300 40.530 1959.440 1700.270 ;
        RECT 1958.840 40.390 1959.440 40.530 ;
        RECT 1958.840 18.010 1958.980 40.390 ;
        RECT 2143.700 18.370 2143.960 18.690 ;
        RECT 1958.780 17.690 1959.040 18.010 ;
        RECT 2143.760 2.400 2143.900 18.370 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1966.110 17.920 1966.430 17.980 ;
        RECT 2161.610 17.920 2161.930 17.980 ;
        RECT 1966.110 17.780 2161.930 17.920 ;
        RECT 1966.110 17.720 1966.430 17.780 ;
        RECT 2161.610 17.720 2161.930 17.780 ;
      LAYER via ;
        RECT 1966.140 17.720 1966.400 17.980 ;
        RECT 2161.640 17.720 2161.900 17.980 ;
      LAYER met2 ;
        RECT 1964.685 1700.410 1964.965 1704.000 ;
        RECT 1964.685 1700.270 1966.340 1700.410 ;
        RECT 1964.685 1700.000 1964.965 1700.270 ;
        RECT 1966.200 18.010 1966.340 1700.270 ;
        RECT 1966.140 17.690 1966.400 18.010 ;
        RECT 2161.640 17.690 2161.900 18.010 ;
        RECT 2161.700 2.400 2161.840 17.690 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1973.010 17.580 1973.330 17.640 ;
        RECT 2179.090 17.580 2179.410 17.640 ;
        RECT 1973.010 17.440 2179.410 17.580 ;
        RECT 1973.010 17.380 1973.330 17.440 ;
        RECT 2179.090 17.380 2179.410 17.440 ;
      LAYER via ;
        RECT 1973.040 17.380 1973.300 17.640 ;
        RECT 2179.120 17.380 2179.380 17.640 ;
      LAYER met2 ;
        RECT 1971.125 1700.410 1971.405 1704.000 ;
        RECT 1971.125 1700.270 1973.240 1700.410 ;
        RECT 1971.125 1700.000 1971.405 1700.270 ;
        RECT 1973.100 17.670 1973.240 1700.270 ;
        RECT 1973.040 17.350 1973.300 17.670 ;
        RECT 2179.120 17.350 2179.380 17.670 ;
        RECT 2179.180 2.400 2179.320 17.350 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2001.605 14.705 2001.775 17.255 ;
      LAYER mcon ;
        RECT 2001.605 17.085 2001.775 17.255 ;
      LAYER met1 ;
        RECT 2001.545 17.240 2001.835 17.285 ;
        RECT 2197.030 17.240 2197.350 17.300 ;
        RECT 2001.545 17.100 2197.350 17.240 ;
        RECT 2001.545 17.055 2001.835 17.100 ;
        RECT 2197.030 17.040 2197.350 17.100 ;
        RECT 1979.910 14.860 1980.230 14.920 ;
        RECT 2001.545 14.860 2001.835 14.905 ;
        RECT 1979.910 14.720 2001.835 14.860 ;
        RECT 1979.910 14.660 1980.230 14.720 ;
        RECT 2001.545 14.675 2001.835 14.720 ;
      LAYER via ;
        RECT 2197.060 17.040 2197.320 17.300 ;
        RECT 1979.940 14.660 1980.200 14.920 ;
      LAYER met2 ;
        RECT 1978.025 1700.410 1978.305 1704.000 ;
        RECT 1978.025 1700.270 1980.140 1700.410 ;
        RECT 1978.025 1700.000 1978.305 1700.270 ;
        RECT 1980.000 14.950 1980.140 1700.270 ;
        RECT 2197.060 17.010 2197.320 17.330 ;
        RECT 1979.940 14.630 1980.200 14.950 ;
        RECT 2197.120 2.400 2197.260 17.010 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1984.970 1690.040 1985.290 1690.100 ;
        RECT 2031.890 1690.040 2032.210 1690.100 ;
        RECT 1984.970 1689.900 2032.210 1690.040 ;
        RECT 1984.970 1689.840 1985.290 1689.900 ;
        RECT 2031.890 1689.840 2032.210 1689.900 ;
        RECT 2031.890 14.180 2032.210 14.240 ;
        RECT 2214.970 14.180 2215.290 14.240 ;
        RECT 2031.890 14.040 2215.290 14.180 ;
        RECT 2031.890 13.980 2032.210 14.040 ;
        RECT 2214.970 13.980 2215.290 14.040 ;
      LAYER via ;
        RECT 1985.000 1689.840 1985.260 1690.100 ;
        RECT 2031.920 1689.840 2032.180 1690.100 ;
        RECT 2031.920 13.980 2032.180 14.240 ;
        RECT 2215.000 13.980 2215.260 14.240 ;
      LAYER met2 ;
        RECT 1984.925 1700.000 1985.205 1704.000 ;
        RECT 1985.060 1690.130 1985.200 1700.000 ;
        RECT 1985.000 1689.810 1985.260 1690.130 ;
        RECT 2031.920 1689.810 2032.180 1690.130 ;
        RECT 2031.980 14.270 2032.120 1689.810 ;
        RECT 2031.920 13.950 2032.180 14.270 ;
        RECT 2215.000 13.950 2215.260 14.270 ;
        RECT 2215.060 2.400 2215.200 13.950 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2111.545 14.705 2111.715 16.235 ;
        RECT 2135.465 15.045 2135.635 16.235 ;
        RECT 2163.065 15.045 2163.235 16.235 ;
        RECT 2209.985 14.705 2210.155 16.235 ;
      LAYER mcon ;
        RECT 2111.545 16.065 2111.715 16.235 ;
        RECT 2135.465 16.065 2135.635 16.235 ;
        RECT 2163.065 16.065 2163.235 16.235 ;
        RECT 2209.985 16.065 2210.155 16.235 ;
      LAYER met1 ;
        RECT 1991.410 1689.360 1991.730 1689.420 ;
        RECT 2045.690 1689.360 2046.010 1689.420 ;
        RECT 1991.410 1689.220 2046.010 1689.360 ;
        RECT 1991.410 1689.160 1991.730 1689.220 ;
        RECT 2045.690 1689.160 2046.010 1689.220 ;
        RECT 2045.690 16.220 2046.010 16.280 ;
        RECT 2062.710 16.220 2063.030 16.280 ;
        RECT 2045.690 16.080 2063.030 16.220 ;
        RECT 2045.690 16.020 2046.010 16.080 ;
        RECT 2062.710 16.020 2063.030 16.080 ;
        RECT 2111.485 16.220 2111.775 16.265 ;
        RECT 2135.405 16.220 2135.695 16.265 ;
        RECT 2111.485 16.080 2135.695 16.220 ;
        RECT 2111.485 16.035 2111.775 16.080 ;
        RECT 2135.405 16.035 2135.695 16.080 ;
        RECT 2163.005 16.220 2163.295 16.265 ;
        RECT 2209.925 16.220 2210.215 16.265 ;
        RECT 2163.005 16.080 2210.215 16.220 ;
        RECT 2163.005 16.035 2163.295 16.080 ;
        RECT 2209.925 16.035 2210.215 16.080 ;
        RECT 2135.405 15.200 2135.695 15.245 ;
        RECT 2163.005 15.200 2163.295 15.245 ;
        RECT 2135.405 15.060 2163.295 15.200 ;
        RECT 2135.405 15.015 2135.695 15.060 ;
        RECT 2163.005 15.015 2163.295 15.060 ;
        RECT 2062.710 14.860 2063.030 14.920 ;
        RECT 2111.485 14.860 2111.775 14.905 ;
        RECT 2062.710 14.720 2111.775 14.860 ;
        RECT 2062.710 14.660 2063.030 14.720 ;
        RECT 2111.485 14.675 2111.775 14.720 ;
        RECT 2209.925 14.860 2210.215 14.905 ;
        RECT 2232.910 14.860 2233.230 14.920 ;
        RECT 2209.925 14.720 2233.230 14.860 ;
        RECT 2209.925 14.675 2210.215 14.720 ;
        RECT 2232.910 14.660 2233.230 14.720 ;
      LAYER via ;
        RECT 1991.440 1689.160 1991.700 1689.420 ;
        RECT 2045.720 1689.160 2045.980 1689.420 ;
        RECT 2045.720 16.020 2045.980 16.280 ;
        RECT 2062.740 16.020 2063.000 16.280 ;
        RECT 2062.740 14.660 2063.000 14.920 ;
        RECT 2232.940 14.660 2233.200 14.920 ;
      LAYER met2 ;
        RECT 1991.365 1700.000 1991.645 1704.000 ;
        RECT 1991.500 1689.450 1991.640 1700.000 ;
        RECT 1991.440 1689.130 1991.700 1689.450 ;
        RECT 2045.720 1689.130 2045.980 1689.450 ;
        RECT 2045.780 16.310 2045.920 1689.130 ;
        RECT 2045.720 15.990 2045.980 16.310 ;
        RECT 2062.740 15.990 2063.000 16.310 ;
        RECT 2062.800 14.950 2062.940 15.990 ;
        RECT 2062.740 14.630 2063.000 14.950 ;
        RECT 2232.940 14.630 2233.200 14.950 ;
        RECT 2233.000 2.400 2233.140 14.630 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 49.540 793.430 49.600 ;
        RECT 1442.630 49.540 1442.950 49.600 ;
        RECT 793.110 49.400 1442.950 49.540 ;
        RECT 793.110 49.340 793.430 49.400 ;
        RECT 1442.630 49.340 1442.950 49.400 ;
        RECT 787.590 2.960 787.910 3.020 ;
        RECT 793.110 2.960 793.430 3.020 ;
        RECT 787.590 2.820 793.430 2.960 ;
        RECT 787.590 2.760 787.910 2.820 ;
        RECT 793.110 2.760 793.430 2.820 ;
      LAYER via ;
        RECT 793.140 49.340 793.400 49.600 ;
        RECT 1442.660 49.340 1442.920 49.600 ;
        RECT 787.620 2.760 787.880 3.020 ;
        RECT 793.140 2.760 793.400 3.020 ;
      LAYER met2 ;
        RECT 1446.265 1700.410 1446.545 1704.000 ;
        RECT 1444.560 1700.270 1446.545 1700.410 ;
        RECT 1444.560 1677.970 1444.700 1700.270 ;
        RECT 1446.265 1700.000 1446.545 1700.270 ;
        RECT 1442.720 1677.830 1444.700 1677.970 ;
        RECT 1442.720 49.630 1442.860 1677.830 ;
        RECT 793.140 49.310 793.400 49.630 ;
        RECT 1442.660 49.310 1442.920 49.630 ;
        RECT 793.200 3.050 793.340 49.310 ;
        RECT 787.620 2.730 787.880 3.050 ;
        RECT 793.140 2.730 793.400 3.050 ;
        RECT 787.680 2.400 787.820 2.730 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2038.865 1683.765 2039.035 1685.635 ;
        RECT 2187.905 1683.765 2188.995 1683.935 ;
      LAYER mcon ;
        RECT 2038.865 1685.465 2039.035 1685.635 ;
        RECT 2188.825 1683.765 2188.995 1683.935 ;
      LAYER met1 ;
        RECT 1998.310 1685.620 1998.630 1685.680 ;
        RECT 2038.805 1685.620 2039.095 1685.665 ;
        RECT 1998.310 1685.480 2039.095 1685.620 ;
        RECT 1998.310 1685.420 1998.630 1685.480 ;
        RECT 2038.805 1685.435 2039.095 1685.480 ;
        RECT 2038.805 1683.920 2039.095 1683.965 ;
        RECT 2187.845 1683.920 2188.135 1683.965 ;
        RECT 2038.805 1683.780 2188.135 1683.920 ;
        RECT 2038.805 1683.735 2039.095 1683.780 ;
        RECT 2187.845 1683.735 2188.135 1683.780 ;
        RECT 2188.765 1683.920 2189.055 1683.965 ;
        RECT 2188.765 1683.780 2234.980 1683.920 ;
        RECT 2188.765 1683.735 2189.055 1683.780 ;
        RECT 2234.840 1683.580 2234.980 1683.780 ;
        RECT 2249.470 1683.580 2249.790 1683.640 ;
        RECT 2234.840 1683.440 2249.790 1683.580 ;
        RECT 2249.470 1683.380 2249.790 1683.440 ;
      LAYER via ;
        RECT 1998.340 1685.420 1998.600 1685.680 ;
        RECT 2249.500 1683.380 2249.760 1683.640 ;
      LAYER met2 ;
        RECT 1998.265 1700.000 1998.545 1704.000 ;
        RECT 1998.400 1685.710 1998.540 1700.000 ;
        RECT 1998.340 1685.390 1998.600 1685.710 ;
        RECT 2249.500 1683.350 2249.760 1683.670 ;
        RECT 2249.560 3.130 2249.700 1683.350 ;
        RECT 2249.560 2.990 2251.080 3.130 ;
        RECT 2250.940 2.400 2251.080 2.990 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2112.005 14.365 2112.175 16.915 ;
        RECT 2135.925 16.065 2136.095 16.915 ;
        RECT 2162.605 14.365 2162.775 16.235 ;
        RECT 2210.905 14.365 2211.075 17.255 ;
      LAYER mcon ;
        RECT 2210.905 17.085 2211.075 17.255 ;
        RECT 2112.005 16.745 2112.175 16.915 ;
        RECT 2135.925 16.745 2136.095 16.915 ;
        RECT 2162.605 16.065 2162.775 16.235 ;
      LAYER met1 ;
        RECT 2005.210 1688.340 2005.530 1688.400 ;
        RECT 2052.590 1688.340 2052.910 1688.400 ;
        RECT 2005.210 1688.200 2052.910 1688.340 ;
        RECT 2005.210 1688.140 2005.530 1688.200 ;
        RECT 2052.590 1688.140 2052.910 1688.200 ;
        RECT 2210.845 17.240 2211.135 17.285 ;
        RECT 2268.330 17.240 2268.650 17.300 ;
        RECT 2210.845 17.100 2268.650 17.240 ;
        RECT 2210.845 17.055 2211.135 17.100 ;
        RECT 2268.330 17.040 2268.650 17.100 ;
        RECT 2111.945 16.900 2112.235 16.945 ;
        RECT 2135.865 16.900 2136.155 16.945 ;
        RECT 2111.945 16.760 2136.155 16.900 ;
        RECT 2111.945 16.715 2112.235 16.760 ;
        RECT 2135.865 16.715 2136.155 16.760 ;
        RECT 2135.865 16.220 2136.155 16.265 ;
        RECT 2162.545 16.220 2162.835 16.265 ;
        RECT 2135.865 16.080 2162.835 16.220 ;
        RECT 2135.865 16.035 2136.155 16.080 ;
        RECT 2162.545 16.035 2162.835 16.080 ;
        RECT 2052.590 14.860 2052.910 14.920 ;
        RECT 2052.590 14.720 2062.480 14.860 ;
        RECT 2052.590 14.660 2052.910 14.720 ;
        RECT 2062.340 14.520 2062.480 14.720 ;
        RECT 2111.945 14.520 2112.235 14.565 ;
        RECT 2062.340 14.380 2112.235 14.520 ;
        RECT 2111.945 14.335 2112.235 14.380 ;
        RECT 2162.545 14.520 2162.835 14.565 ;
        RECT 2210.845 14.520 2211.135 14.565 ;
        RECT 2162.545 14.380 2211.135 14.520 ;
        RECT 2162.545 14.335 2162.835 14.380 ;
        RECT 2210.845 14.335 2211.135 14.380 ;
      LAYER via ;
        RECT 2005.240 1688.140 2005.500 1688.400 ;
        RECT 2052.620 1688.140 2052.880 1688.400 ;
        RECT 2268.360 17.040 2268.620 17.300 ;
        RECT 2052.620 14.660 2052.880 14.920 ;
      LAYER met2 ;
        RECT 2005.165 1700.000 2005.445 1704.000 ;
        RECT 2005.300 1688.430 2005.440 1700.000 ;
        RECT 2005.240 1688.110 2005.500 1688.430 ;
        RECT 2052.620 1688.110 2052.880 1688.430 ;
        RECT 2052.680 14.950 2052.820 1688.110 ;
        RECT 2268.360 17.010 2268.620 17.330 ;
        RECT 2052.620 14.630 2052.880 14.950 ;
        RECT 2268.420 2.400 2268.560 17.010 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2011.650 1684.600 2011.970 1684.660 ;
        RECT 2011.650 1684.460 2016.020 1684.600 ;
        RECT 2011.650 1684.400 2011.970 1684.460 ;
        RECT 2015.880 1684.260 2016.020 1684.460 ;
        RECT 2283.970 1684.260 2284.290 1684.320 ;
        RECT 2015.880 1684.120 2284.290 1684.260 ;
        RECT 2283.970 1684.060 2284.290 1684.120 ;
      LAYER via ;
        RECT 2011.680 1684.400 2011.940 1684.660 ;
        RECT 2284.000 1684.060 2284.260 1684.320 ;
      LAYER met2 ;
        RECT 2011.605 1700.000 2011.885 1704.000 ;
        RECT 2011.740 1684.690 2011.880 1700.000 ;
        RECT 2011.680 1684.370 2011.940 1684.690 ;
        RECT 2284.000 1684.030 2284.260 1684.350 ;
        RECT 2284.060 16.730 2284.200 1684.030 ;
        RECT 2284.060 16.590 2286.500 16.730 ;
        RECT 2286.360 2.400 2286.500 16.590 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2018.550 1689.020 2018.870 1689.080 ;
        RECT 2059.490 1689.020 2059.810 1689.080 ;
        RECT 2018.550 1688.880 2059.810 1689.020 ;
        RECT 2018.550 1688.820 2018.870 1688.880 ;
        RECT 2059.490 1688.820 2059.810 1688.880 ;
        RECT 2059.490 15.880 2059.810 15.940 ;
        RECT 2059.490 15.740 2061.100 15.880 ;
        RECT 2059.490 15.680 2059.810 15.740 ;
        RECT 2060.960 15.540 2061.100 15.740 ;
        RECT 2304.210 15.540 2304.530 15.600 ;
        RECT 2060.960 15.400 2304.530 15.540 ;
        RECT 2304.210 15.340 2304.530 15.400 ;
      LAYER via ;
        RECT 2018.580 1688.820 2018.840 1689.080 ;
        RECT 2059.520 1688.820 2059.780 1689.080 ;
        RECT 2059.520 15.680 2059.780 15.940 ;
        RECT 2304.240 15.340 2304.500 15.600 ;
      LAYER met2 ;
        RECT 2018.505 1700.000 2018.785 1704.000 ;
        RECT 2018.640 1689.110 2018.780 1700.000 ;
        RECT 2018.580 1688.790 2018.840 1689.110 ;
        RECT 2059.520 1688.790 2059.780 1689.110 ;
        RECT 2059.580 15.970 2059.720 1688.790 ;
        RECT 2059.520 15.650 2059.780 15.970 ;
        RECT 2304.240 15.310 2304.500 15.630 ;
        RECT 2304.300 2.400 2304.440 15.310 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2026.830 1684.600 2027.150 1684.660 ;
        RECT 2318.470 1684.600 2318.790 1684.660 ;
        RECT 2026.830 1684.460 2318.790 1684.600 ;
        RECT 2026.830 1684.400 2027.150 1684.460 ;
        RECT 2318.470 1684.400 2318.790 1684.460 ;
      LAYER via ;
        RECT 2026.860 1684.400 2027.120 1684.660 ;
        RECT 2318.500 1684.400 2318.760 1684.660 ;
      LAYER met2 ;
        RECT 2025.405 1700.410 2025.685 1704.000 ;
        RECT 2025.405 1700.270 2027.060 1700.410 ;
        RECT 2025.405 1700.000 2025.685 1700.270 ;
        RECT 2026.920 1684.690 2027.060 1700.270 ;
        RECT 2026.860 1684.370 2027.120 1684.690 ;
        RECT 2318.500 1684.370 2318.760 1684.690 ;
        RECT 2318.560 17.410 2318.700 1684.370 ;
        RECT 2318.560 17.270 2322.380 17.410 ;
        RECT 2322.240 2.400 2322.380 17.270 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2033.730 1689.700 2034.050 1689.760 ;
        RECT 2033.730 1689.560 2075.360 1689.700 ;
        RECT 2033.730 1689.500 2034.050 1689.560 ;
        RECT 2075.220 1689.360 2075.360 1689.560 ;
        RECT 2087.090 1689.360 2087.410 1689.420 ;
        RECT 2075.220 1689.220 2087.410 1689.360 ;
        RECT 2087.090 1689.160 2087.410 1689.220 ;
        RECT 2087.090 15.880 2087.410 15.940 ;
        RECT 2339.630 15.880 2339.950 15.940 ;
        RECT 2087.090 15.740 2339.950 15.880 ;
        RECT 2087.090 15.680 2087.410 15.740 ;
        RECT 2339.630 15.680 2339.950 15.740 ;
      LAYER via ;
        RECT 2033.760 1689.500 2034.020 1689.760 ;
        RECT 2087.120 1689.160 2087.380 1689.420 ;
        RECT 2087.120 15.680 2087.380 15.940 ;
        RECT 2339.660 15.680 2339.920 15.940 ;
      LAYER met2 ;
        RECT 2031.845 1700.410 2032.125 1704.000 ;
        RECT 2031.845 1700.270 2033.960 1700.410 ;
        RECT 2031.845 1700.000 2032.125 1700.270 ;
        RECT 2033.820 1689.790 2033.960 1700.270 ;
        RECT 2033.760 1689.470 2034.020 1689.790 ;
        RECT 2087.120 1689.130 2087.380 1689.450 ;
        RECT 2087.180 15.970 2087.320 1689.130 ;
        RECT 2087.120 15.650 2087.380 15.970 ;
        RECT 2339.660 15.650 2339.920 15.970 ;
        RECT 2339.720 2.400 2339.860 15.650 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2087.165 1684.785 2087.335 1686.315 ;
      LAYER mcon ;
        RECT 2087.165 1686.145 2087.335 1686.315 ;
      LAYER met1 ;
        RECT 2040.170 1686.300 2040.490 1686.360 ;
        RECT 2087.105 1686.300 2087.395 1686.345 ;
        RECT 2040.170 1686.160 2087.395 1686.300 ;
        RECT 2040.170 1686.100 2040.490 1686.160 ;
        RECT 2087.105 1686.115 2087.395 1686.160 ;
        RECT 2087.105 1684.940 2087.395 1684.985 ;
        RECT 2352.970 1684.940 2353.290 1685.000 ;
        RECT 2087.105 1684.800 2353.290 1684.940 ;
        RECT 2087.105 1684.755 2087.395 1684.800 ;
        RECT 2352.970 1684.740 2353.290 1684.800 ;
      LAYER via ;
        RECT 2040.200 1686.100 2040.460 1686.360 ;
        RECT 2353.000 1684.740 2353.260 1685.000 ;
      LAYER met2 ;
        RECT 2038.745 1700.410 2039.025 1704.000 ;
        RECT 2038.745 1700.270 2040.400 1700.410 ;
        RECT 2038.745 1700.000 2039.025 1700.270 ;
        RECT 2040.260 1686.390 2040.400 1700.270 ;
        RECT 2040.200 1686.070 2040.460 1686.390 ;
        RECT 2353.000 1684.710 2353.260 1685.030 ;
        RECT 2353.060 16.730 2353.200 1684.710 ;
        RECT 2353.060 16.590 2357.800 16.730 ;
        RECT 2357.660 2.400 2357.800 16.590 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2100.890 1689.020 2101.210 1689.080 ;
        RECT 2069.700 1688.880 2101.210 1689.020 ;
        RECT 2045.230 1688.680 2045.550 1688.740 ;
        RECT 2069.700 1688.680 2069.840 1688.880 ;
        RECT 2100.890 1688.820 2101.210 1688.880 ;
        RECT 2045.230 1688.540 2069.840 1688.680 ;
        RECT 2045.230 1688.480 2045.550 1688.540 ;
        RECT 2100.890 16.560 2101.210 16.620 ;
        RECT 2375.510 16.560 2375.830 16.620 ;
        RECT 2100.890 16.420 2375.830 16.560 ;
        RECT 2100.890 16.360 2101.210 16.420 ;
        RECT 2375.510 16.360 2375.830 16.420 ;
      LAYER via ;
        RECT 2045.260 1688.480 2045.520 1688.740 ;
        RECT 2100.920 1688.820 2101.180 1689.080 ;
        RECT 2100.920 16.360 2101.180 16.620 ;
        RECT 2375.540 16.360 2375.800 16.620 ;
      LAYER met2 ;
        RECT 2045.185 1700.000 2045.465 1704.000 ;
        RECT 2045.320 1688.770 2045.460 1700.000 ;
        RECT 2100.920 1688.790 2101.180 1689.110 ;
        RECT 2045.260 1688.450 2045.520 1688.770 ;
        RECT 2100.980 16.650 2101.120 1688.790 ;
        RECT 2100.920 16.330 2101.180 16.650 ;
        RECT 2375.540 16.330 2375.800 16.650 ;
        RECT 2375.600 2.400 2375.740 16.330 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2052.130 1685.620 2052.450 1685.680 ;
        RECT 2387.470 1685.620 2387.790 1685.680 ;
        RECT 2052.130 1685.480 2387.790 1685.620 ;
        RECT 2052.130 1685.420 2052.450 1685.480 ;
        RECT 2387.470 1685.420 2387.790 1685.480 ;
        RECT 2387.470 20.980 2387.790 21.040 ;
        RECT 2393.450 20.980 2393.770 21.040 ;
        RECT 2387.470 20.840 2393.770 20.980 ;
        RECT 2387.470 20.780 2387.790 20.840 ;
        RECT 2393.450 20.780 2393.770 20.840 ;
      LAYER via ;
        RECT 2052.160 1685.420 2052.420 1685.680 ;
        RECT 2387.500 1685.420 2387.760 1685.680 ;
        RECT 2387.500 20.780 2387.760 21.040 ;
        RECT 2393.480 20.780 2393.740 21.040 ;
      LAYER met2 ;
        RECT 2052.085 1700.000 2052.365 1704.000 ;
        RECT 2052.220 1685.710 2052.360 1700.000 ;
        RECT 2052.160 1685.390 2052.420 1685.710 ;
        RECT 2387.500 1685.390 2387.760 1685.710 ;
        RECT 2387.560 21.070 2387.700 1685.390 ;
        RECT 2387.500 20.750 2387.760 21.070 ;
        RECT 2393.480 20.750 2393.740 21.070 ;
        RECT 2393.540 2.400 2393.680 20.750 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2163.525 1687.165 2163.695 1689.375 ;
        RECT 2186.525 1683.085 2186.695 1689.375 ;
        RECT 2233.445 14.705 2233.615 17.595 ;
      LAYER mcon ;
        RECT 2163.525 1689.205 2163.695 1689.375 ;
        RECT 2186.525 1689.205 2186.695 1689.375 ;
        RECT 2233.445 17.425 2233.615 17.595 ;
      LAYER met1 ;
        RECT 2163.465 1689.360 2163.755 1689.405 ;
        RECT 2186.465 1689.360 2186.755 1689.405 ;
        RECT 2163.465 1689.220 2186.755 1689.360 ;
        RECT 2163.465 1689.175 2163.755 1689.220 ;
        RECT 2186.465 1689.175 2186.755 1689.220 ;
        RECT 2059.030 1687.660 2059.350 1687.720 ;
        RECT 2059.030 1687.520 2141.140 1687.660 ;
        RECT 2059.030 1687.460 2059.350 1687.520 ;
        RECT 2141.000 1687.320 2141.140 1687.520 ;
        RECT 2163.465 1687.320 2163.755 1687.365 ;
        RECT 2141.000 1687.180 2163.755 1687.320 ;
        RECT 2163.465 1687.135 2163.755 1687.180 ;
        RECT 2186.465 1683.240 2186.755 1683.285 ;
        RECT 2190.590 1683.240 2190.910 1683.300 ;
        RECT 2186.465 1683.100 2190.910 1683.240 ;
        RECT 2186.465 1683.055 2186.755 1683.100 ;
        RECT 2190.590 1683.040 2190.910 1683.100 ;
        RECT 2190.590 17.580 2190.910 17.640 ;
        RECT 2233.385 17.580 2233.675 17.625 ;
        RECT 2190.590 17.440 2233.675 17.580 ;
        RECT 2190.590 17.380 2190.910 17.440 ;
        RECT 2233.385 17.395 2233.675 17.440 ;
        RECT 2233.385 14.860 2233.675 14.905 ;
        RECT 2411.390 14.860 2411.710 14.920 ;
        RECT 2233.385 14.720 2411.710 14.860 ;
        RECT 2233.385 14.675 2233.675 14.720 ;
        RECT 2411.390 14.660 2411.710 14.720 ;
      LAYER via ;
        RECT 2059.060 1687.460 2059.320 1687.720 ;
        RECT 2190.620 1683.040 2190.880 1683.300 ;
        RECT 2190.620 17.380 2190.880 17.640 ;
        RECT 2411.420 14.660 2411.680 14.920 ;
      LAYER met2 ;
        RECT 2058.985 1700.000 2059.265 1704.000 ;
        RECT 2059.120 1687.750 2059.260 1700.000 ;
        RECT 2059.060 1687.430 2059.320 1687.750 ;
        RECT 2190.620 1683.010 2190.880 1683.330 ;
        RECT 2190.680 17.670 2190.820 1683.010 ;
        RECT 2190.620 17.350 2190.880 17.670 ;
        RECT 2411.420 14.630 2411.680 14.950 ;
        RECT 2411.480 2.400 2411.620 14.630 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 49.200 807.230 49.260 ;
        RECT 1449.530 49.200 1449.850 49.260 ;
        RECT 806.910 49.060 1449.850 49.200 ;
        RECT 806.910 49.000 807.230 49.060 ;
        RECT 1449.530 49.000 1449.850 49.060 ;
        RECT 805.530 2.960 805.850 3.020 ;
        RECT 806.910 2.960 807.230 3.020 ;
        RECT 805.530 2.820 807.230 2.960 ;
        RECT 805.530 2.760 805.850 2.820 ;
        RECT 806.910 2.760 807.230 2.820 ;
      LAYER via ;
        RECT 806.940 49.000 807.200 49.260 ;
        RECT 1449.560 49.000 1449.820 49.260 ;
        RECT 805.560 2.760 805.820 3.020 ;
        RECT 806.940 2.760 807.200 3.020 ;
      LAYER met2 ;
        RECT 1452.705 1700.410 1452.985 1704.000 ;
        RECT 1451.000 1700.270 1452.985 1700.410 ;
        RECT 1451.000 1677.970 1451.140 1700.270 ;
        RECT 1452.705 1700.000 1452.985 1700.270 ;
        RECT 1449.620 1677.830 1451.140 1677.970 ;
        RECT 1449.620 49.290 1449.760 1677.830 ;
        RECT 806.940 48.970 807.200 49.290 ;
        RECT 1449.560 48.970 1449.820 49.290 ;
        RECT 807.000 3.050 807.140 48.970 ;
        RECT 805.560 2.730 805.820 3.050 ;
        RECT 806.940 2.730 807.200 3.050 ;
        RECT 805.620 2.400 805.760 2.730 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1120.705 21.165 1120.875 24.055 ;
      LAYER mcon ;
        RECT 1120.705 23.885 1120.875 24.055 ;
      LAYER met1 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 1120.645 24.040 1120.935 24.085 ;
        RECT 2.830 23.900 1120.935 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 1120.645 23.855 1120.935 23.900 ;
        RECT 1120.645 21.320 1120.935 21.365 ;
        RECT 1145.470 21.320 1145.790 21.380 ;
        RECT 1120.645 21.180 1145.790 21.320 ;
        RECT 1120.645 21.135 1120.935 21.180 ;
        RECT 1145.470 21.120 1145.790 21.180 ;
      LAYER via ;
        RECT 2.860 23.840 3.120 24.100 ;
        RECT 1145.500 21.120 1145.760 21.380 ;
      LAYER met2 ;
        RECT 1150.025 1700.410 1150.305 1704.000 ;
        RECT 1145.560 1700.270 1150.305 1700.410 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 1145.560 21.410 1145.700 1700.270 ;
        RECT 1150.025 1700.000 1150.305 1700.270 ;
        RECT 1145.500 21.090 1145.760 21.410 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1146.465 1490.645 1146.635 1497.955 ;
        RECT 1146.925 1365.525 1147.095 1400.715 ;
        RECT 1146.925 1317.245 1147.095 1352.435 ;
        RECT 1146.925 1268.965 1147.095 1304.155 ;
        RECT 1146.465 1076.185 1146.635 1103.895 ;
        RECT 1146.465 531.505 1146.635 579.615 ;
        RECT 1146.465 434.945 1146.635 483.055 ;
        RECT 1146.465 324.785 1146.635 372.555 ;
        RECT 1146.465 193.545 1146.635 207.315 ;
        RECT 1146.005 41.565 1146.175 89.675 ;
        RECT 13.945 23.545 14.115 24.395 ;
        RECT 62.245 23.545 62.415 24.395 ;
        RECT 96.745 23.545 96.915 24.395 ;
        RECT 158.845 23.545 159.015 24.395 ;
        RECT 207.145 23.545 207.315 24.395 ;
        RECT 255.445 23.545 255.615 24.395 ;
        RECT 303.745 23.545 303.915 24.395 ;
        RECT 641.845 23.545 642.015 24.395 ;
        RECT 690.145 23.545 690.315 24.395 ;
        RECT 738.445 23.545 738.615 24.395 ;
        RECT 786.745 23.545 786.915 24.395 ;
        RECT 835.045 23.545 835.215 24.395 ;
        RECT 869.545 23.545 869.715 24.395 ;
        RECT 931.645 23.545 931.815 24.395 ;
        RECT 979.945 23.545 980.115 24.395 ;
        RECT 1028.245 22.865 1028.415 24.395 ;
        RECT 1076.085 22.865 1076.255 24.395 ;
      LAYER mcon ;
        RECT 1146.465 1497.785 1146.635 1497.955 ;
        RECT 1146.925 1400.545 1147.095 1400.715 ;
        RECT 1146.925 1352.265 1147.095 1352.435 ;
        RECT 1146.925 1303.985 1147.095 1304.155 ;
        RECT 1146.465 1103.725 1146.635 1103.895 ;
        RECT 1146.465 579.445 1146.635 579.615 ;
        RECT 1146.465 482.885 1146.635 483.055 ;
        RECT 1146.465 372.385 1146.635 372.555 ;
        RECT 1146.465 207.145 1146.635 207.315 ;
        RECT 1146.005 89.505 1146.175 89.675 ;
        RECT 13.945 24.225 14.115 24.395 ;
        RECT 62.245 24.225 62.415 24.395 ;
        RECT 96.745 24.225 96.915 24.395 ;
        RECT 158.845 24.225 159.015 24.395 ;
        RECT 207.145 24.225 207.315 24.395 ;
        RECT 255.445 24.225 255.615 24.395 ;
        RECT 303.745 24.225 303.915 24.395 ;
        RECT 641.845 24.225 642.015 24.395 ;
        RECT 690.145 24.225 690.315 24.395 ;
        RECT 738.445 24.225 738.615 24.395 ;
        RECT 786.745 24.225 786.915 24.395 ;
        RECT 835.045 24.225 835.215 24.395 ;
        RECT 869.545 24.225 869.715 24.395 ;
        RECT 931.645 24.225 931.815 24.395 ;
        RECT 979.945 24.225 980.115 24.395 ;
        RECT 1028.245 24.225 1028.415 24.395 ;
        RECT 1076.085 24.225 1076.255 24.395 ;
      LAYER met1 ;
        RECT 1146.390 1607.760 1146.710 1607.820 ;
        RECT 1147.310 1607.760 1147.630 1607.820 ;
        RECT 1146.390 1607.620 1147.630 1607.760 ;
        RECT 1146.390 1607.560 1146.710 1607.620 ;
        RECT 1147.310 1607.560 1147.630 1607.620 ;
        RECT 1147.310 1569.680 1147.630 1569.740 ;
        RECT 1148.230 1569.680 1148.550 1569.740 ;
        RECT 1147.310 1569.540 1148.550 1569.680 ;
        RECT 1147.310 1569.480 1147.630 1569.540 ;
        RECT 1148.230 1569.480 1148.550 1569.540 ;
        RECT 1147.310 1545.540 1147.630 1545.600 ;
        RECT 1148.230 1545.540 1148.550 1545.600 ;
        RECT 1147.310 1545.400 1148.550 1545.540 ;
        RECT 1147.310 1545.340 1147.630 1545.400 ;
        RECT 1148.230 1545.340 1148.550 1545.400 ;
        RECT 1146.405 1497.940 1146.695 1497.985 ;
        RECT 1147.310 1497.940 1147.630 1498.000 ;
        RECT 1146.405 1497.800 1147.630 1497.940 ;
        RECT 1146.405 1497.755 1146.695 1497.800 ;
        RECT 1147.310 1497.740 1147.630 1497.800 ;
        RECT 1146.390 1490.800 1146.710 1490.860 ;
        RECT 1146.195 1490.660 1146.710 1490.800 ;
        RECT 1146.390 1490.600 1146.710 1490.660 ;
        RECT 1146.850 1462.240 1147.170 1462.300 ;
        RECT 1147.770 1462.240 1148.090 1462.300 ;
        RECT 1146.850 1462.100 1148.090 1462.240 ;
        RECT 1146.850 1462.040 1147.170 1462.100 ;
        RECT 1147.770 1462.040 1148.090 1462.100 ;
        RECT 1146.850 1414.780 1147.170 1415.040 ;
        RECT 1146.940 1414.020 1147.080 1414.780 ;
        RECT 1146.850 1413.760 1147.170 1414.020 ;
        RECT 1146.850 1400.700 1147.170 1400.760 ;
        RECT 1146.655 1400.560 1147.170 1400.700 ;
        RECT 1146.850 1400.500 1147.170 1400.560 ;
        RECT 1146.850 1365.680 1147.170 1365.740 ;
        RECT 1146.655 1365.540 1147.170 1365.680 ;
        RECT 1146.850 1365.480 1147.170 1365.540 ;
        RECT 1146.850 1352.420 1147.170 1352.480 ;
        RECT 1146.655 1352.280 1147.170 1352.420 ;
        RECT 1146.850 1352.220 1147.170 1352.280 ;
        RECT 1146.850 1317.400 1147.170 1317.460 ;
        RECT 1146.655 1317.260 1147.170 1317.400 ;
        RECT 1146.850 1317.200 1147.170 1317.260 ;
        RECT 1146.850 1304.140 1147.170 1304.200 ;
        RECT 1146.655 1304.000 1147.170 1304.140 ;
        RECT 1146.850 1303.940 1147.170 1304.000 ;
        RECT 1146.850 1269.120 1147.170 1269.180 ;
        RECT 1146.655 1268.980 1147.170 1269.120 ;
        RECT 1146.850 1268.920 1147.170 1268.980 ;
        RECT 1146.850 1221.860 1147.170 1221.920 ;
        RECT 1146.480 1221.720 1147.170 1221.860 ;
        RECT 1146.480 1221.240 1146.620 1221.720 ;
        RECT 1146.850 1221.660 1147.170 1221.720 ;
        RECT 1146.390 1220.980 1146.710 1221.240 ;
        RECT 1146.850 1152.500 1147.170 1152.560 ;
        RECT 1147.770 1152.500 1148.090 1152.560 ;
        RECT 1146.850 1152.360 1148.090 1152.500 ;
        RECT 1146.850 1152.300 1147.170 1152.360 ;
        RECT 1147.770 1152.300 1148.090 1152.360 ;
        RECT 1146.850 1125.300 1147.170 1125.360 ;
        RECT 1146.480 1125.160 1147.170 1125.300 ;
        RECT 1146.480 1124.680 1146.620 1125.160 ;
        RECT 1146.850 1125.100 1147.170 1125.160 ;
        RECT 1146.390 1124.420 1146.710 1124.680 ;
        RECT 1146.390 1103.880 1146.710 1103.940 ;
        RECT 1146.195 1103.740 1146.710 1103.880 ;
        RECT 1146.390 1103.680 1146.710 1103.740 ;
        RECT 1146.390 1076.340 1146.710 1076.400 ;
        RECT 1146.195 1076.200 1146.710 1076.340 ;
        RECT 1146.390 1076.140 1146.710 1076.200 ;
        RECT 1146.390 1014.460 1146.710 1014.520 ;
        RECT 1146.850 1014.460 1147.170 1014.520 ;
        RECT 1146.390 1014.320 1147.170 1014.460 ;
        RECT 1146.390 1014.260 1146.710 1014.320 ;
        RECT 1146.850 1014.260 1147.170 1014.320 ;
        RECT 1146.850 966.180 1147.170 966.240 ;
        RECT 1147.770 966.180 1148.090 966.240 ;
        RECT 1146.850 966.040 1148.090 966.180 ;
        RECT 1146.850 965.980 1147.170 966.040 ;
        RECT 1147.770 965.980 1148.090 966.040 ;
        RECT 1146.850 869.620 1147.170 869.680 ;
        RECT 1147.770 869.620 1148.090 869.680 ;
        RECT 1146.850 869.480 1148.090 869.620 ;
        RECT 1146.850 869.420 1147.170 869.480 ;
        RECT 1147.770 869.420 1148.090 869.480 ;
        RECT 1146.390 786.800 1146.710 787.060 ;
        RECT 1146.480 786.660 1146.620 786.800 ;
        RECT 1146.850 786.660 1147.170 786.720 ;
        RECT 1146.480 786.520 1147.170 786.660 ;
        RECT 1146.850 786.460 1147.170 786.520 ;
        RECT 1146.850 772.720 1147.170 772.780 ;
        RECT 1147.770 772.720 1148.090 772.780 ;
        RECT 1146.850 772.580 1148.090 772.720 ;
        RECT 1146.850 772.520 1147.170 772.580 ;
        RECT 1147.770 772.520 1148.090 772.580 ;
        RECT 1146.390 689.900 1146.710 690.160 ;
        RECT 1146.480 689.760 1146.620 689.900 ;
        RECT 1146.850 689.760 1147.170 689.820 ;
        RECT 1146.480 689.620 1147.170 689.760 ;
        RECT 1146.850 689.560 1147.170 689.620 ;
        RECT 1146.850 676.160 1147.170 676.220 ;
        RECT 1147.770 676.160 1148.090 676.220 ;
        RECT 1146.850 676.020 1148.090 676.160 ;
        RECT 1146.850 675.960 1147.170 676.020 ;
        RECT 1147.770 675.960 1148.090 676.020 ;
        RECT 1146.390 593.340 1146.710 593.600 ;
        RECT 1146.480 593.200 1146.620 593.340 ;
        RECT 1146.850 593.200 1147.170 593.260 ;
        RECT 1146.480 593.060 1147.170 593.200 ;
        RECT 1146.850 593.000 1147.170 593.060 ;
        RECT 1146.405 579.600 1146.695 579.645 ;
        RECT 1146.850 579.600 1147.170 579.660 ;
        RECT 1146.405 579.460 1147.170 579.600 ;
        RECT 1146.405 579.415 1146.695 579.460 ;
        RECT 1146.850 579.400 1147.170 579.460 ;
        RECT 1146.390 531.660 1146.710 531.720 ;
        RECT 1146.195 531.520 1146.710 531.660 ;
        RECT 1146.390 531.460 1146.710 531.520 ;
        RECT 1146.390 496.780 1146.710 497.040 ;
        RECT 1146.480 496.640 1146.620 496.780 ;
        RECT 1146.850 496.640 1147.170 496.700 ;
        RECT 1146.480 496.500 1147.170 496.640 ;
        RECT 1146.850 496.440 1147.170 496.500 ;
        RECT 1146.405 483.040 1146.695 483.085 ;
        RECT 1146.850 483.040 1147.170 483.100 ;
        RECT 1146.405 482.900 1147.170 483.040 ;
        RECT 1146.405 482.855 1146.695 482.900 ;
        RECT 1146.850 482.840 1147.170 482.900 ;
        RECT 1146.390 435.100 1146.710 435.160 ;
        RECT 1146.195 434.960 1146.710 435.100 ;
        RECT 1146.390 434.900 1146.710 434.960 ;
        RECT 1146.390 400.220 1146.710 400.480 ;
        RECT 1146.480 399.740 1146.620 400.220 ;
        RECT 1146.850 399.740 1147.170 399.800 ;
        RECT 1146.480 399.600 1147.170 399.740 ;
        RECT 1146.850 399.540 1147.170 399.600 ;
        RECT 1146.405 372.540 1146.695 372.585 ;
        RECT 1146.850 372.540 1147.170 372.600 ;
        RECT 1146.405 372.400 1147.170 372.540 ;
        RECT 1146.405 372.355 1146.695 372.400 ;
        RECT 1146.850 372.340 1147.170 372.400 ;
        RECT 1146.390 324.940 1146.710 325.000 ;
        RECT 1146.195 324.800 1146.710 324.940 ;
        RECT 1146.390 324.740 1146.710 324.800 ;
        RECT 1146.390 324.260 1146.710 324.320 ;
        RECT 1147.310 324.260 1147.630 324.320 ;
        RECT 1146.390 324.120 1147.630 324.260 ;
        RECT 1146.390 324.060 1146.710 324.120 ;
        RECT 1147.310 324.060 1147.630 324.120 ;
        RECT 1146.850 255.580 1147.170 255.640 ;
        RECT 1146.480 255.440 1147.170 255.580 ;
        RECT 1146.480 255.300 1146.620 255.440 ;
        RECT 1146.850 255.380 1147.170 255.440 ;
        RECT 1146.390 255.040 1146.710 255.300 ;
        RECT 1146.390 207.300 1146.710 207.360 ;
        RECT 1146.195 207.160 1146.710 207.300 ;
        RECT 1146.390 207.100 1146.710 207.160 ;
        RECT 1146.405 193.700 1146.695 193.745 ;
        RECT 1146.850 193.700 1147.170 193.760 ;
        RECT 1146.405 193.560 1147.170 193.700 ;
        RECT 1146.405 193.515 1146.695 193.560 ;
        RECT 1146.850 193.500 1147.170 193.560 ;
        RECT 1146.390 158.820 1146.710 159.080 ;
        RECT 1146.480 158.340 1146.620 158.820 ;
        RECT 1146.850 158.340 1147.170 158.400 ;
        RECT 1146.480 158.200 1147.170 158.340 ;
        RECT 1146.850 158.140 1147.170 158.200 ;
        RECT 1145.945 89.660 1146.235 89.705 ;
        RECT 1146.850 89.660 1147.170 89.720 ;
        RECT 1145.945 89.520 1147.170 89.660 ;
        RECT 1145.945 89.475 1146.235 89.520 ;
        RECT 1146.850 89.460 1147.170 89.520 ;
        RECT 1145.930 41.720 1146.250 41.780 ;
        RECT 1145.735 41.580 1146.250 41.720 ;
        RECT 1145.930 41.520 1146.250 41.580 ;
        RECT 13.885 24.380 14.175 24.425 ;
        RECT 62.185 24.380 62.475 24.425 ;
        RECT 13.885 24.240 62.475 24.380 ;
        RECT 13.885 24.195 14.175 24.240 ;
        RECT 62.185 24.195 62.475 24.240 ;
        RECT 96.685 24.380 96.975 24.425 ;
        RECT 158.785 24.380 159.075 24.425 ;
        RECT 96.685 24.240 159.075 24.380 ;
        RECT 96.685 24.195 96.975 24.240 ;
        RECT 158.785 24.195 159.075 24.240 ;
        RECT 207.085 24.380 207.375 24.425 ;
        RECT 255.385 24.380 255.675 24.425 ;
        RECT 207.085 24.240 255.675 24.380 ;
        RECT 207.085 24.195 207.375 24.240 ;
        RECT 255.385 24.195 255.675 24.240 ;
        RECT 303.685 24.380 303.975 24.425 ;
        RECT 641.785 24.380 642.075 24.425 ;
        RECT 303.685 24.240 642.075 24.380 ;
        RECT 303.685 24.195 303.975 24.240 ;
        RECT 641.785 24.195 642.075 24.240 ;
        RECT 690.085 24.380 690.375 24.425 ;
        RECT 738.385 24.380 738.675 24.425 ;
        RECT 690.085 24.240 738.675 24.380 ;
        RECT 690.085 24.195 690.375 24.240 ;
        RECT 738.385 24.195 738.675 24.240 ;
        RECT 786.685 24.380 786.975 24.425 ;
        RECT 834.985 24.380 835.275 24.425 ;
        RECT 786.685 24.240 835.275 24.380 ;
        RECT 786.685 24.195 786.975 24.240 ;
        RECT 834.985 24.195 835.275 24.240 ;
        RECT 869.485 24.380 869.775 24.425 ;
        RECT 931.585 24.380 931.875 24.425 ;
        RECT 869.485 24.240 931.875 24.380 ;
        RECT 869.485 24.195 869.775 24.240 ;
        RECT 931.585 24.195 931.875 24.240 ;
        RECT 979.885 24.380 980.175 24.425 ;
        RECT 1028.185 24.380 1028.475 24.425 ;
        RECT 979.885 24.240 1028.475 24.380 ;
        RECT 979.885 24.195 980.175 24.240 ;
        RECT 1028.185 24.195 1028.475 24.240 ;
        RECT 1076.025 24.380 1076.315 24.425 ;
        RECT 1145.930 24.380 1146.250 24.440 ;
        RECT 1076.025 24.240 1146.250 24.380 ;
        RECT 1076.025 24.195 1076.315 24.240 ;
        RECT 1145.930 24.180 1146.250 24.240 ;
        RECT 8.350 23.700 8.670 23.760 ;
        RECT 13.885 23.700 14.175 23.745 ;
        RECT 8.350 23.560 14.175 23.700 ;
        RECT 8.350 23.500 8.670 23.560 ;
        RECT 13.885 23.515 14.175 23.560 ;
        RECT 62.185 23.700 62.475 23.745 ;
        RECT 96.685 23.700 96.975 23.745 ;
        RECT 62.185 23.560 96.975 23.700 ;
        RECT 62.185 23.515 62.475 23.560 ;
        RECT 96.685 23.515 96.975 23.560 ;
        RECT 158.785 23.700 159.075 23.745 ;
        RECT 207.085 23.700 207.375 23.745 ;
        RECT 158.785 23.560 207.375 23.700 ;
        RECT 158.785 23.515 159.075 23.560 ;
        RECT 207.085 23.515 207.375 23.560 ;
        RECT 255.385 23.700 255.675 23.745 ;
        RECT 303.685 23.700 303.975 23.745 ;
        RECT 255.385 23.560 303.975 23.700 ;
        RECT 255.385 23.515 255.675 23.560 ;
        RECT 303.685 23.515 303.975 23.560 ;
        RECT 641.785 23.700 642.075 23.745 ;
        RECT 690.085 23.700 690.375 23.745 ;
        RECT 641.785 23.560 690.375 23.700 ;
        RECT 641.785 23.515 642.075 23.560 ;
        RECT 690.085 23.515 690.375 23.560 ;
        RECT 738.385 23.700 738.675 23.745 ;
        RECT 786.685 23.700 786.975 23.745 ;
        RECT 738.385 23.560 786.975 23.700 ;
        RECT 738.385 23.515 738.675 23.560 ;
        RECT 786.685 23.515 786.975 23.560 ;
        RECT 834.985 23.700 835.275 23.745 ;
        RECT 869.485 23.700 869.775 23.745 ;
        RECT 834.985 23.560 869.775 23.700 ;
        RECT 834.985 23.515 835.275 23.560 ;
        RECT 869.485 23.515 869.775 23.560 ;
        RECT 931.585 23.700 931.875 23.745 ;
        RECT 979.885 23.700 980.175 23.745 ;
        RECT 931.585 23.560 980.175 23.700 ;
        RECT 931.585 23.515 931.875 23.560 ;
        RECT 979.885 23.515 980.175 23.560 ;
        RECT 1028.185 23.020 1028.475 23.065 ;
        RECT 1076.025 23.020 1076.315 23.065 ;
        RECT 1028.185 22.880 1076.315 23.020 ;
        RECT 1028.185 22.835 1028.475 22.880 ;
        RECT 1076.025 22.835 1076.315 22.880 ;
      LAYER via ;
        RECT 1146.420 1607.560 1146.680 1607.820 ;
        RECT 1147.340 1607.560 1147.600 1607.820 ;
        RECT 1147.340 1569.480 1147.600 1569.740 ;
        RECT 1148.260 1569.480 1148.520 1569.740 ;
        RECT 1147.340 1545.340 1147.600 1545.600 ;
        RECT 1148.260 1545.340 1148.520 1545.600 ;
        RECT 1147.340 1497.740 1147.600 1498.000 ;
        RECT 1146.420 1490.600 1146.680 1490.860 ;
        RECT 1146.880 1462.040 1147.140 1462.300 ;
        RECT 1147.800 1462.040 1148.060 1462.300 ;
        RECT 1146.880 1414.780 1147.140 1415.040 ;
        RECT 1146.880 1413.760 1147.140 1414.020 ;
        RECT 1146.880 1400.500 1147.140 1400.760 ;
        RECT 1146.880 1365.480 1147.140 1365.740 ;
        RECT 1146.880 1352.220 1147.140 1352.480 ;
        RECT 1146.880 1317.200 1147.140 1317.460 ;
        RECT 1146.880 1303.940 1147.140 1304.200 ;
        RECT 1146.880 1268.920 1147.140 1269.180 ;
        RECT 1146.880 1221.660 1147.140 1221.920 ;
        RECT 1146.420 1220.980 1146.680 1221.240 ;
        RECT 1146.880 1152.300 1147.140 1152.560 ;
        RECT 1147.800 1152.300 1148.060 1152.560 ;
        RECT 1146.880 1125.100 1147.140 1125.360 ;
        RECT 1146.420 1124.420 1146.680 1124.680 ;
        RECT 1146.420 1103.680 1146.680 1103.940 ;
        RECT 1146.420 1076.140 1146.680 1076.400 ;
        RECT 1146.420 1014.260 1146.680 1014.520 ;
        RECT 1146.880 1014.260 1147.140 1014.520 ;
        RECT 1146.880 965.980 1147.140 966.240 ;
        RECT 1147.800 965.980 1148.060 966.240 ;
        RECT 1146.880 869.420 1147.140 869.680 ;
        RECT 1147.800 869.420 1148.060 869.680 ;
        RECT 1146.420 786.800 1146.680 787.060 ;
        RECT 1146.880 786.460 1147.140 786.720 ;
        RECT 1146.880 772.520 1147.140 772.780 ;
        RECT 1147.800 772.520 1148.060 772.780 ;
        RECT 1146.420 689.900 1146.680 690.160 ;
        RECT 1146.880 689.560 1147.140 689.820 ;
        RECT 1146.880 675.960 1147.140 676.220 ;
        RECT 1147.800 675.960 1148.060 676.220 ;
        RECT 1146.420 593.340 1146.680 593.600 ;
        RECT 1146.880 593.000 1147.140 593.260 ;
        RECT 1146.880 579.400 1147.140 579.660 ;
        RECT 1146.420 531.460 1146.680 531.720 ;
        RECT 1146.420 496.780 1146.680 497.040 ;
        RECT 1146.880 496.440 1147.140 496.700 ;
        RECT 1146.880 482.840 1147.140 483.100 ;
        RECT 1146.420 434.900 1146.680 435.160 ;
        RECT 1146.420 400.220 1146.680 400.480 ;
        RECT 1146.880 399.540 1147.140 399.800 ;
        RECT 1146.880 372.340 1147.140 372.600 ;
        RECT 1146.420 324.740 1146.680 325.000 ;
        RECT 1146.420 324.060 1146.680 324.320 ;
        RECT 1147.340 324.060 1147.600 324.320 ;
        RECT 1146.880 255.380 1147.140 255.640 ;
        RECT 1146.420 255.040 1146.680 255.300 ;
        RECT 1146.420 207.100 1146.680 207.360 ;
        RECT 1146.880 193.500 1147.140 193.760 ;
        RECT 1146.420 158.820 1146.680 159.080 ;
        RECT 1146.880 158.140 1147.140 158.400 ;
        RECT 1146.880 89.460 1147.140 89.720 ;
        RECT 1145.960 41.520 1146.220 41.780 ;
        RECT 1145.960 24.180 1146.220 24.440 ;
        RECT 8.380 23.500 8.640 23.760 ;
      LAYER met2 ;
        RECT 1151.865 1700.410 1152.145 1704.000 ;
        RECT 1150.620 1700.270 1152.145 1700.410 ;
        RECT 1150.620 1677.970 1150.760 1700.270 ;
        RECT 1151.865 1700.000 1152.145 1700.270 ;
        RECT 1146.480 1677.830 1150.760 1677.970 ;
        RECT 1146.480 1607.850 1146.620 1677.830 ;
        RECT 1146.420 1607.530 1146.680 1607.850 ;
        RECT 1147.340 1607.530 1147.600 1607.850 ;
        RECT 1147.400 1569.770 1147.540 1607.530 ;
        RECT 1147.340 1569.450 1147.600 1569.770 ;
        RECT 1148.260 1569.450 1148.520 1569.770 ;
        RECT 1148.320 1545.630 1148.460 1569.450 ;
        RECT 1147.340 1545.310 1147.600 1545.630 ;
        RECT 1148.260 1545.310 1148.520 1545.630 ;
        RECT 1147.400 1498.030 1147.540 1545.310 ;
        RECT 1147.340 1497.710 1147.600 1498.030 ;
        RECT 1146.420 1490.570 1146.680 1490.890 ;
        RECT 1146.480 1490.290 1146.620 1490.570 ;
        RECT 1146.870 1490.290 1147.150 1490.405 ;
        RECT 1146.480 1490.150 1147.150 1490.290 ;
        RECT 1146.870 1490.035 1147.150 1490.150 ;
        RECT 1147.790 1490.035 1148.070 1490.405 ;
        RECT 1147.860 1462.330 1148.000 1490.035 ;
        RECT 1146.880 1462.010 1147.140 1462.330 ;
        RECT 1147.800 1462.010 1148.060 1462.330 ;
        RECT 1146.940 1415.070 1147.080 1462.010 ;
        RECT 1146.880 1414.750 1147.140 1415.070 ;
        RECT 1146.880 1413.730 1147.140 1414.050 ;
        RECT 1146.940 1400.790 1147.080 1413.730 ;
        RECT 1146.880 1400.470 1147.140 1400.790 ;
        RECT 1146.880 1365.450 1147.140 1365.770 ;
        RECT 1146.940 1352.510 1147.080 1365.450 ;
        RECT 1146.880 1352.190 1147.140 1352.510 ;
        RECT 1146.880 1317.170 1147.140 1317.490 ;
        RECT 1146.940 1304.230 1147.080 1317.170 ;
        RECT 1146.880 1303.910 1147.140 1304.230 ;
        RECT 1146.880 1268.890 1147.140 1269.210 ;
        RECT 1146.940 1221.950 1147.080 1268.890 ;
        RECT 1146.880 1221.630 1147.140 1221.950 ;
        RECT 1146.420 1220.950 1146.680 1221.270 ;
        RECT 1146.480 1200.725 1146.620 1220.950 ;
        RECT 1146.410 1200.355 1146.690 1200.725 ;
        RECT 1147.790 1200.355 1148.070 1200.725 ;
        RECT 1147.860 1152.590 1148.000 1200.355 ;
        RECT 1146.880 1152.270 1147.140 1152.590 ;
        RECT 1147.800 1152.270 1148.060 1152.590 ;
        RECT 1146.940 1125.390 1147.080 1152.270 ;
        RECT 1146.880 1125.070 1147.140 1125.390 ;
        RECT 1146.420 1124.390 1146.680 1124.710 ;
        RECT 1146.480 1103.970 1146.620 1124.390 ;
        RECT 1146.420 1103.650 1146.680 1103.970 ;
        RECT 1146.420 1076.110 1146.680 1076.430 ;
        RECT 1146.480 1055.770 1146.620 1076.110 ;
        RECT 1146.480 1055.630 1147.080 1055.770 ;
        RECT 1146.940 1014.550 1147.080 1055.630 ;
        RECT 1146.420 1014.405 1146.680 1014.550 ;
        RECT 1146.410 1014.035 1146.690 1014.405 ;
        RECT 1146.880 1014.230 1147.140 1014.550 ;
        RECT 1147.790 1014.035 1148.070 1014.405 ;
        RECT 1147.860 966.270 1148.000 1014.035 ;
        RECT 1146.880 965.950 1147.140 966.270 ;
        RECT 1147.800 965.950 1148.060 966.270 ;
        RECT 1146.940 931.330 1147.080 965.950 ;
        RECT 1146.480 931.190 1147.080 931.330 ;
        RECT 1146.480 917.845 1146.620 931.190 ;
        RECT 1146.410 917.475 1146.690 917.845 ;
        RECT 1147.790 917.475 1148.070 917.845 ;
        RECT 1147.860 869.710 1148.000 917.475 ;
        RECT 1146.880 869.390 1147.140 869.710 ;
        RECT 1147.800 869.390 1148.060 869.710 ;
        RECT 1146.940 834.770 1147.080 869.390 ;
        RECT 1146.480 834.630 1147.080 834.770 ;
        RECT 1146.480 787.090 1146.620 834.630 ;
        RECT 1146.420 786.770 1146.680 787.090 ;
        RECT 1146.880 786.430 1147.140 786.750 ;
        RECT 1146.940 772.810 1147.080 786.430 ;
        RECT 1146.880 772.490 1147.140 772.810 ;
        RECT 1147.800 772.490 1148.060 772.810 ;
        RECT 1147.860 724.725 1148.000 772.490 ;
        RECT 1146.410 724.355 1146.690 724.725 ;
        RECT 1147.790 724.355 1148.070 724.725 ;
        RECT 1146.480 690.190 1146.620 724.355 ;
        RECT 1146.420 689.870 1146.680 690.190 ;
        RECT 1146.880 689.530 1147.140 689.850 ;
        RECT 1146.940 676.250 1147.080 689.530 ;
        RECT 1146.880 675.930 1147.140 676.250 ;
        RECT 1147.800 675.930 1148.060 676.250 ;
        RECT 1147.860 628.165 1148.000 675.930 ;
        RECT 1146.410 627.795 1146.690 628.165 ;
        RECT 1147.790 627.795 1148.070 628.165 ;
        RECT 1146.480 593.630 1146.620 627.795 ;
        RECT 1146.420 593.310 1146.680 593.630 ;
        RECT 1146.880 592.970 1147.140 593.290 ;
        RECT 1146.940 579.690 1147.080 592.970 ;
        RECT 1146.880 579.370 1147.140 579.690 ;
        RECT 1146.420 531.430 1146.680 531.750 ;
        RECT 1146.480 497.070 1146.620 531.430 ;
        RECT 1146.420 496.750 1146.680 497.070 ;
        RECT 1146.880 496.410 1147.140 496.730 ;
        RECT 1146.940 483.130 1147.080 496.410 ;
        RECT 1146.880 482.810 1147.140 483.130 ;
        RECT 1146.420 434.870 1146.680 435.190 ;
        RECT 1146.480 400.510 1146.620 434.870 ;
        RECT 1146.420 400.190 1146.680 400.510 ;
        RECT 1146.880 399.510 1147.140 399.830 ;
        RECT 1146.940 372.630 1147.080 399.510 ;
        RECT 1146.880 372.310 1147.140 372.630 ;
        RECT 1146.420 324.710 1146.680 325.030 ;
        RECT 1146.480 324.350 1146.620 324.710 ;
        RECT 1146.420 324.030 1146.680 324.350 ;
        RECT 1147.340 324.030 1147.600 324.350 ;
        RECT 1147.400 303.010 1147.540 324.030 ;
        RECT 1146.940 302.870 1147.540 303.010 ;
        RECT 1146.940 255.670 1147.080 302.870 ;
        RECT 1146.880 255.350 1147.140 255.670 ;
        RECT 1146.420 255.010 1146.680 255.330 ;
        RECT 1146.480 207.390 1146.620 255.010 ;
        RECT 1146.420 207.070 1146.680 207.390 ;
        RECT 1146.880 193.530 1147.140 193.790 ;
        RECT 1146.480 193.470 1147.140 193.530 ;
        RECT 1146.480 193.390 1147.080 193.470 ;
        RECT 1146.480 159.110 1146.620 193.390 ;
        RECT 1146.420 158.790 1146.680 159.110 ;
        RECT 1146.880 158.110 1147.140 158.430 ;
        RECT 1146.940 111.365 1147.080 158.110 ;
        RECT 1146.870 110.995 1147.150 111.365 ;
        RECT 1146.870 89.915 1147.150 90.285 ;
        RECT 1146.940 89.750 1147.080 89.915 ;
        RECT 1146.880 89.430 1147.140 89.750 ;
        RECT 1145.960 41.490 1146.220 41.810 ;
        RECT 1146.020 24.470 1146.160 41.490 ;
        RECT 1145.960 24.150 1146.220 24.470 ;
        RECT 8.380 23.470 8.640 23.790 ;
        RECT 8.440 2.400 8.580 23.470 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 1146.870 1490.080 1147.150 1490.360 ;
        RECT 1147.790 1490.080 1148.070 1490.360 ;
        RECT 1146.410 1200.400 1146.690 1200.680 ;
        RECT 1147.790 1200.400 1148.070 1200.680 ;
        RECT 1146.410 1014.080 1146.690 1014.360 ;
        RECT 1147.790 1014.080 1148.070 1014.360 ;
        RECT 1146.410 917.520 1146.690 917.800 ;
        RECT 1147.790 917.520 1148.070 917.800 ;
        RECT 1146.410 724.400 1146.690 724.680 ;
        RECT 1147.790 724.400 1148.070 724.680 ;
        RECT 1146.410 627.840 1146.690 628.120 ;
        RECT 1147.790 627.840 1148.070 628.120 ;
        RECT 1146.870 111.040 1147.150 111.320 ;
        RECT 1146.870 89.960 1147.150 90.240 ;
      LAYER met3 ;
        RECT 1146.845 1490.370 1147.175 1490.385 ;
        RECT 1147.765 1490.370 1148.095 1490.385 ;
        RECT 1146.845 1490.070 1148.095 1490.370 ;
        RECT 1146.845 1490.055 1147.175 1490.070 ;
        RECT 1147.765 1490.055 1148.095 1490.070 ;
        RECT 1146.385 1200.690 1146.715 1200.705 ;
        RECT 1147.765 1200.690 1148.095 1200.705 ;
        RECT 1146.385 1200.390 1148.095 1200.690 ;
        RECT 1146.385 1200.375 1146.715 1200.390 ;
        RECT 1147.765 1200.375 1148.095 1200.390 ;
        RECT 1146.385 1014.370 1146.715 1014.385 ;
        RECT 1147.765 1014.370 1148.095 1014.385 ;
        RECT 1146.385 1014.070 1148.095 1014.370 ;
        RECT 1146.385 1014.055 1146.715 1014.070 ;
        RECT 1147.765 1014.055 1148.095 1014.070 ;
        RECT 1146.385 917.810 1146.715 917.825 ;
        RECT 1147.765 917.810 1148.095 917.825 ;
        RECT 1146.385 917.510 1148.095 917.810 ;
        RECT 1146.385 917.495 1146.715 917.510 ;
        RECT 1147.765 917.495 1148.095 917.510 ;
        RECT 1146.385 724.690 1146.715 724.705 ;
        RECT 1147.765 724.690 1148.095 724.705 ;
        RECT 1146.385 724.390 1148.095 724.690 ;
        RECT 1146.385 724.375 1146.715 724.390 ;
        RECT 1147.765 724.375 1148.095 724.390 ;
        RECT 1146.385 628.130 1146.715 628.145 ;
        RECT 1147.765 628.130 1148.095 628.145 ;
        RECT 1146.385 627.830 1148.095 628.130 ;
        RECT 1146.385 627.815 1146.715 627.830 ;
        RECT 1147.765 627.815 1148.095 627.830 ;
        RECT 1146.845 111.340 1147.175 111.345 ;
        RECT 1146.590 111.330 1147.175 111.340 ;
        RECT 1146.390 111.030 1147.175 111.330 ;
        RECT 1146.590 111.020 1147.175 111.030 ;
        RECT 1146.845 111.015 1147.175 111.020 ;
        RECT 1146.845 90.260 1147.175 90.265 ;
        RECT 1146.590 90.250 1147.175 90.260 ;
        RECT 1146.590 89.950 1147.400 90.250 ;
        RECT 1146.590 89.940 1147.175 89.950 ;
        RECT 1146.845 89.935 1147.175 89.940 ;
      LAYER via3 ;
        RECT 1146.620 111.020 1146.940 111.340 ;
        RECT 1146.620 89.940 1146.940 90.260 ;
      LAYER met4 ;
        RECT 1146.615 111.015 1146.945 111.345 ;
        RECT 1146.630 90.265 1146.930 111.015 ;
        RECT 1146.615 89.935 1146.945 90.265 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1121.165 23.885 1121.335 24.735 ;
      LAYER mcon ;
        RECT 1121.165 24.565 1121.335 24.735 ;
      LAYER met1 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 1121.105 24.720 1121.395 24.765 ;
        RECT 14.330 24.580 1121.395 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 1121.105 24.535 1121.395 24.580 ;
        RECT 1152.370 24.380 1152.690 24.440 ;
        RECT 1146.940 24.240 1152.690 24.380 ;
        RECT 1121.105 24.040 1121.395 24.085 ;
        RECT 1146.940 24.040 1147.080 24.240 ;
        RECT 1152.370 24.180 1152.690 24.240 ;
        RECT 1121.105 23.900 1147.080 24.040 ;
        RECT 1121.105 23.855 1121.395 23.900 ;
      LAYER via ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 1152.400 24.180 1152.660 24.440 ;
      LAYER met2 ;
        RECT 1154.165 1700.410 1154.445 1704.000 ;
        RECT 1152.460 1700.270 1154.445 1700.410 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 1152.460 24.470 1152.600 1700.270 ;
        RECT 1154.165 1700.000 1154.445 1700.270 ;
        RECT 1152.400 24.150 1152.660 24.470 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1159.730 1678.140 1160.050 1678.200 ;
        RECT 1162.030 1678.140 1162.350 1678.200 ;
        RECT 1159.730 1678.000 1162.350 1678.140 ;
        RECT 1159.730 1677.940 1160.050 1678.000 ;
        RECT 1162.030 1677.940 1162.350 1678.000 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1159.730 25.060 1160.050 25.120 ;
        RECT 38.250 24.920 1160.050 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1159.730 24.860 1160.050 24.920 ;
      LAYER via ;
        RECT 1159.760 1677.940 1160.020 1678.200 ;
        RECT 1162.060 1677.940 1162.320 1678.200 ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1159.760 24.860 1160.020 25.120 ;
      LAYER met2 ;
        RECT 1163.365 1700.410 1163.645 1704.000 ;
        RECT 1162.120 1700.270 1163.645 1700.410 ;
        RECT 1162.120 1678.230 1162.260 1700.270 ;
        RECT 1163.365 1700.000 1163.645 1700.270 ;
        RECT 1159.760 1677.910 1160.020 1678.230 ;
        RECT 1162.060 1677.910 1162.320 1678.230 ;
        RECT 1159.820 25.150 1159.960 1677.910 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 1159.760 24.830 1160.020 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1235.630 1678.140 1235.950 1678.200 ;
        RECT 1238.390 1678.140 1238.710 1678.200 ;
        RECT 1235.630 1678.000 1238.710 1678.140 ;
        RECT 1235.630 1677.940 1235.950 1678.000 ;
        RECT 1238.390 1677.940 1238.710 1678.000 ;
        RECT 240.650 25.740 240.970 25.800 ;
        RECT 1235.630 25.740 1235.950 25.800 ;
        RECT 240.650 25.600 1235.950 25.740 ;
        RECT 240.650 25.540 240.970 25.600 ;
        RECT 1235.630 25.540 1235.950 25.600 ;
      LAYER via ;
        RECT 1235.660 1677.940 1235.920 1678.200 ;
        RECT 1238.420 1677.940 1238.680 1678.200 ;
        RECT 240.680 25.540 240.940 25.800 ;
        RECT 1235.660 25.540 1235.920 25.800 ;
      LAYER met2 ;
        RECT 1239.725 1700.410 1240.005 1704.000 ;
        RECT 1238.480 1700.270 1240.005 1700.410 ;
        RECT 1238.480 1678.230 1238.620 1700.270 ;
        RECT 1239.725 1700.000 1240.005 1700.270 ;
        RECT 1235.660 1677.910 1235.920 1678.230 ;
        RECT 1238.420 1677.910 1238.680 1678.230 ;
        RECT 1235.720 25.830 1235.860 1677.910 ;
        RECT 240.680 25.510 240.940 25.830 ;
        RECT 1235.660 25.510 1235.920 25.830 ;
        RECT 240.740 2.400 240.880 25.510 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1243.985 1497.445 1244.155 1559.835 ;
        RECT 1243.525 427.805 1243.695 473.195 ;
        RECT 1243.985 331.245 1244.155 379.355 ;
      LAYER mcon ;
        RECT 1243.985 1559.665 1244.155 1559.835 ;
        RECT 1243.525 473.025 1243.695 473.195 ;
        RECT 1243.985 379.185 1244.155 379.355 ;
      LAYER met1 ;
        RECT 1244.370 1628.500 1244.690 1628.560 ;
        RECT 1246.210 1628.500 1246.530 1628.560 ;
        RECT 1244.370 1628.360 1246.530 1628.500 ;
        RECT 1244.370 1628.300 1244.690 1628.360 ;
        RECT 1246.210 1628.300 1246.530 1628.360 ;
        RECT 1243.910 1611.160 1244.230 1611.220 ;
        RECT 1246.210 1611.160 1246.530 1611.220 ;
        RECT 1243.910 1611.020 1246.530 1611.160 ;
        RECT 1243.910 1610.960 1244.230 1611.020 ;
        RECT 1246.210 1610.960 1246.530 1611.020 ;
        RECT 1243.925 1559.820 1244.215 1559.865 ;
        RECT 1244.370 1559.820 1244.690 1559.880 ;
        RECT 1243.925 1559.680 1244.690 1559.820 ;
        RECT 1243.925 1559.635 1244.215 1559.680 ;
        RECT 1244.370 1559.620 1244.690 1559.680 ;
        RECT 1243.910 1497.600 1244.230 1497.660 ;
        RECT 1243.715 1497.460 1244.230 1497.600 ;
        RECT 1243.910 1497.400 1244.230 1497.460 ;
        RECT 1243.910 883.900 1244.230 883.960 ;
        RECT 1243.540 883.760 1244.230 883.900 ;
        RECT 1243.540 883.280 1243.680 883.760 ;
        RECT 1243.910 883.700 1244.230 883.760 ;
        RECT 1243.450 883.020 1243.770 883.280 ;
        RECT 1243.450 473.180 1243.770 473.240 ;
        RECT 1243.255 473.040 1243.770 473.180 ;
        RECT 1243.450 472.980 1243.770 473.040 ;
        RECT 1243.465 427.960 1243.755 428.005 ;
        RECT 1243.910 427.960 1244.230 428.020 ;
        RECT 1243.465 427.820 1244.230 427.960 ;
        RECT 1243.465 427.775 1243.755 427.820 ;
        RECT 1243.910 427.760 1244.230 427.820 ;
        RECT 1243.910 379.340 1244.230 379.400 ;
        RECT 1243.715 379.200 1244.230 379.340 ;
        RECT 1243.910 379.140 1244.230 379.200 ;
        RECT 1243.910 331.400 1244.230 331.460 ;
        RECT 1243.715 331.260 1244.230 331.400 ;
        RECT 1243.910 331.200 1244.230 331.260 ;
        RECT 1243.910 97.140 1244.230 97.200 ;
        RECT 1243.540 97.000 1244.230 97.140 ;
        RECT 1243.540 96.860 1243.680 97.000 ;
        RECT 1243.910 96.940 1244.230 97.000 ;
        RECT 1243.450 96.600 1243.770 96.860 ;
        RECT 258.130 26.080 258.450 26.140 ;
        RECT 1243.450 26.080 1243.770 26.140 ;
        RECT 258.130 25.940 1243.770 26.080 ;
        RECT 258.130 25.880 258.450 25.940 ;
        RECT 1243.450 25.880 1243.770 25.940 ;
      LAYER via ;
        RECT 1244.400 1628.300 1244.660 1628.560 ;
        RECT 1246.240 1628.300 1246.500 1628.560 ;
        RECT 1243.940 1610.960 1244.200 1611.220 ;
        RECT 1246.240 1610.960 1246.500 1611.220 ;
        RECT 1244.400 1559.620 1244.660 1559.880 ;
        RECT 1243.940 1497.400 1244.200 1497.660 ;
        RECT 1243.940 883.700 1244.200 883.960 ;
        RECT 1243.480 883.020 1243.740 883.280 ;
        RECT 1243.480 472.980 1243.740 473.240 ;
        RECT 1243.940 427.760 1244.200 428.020 ;
        RECT 1243.940 379.140 1244.200 379.400 ;
        RECT 1243.940 331.200 1244.200 331.460 ;
        RECT 1243.940 96.940 1244.200 97.200 ;
        RECT 1243.480 96.600 1243.740 96.860 ;
        RECT 258.160 25.880 258.420 26.140 ;
        RECT 1243.480 25.880 1243.740 26.140 ;
      LAYER met2 ;
        RECT 1246.165 1700.410 1246.445 1704.000 ;
        RECT 1244.460 1700.270 1246.445 1700.410 ;
        RECT 1244.460 1628.590 1244.600 1700.270 ;
        RECT 1246.165 1700.000 1246.445 1700.270 ;
        RECT 1244.400 1628.270 1244.660 1628.590 ;
        RECT 1246.240 1628.270 1246.500 1628.590 ;
        RECT 1246.300 1611.250 1246.440 1628.270 ;
        RECT 1243.940 1610.930 1244.200 1611.250 ;
        RECT 1246.240 1610.930 1246.500 1611.250 ;
        RECT 1244.000 1587.530 1244.140 1610.930 ;
        RECT 1244.000 1587.390 1244.600 1587.530 ;
        RECT 1244.460 1559.910 1244.600 1587.390 ;
        RECT 1244.400 1559.590 1244.660 1559.910 ;
        RECT 1243.940 1497.370 1244.200 1497.690 ;
        RECT 1244.000 1486.890 1244.140 1497.370 ;
        RECT 1243.540 1486.750 1244.140 1486.890 ;
        RECT 1243.540 1438.610 1243.680 1486.750 ;
        RECT 1243.540 1438.470 1244.140 1438.610 ;
        RECT 1244.000 1388.970 1244.140 1438.470 ;
        RECT 1243.540 1388.830 1244.140 1388.970 ;
        RECT 1243.540 1352.930 1243.680 1388.830 ;
        RECT 1243.540 1352.790 1244.140 1352.930 ;
        RECT 1244.000 1292.410 1244.140 1352.790 ;
        RECT 1243.540 1292.270 1244.140 1292.410 ;
        RECT 1243.540 1256.370 1243.680 1292.270 ;
        RECT 1243.540 1256.230 1244.140 1256.370 ;
        RECT 1244.000 1197.210 1244.140 1256.230 ;
        RECT 1243.540 1197.070 1244.140 1197.210 ;
        RECT 1243.540 1148.930 1243.680 1197.070 ;
        RECT 1243.540 1148.790 1244.140 1148.930 ;
        RECT 1244.000 1089.770 1244.140 1148.790 ;
        RECT 1243.540 1089.630 1244.140 1089.770 ;
        RECT 1243.540 1053.730 1243.680 1089.630 ;
        RECT 1243.540 1053.590 1244.140 1053.730 ;
        RECT 1244.000 993.210 1244.140 1053.590 ;
        RECT 1243.540 993.070 1244.140 993.210 ;
        RECT 1243.540 957.170 1243.680 993.070 ;
        RECT 1243.540 957.030 1244.140 957.170 ;
        RECT 1244.000 883.990 1244.140 957.030 ;
        RECT 1243.940 883.670 1244.200 883.990 ;
        RECT 1243.480 882.990 1243.740 883.310 ;
        RECT 1243.540 859.250 1243.680 882.990 ;
        RECT 1243.540 859.110 1244.140 859.250 ;
        RECT 1244.000 810.970 1244.140 859.110 ;
        RECT 1243.540 810.830 1244.140 810.970 ;
        RECT 1243.540 762.690 1243.680 810.830 ;
        RECT 1243.540 762.550 1244.140 762.690 ;
        RECT 1244.000 617.850 1244.140 762.550 ;
        RECT 1243.540 617.710 1244.140 617.850 ;
        RECT 1243.540 569.570 1243.680 617.710 ;
        RECT 1243.540 569.430 1244.140 569.570 ;
        RECT 1244.000 521.290 1244.140 569.430 ;
        RECT 1243.540 521.150 1244.140 521.290 ;
        RECT 1243.540 473.270 1243.680 521.150 ;
        RECT 1243.480 472.950 1243.740 473.270 ;
        RECT 1243.940 427.730 1244.200 428.050 ;
        RECT 1244.000 379.430 1244.140 427.730 ;
        RECT 1243.940 379.110 1244.200 379.430 ;
        RECT 1243.940 331.170 1244.200 331.490 ;
        RECT 1244.000 313.890 1244.140 331.170 ;
        RECT 1243.540 313.750 1244.140 313.890 ;
        RECT 1243.540 279.210 1243.680 313.750 ;
        RECT 1243.540 279.070 1244.140 279.210 ;
        RECT 1244.000 97.230 1244.140 279.070 ;
        RECT 1243.940 96.910 1244.200 97.230 ;
        RECT 1243.480 96.570 1243.740 96.890 ;
        RECT 1243.540 26.170 1243.680 96.570 ;
        RECT 258.160 25.850 258.420 26.170 ;
        RECT 1243.480 25.850 1243.740 26.170 ;
        RECT 258.220 2.400 258.360 25.850 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1250.425 1497.445 1250.595 1579.895 ;
      LAYER mcon ;
        RECT 1250.425 1579.725 1250.595 1579.895 ;
      LAYER met1 ;
        RECT 1249.890 1580.560 1250.210 1580.620 ;
        RECT 1250.810 1580.560 1251.130 1580.620 ;
        RECT 1249.890 1580.420 1251.130 1580.560 ;
        RECT 1249.890 1580.360 1250.210 1580.420 ;
        RECT 1250.810 1580.360 1251.130 1580.420 ;
        RECT 1250.365 1579.880 1250.655 1579.925 ;
        RECT 1250.810 1579.880 1251.130 1579.940 ;
        RECT 1250.365 1579.740 1251.130 1579.880 ;
        RECT 1250.365 1579.695 1250.655 1579.740 ;
        RECT 1250.810 1579.680 1251.130 1579.740 ;
        RECT 1250.350 1497.600 1250.670 1497.660 ;
        RECT 1250.155 1497.460 1250.670 1497.600 ;
        RECT 1250.350 1497.400 1250.670 1497.460 ;
        RECT 1249.890 283.120 1250.210 283.180 ;
        RECT 1250.350 283.120 1250.670 283.180 ;
        RECT 1249.890 282.980 1250.670 283.120 ;
        RECT 1249.890 282.920 1250.210 282.980 ;
        RECT 1250.350 282.920 1250.670 282.980 ;
        RECT 1249.890 96.800 1250.210 96.860 ;
        RECT 1250.350 96.800 1250.670 96.860 ;
        RECT 1249.890 96.660 1250.670 96.800 ;
        RECT 1249.890 96.600 1250.210 96.660 ;
        RECT 1250.350 96.600 1250.670 96.660 ;
      LAYER via ;
        RECT 1249.920 1580.360 1250.180 1580.620 ;
        RECT 1250.840 1580.360 1251.100 1580.620 ;
        RECT 1250.840 1579.680 1251.100 1579.940 ;
        RECT 1250.380 1497.400 1250.640 1497.660 ;
        RECT 1249.920 282.920 1250.180 283.180 ;
        RECT 1250.380 282.920 1250.640 283.180 ;
        RECT 1249.920 96.600 1250.180 96.860 ;
        RECT 1250.380 96.600 1250.640 96.860 ;
      LAYER met2 ;
        RECT 1253.065 1700.410 1253.345 1704.000 ;
        RECT 1251.360 1700.270 1253.345 1700.410 ;
        RECT 1251.360 1677.970 1251.500 1700.270 ;
        RECT 1253.065 1700.000 1253.345 1700.270 ;
        RECT 1250.900 1677.830 1251.500 1677.970 ;
        RECT 1250.900 1676.725 1251.040 1677.830 ;
        RECT 1250.830 1676.355 1251.110 1676.725 ;
        RECT 1251.290 1675.675 1251.570 1676.045 ;
        RECT 1251.360 1628.445 1251.500 1675.675 ;
        RECT 1249.910 1628.075 1250.190 1628.445 ;
        RECT 1251.290 1628.075 1251.570 1628.445 ;
        RECT 1249.980 1580.650 1250.120 1628.075 ;
        RECT 1249.920 1580.330 1250.180 1580.650 ;
        RECT 1250.840 1580.330 1251.100 1580.650 ;
        RECT 1250.900 1579.970 1251.040 1580.330 ;
        RECT 1250.840 1579.650 1251.100 1579.970 ;
        RECT 1250.380 1497.370 1250.640 1497.690 ;
        RECT 1250.440 1486.890 1250.580 1497.370 ;
        RECT 1249.980 1486.750 1250.580 1486.890 ;
        RECT 1249.980 1438.610 1250.120 1486.750 ;
        RECT 1249.980 1438.470 1250.580 1438.610 ;
        RECT 1250.440 1388.970 1250.580 1438.470 ;
        RECT 1249.980 1388.830 1250.580 1388.970 ;
        RECT 1249.980 1352.930 1250.120 1388.830 ;
        RECT 1249.980 1352.790 1250.580 1352.930 ;
        RECT 1250.440 1292.410 1250.580 1352.790 ;
        RECT 1249.980 1292.270 1250.580 1292.410 ;
        RECT 1249.980 1256.370 1250.120 1292.270 ;
        RECT 1249.980 1256.230 1250.580 1256.370 ;
        RECT 1250.440 1197.210 1250.580 1256.230 ;
        RECT 1249.980 1197.070 1250.580 1197.210 ;
        RECT 1249.980 1148.930 1250.120 1197.070 ;
        RECT 1249.980 1148.790 1250.580 1148.930 ;
        RECT 1250.440 1089.770 1250.580 1148.790 ;
        RECT 1249.980 1089.630 1250.580 1089.770 ;
        RECT 1249.980 1053.730 1250.120 1089.630 ;
        RECT 1249.980 1053.590 1250.580 1053.730 ;
        RECT 1250.440 993.210 1250.580 1053.590 ;
        RECT 1249.980 993.070 1250.580 993.210 ;
        RECT 1249.980 957.170 1250.120 993.070 ;
        RECT 1249.980 957.030 1250.580 957.170 ;
        RECT 1250.440 893.930 1250.580 957.030 ;
        RECT 1249.980 893.790 1250.580 893.930 ;
        RECT 1249.980 859.250 1250.120 893.790 ;
        RECT 1249.980 859.110 1250.580 859.250 ;
        RECT 1250.440 810.970 1250.580 859.110 ;
        RECT 1249.980 810.830 1250.580 810.970 ;
        RECT 1249.980 762.690 1250.120 810.830 ;
        RECT 1249.980 762.550 1250.580 762.690 ;
        RECT 1250.440 617.850 1250.580 762.550 ;
        RECT 1249.980 617.710 1250.580 617.850 ;
        RECT 1249.980 569.570 1250.120 617.710 ;
        RECT 1249.980 569.430 1250.580 569.570 ;
        RECT 1250.440 521.290 1250.580 569.430 ;
        RECT 1249.980 521.150 1250.580 521.290 ;
        RECT 1249.980 473.010 1250.120 521.150 ;
        RECT 1249.980 472.870 1250.580 473.010 ;
        RECT 1250.440 283.210 1250.580 472.870 ;
        RECT 1249.920 282.890 1250.180 283.210 ;
        RECT 1250.380 282.890 1250.640 283.210 ;
        RECT 1249.980 279.210 1250.120 282.890 ;
        RECT 1249.980 279.070 1250.580 279.210 ;
        RECT 1250.440 96.890 1250.580 279.070 ;
        RECT 1249.920 96.570 1250.180 96.890 ;
        RECT 1250.380 96.570 1250.640 96.890 ;
        RECT 1249.980 31.125 1250.120 96.570 ;
        RECT 276.090 30.755 276.370 31.125 ;
        RECT 1249.910 30.755 1250.190 31.125 ;
        RECT 276.160 2.400 276.300 30.755 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 1250.830 1676.400 1251.110 1676.680 ;
        RECT 1251.290 1675.720 1251.570 1676.000 ;
        RECT 1249.910 1628.120 1250.190 1628.400 ;
        RECT 1251.290 1628.120 1251.570 1628.400 ;
        RECT 276.090 30.800 276.370 31.080 ;
        RECT 1249.910 30.800 1250.190 31.080 ;
      LAYER met3 ;
        RECT 1250.805 1676.690 1251.135 1676.705 ;
        RECT 1250.590 1676.375 1251.135 1676.690 ;
        RECT 1250.590 1676.010 1250.890 1676.375 ;
        RECT 1251.265 1676.010 1251.595 1676.025 ;
        RECT 1250.590 1675.710 1251.595 1676.010 ;
        RECT 1251.265 1675.695 1251.595 1675.710 ;
        RECT 1249.885 1628.410 1250.215 1628.425 ;
        RECT 1251.265 1628.410 1251.595 1628.425 ;
        RECT 1249.885 1628.110 1251.595 1628.410 ;
        RECT 1249.885 1628.095 1250.215 1628.110 ;
        RECT 1251.265 1628.095 1251.595 1628.110 ;
        RECT 276.065 31.090 276.395 31.105 ;
        RECT 1249.885 31.090 1250.215 31.105 ;
        RECT 276.065 30.790 1250.215 31.090 ;
        RECT 276.065 30.775 276.395 30.790 ;
        RECT 1249.885 30.775 1250.215 30.790 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1257.325 1304.325 1257.495 1369.435 ;
        RECT 1257.325 1255.365 1257.495 1297.015 ;
        RECT 1257.325 1200.625 1257.495 1207.595 ;
        RECT 1257.325 1152.345 1257.495 1200.115 ;
        RECT 1256.865 807.245 1257.035 855.355 ;
        RECT 1257.785 676.005 1257.955 717.655 ;
        RECT 1257.325 620.925 1257.495 669.375 ;
        RECT 1257.325 476.425 1257.495 524.195 ;
        RECT 1256.865 89.845 1257.035 137.955 ;
      LAYER mcon ;
        RECT 1257.325 1369.265 1257.495 1369.435 ;
        RECT 1257.325 1296.845 1257.495 1297.015 ;
        RECT 1257.325 1207.425 1257.495 1207.595 ;
        RECT 1257.325 1199.945 1257.495 1200.115 ;
        RECT 1256.865 855.185 1257.035 855.355 ;
        RECT 1257.785 717.485 1257.955 717.655 ;
        RECT 1257.325 669.205 1257.495 669.375 ;
        RECT 1257.325 524.025 1257.495 524.195 ;
        RECT 1256.865 137.785 1257.035 137.955 ;
      LAYER met1 ;
        RECT 1257.250 1642.100 1257.570 1642.160 ;
        RECT 1258.170 1642.100 1258.490 1642.160 ;
        RECT 1257.250 1641.960 1258.490 1642.100 ;
        RECT 1257.250 1641.900 1257.570 1641.960 ;
        RECT 1258.170 1641.900 1258.490 1641.960 ;
        RECT 1258.170 1594.500 1258.490 1594.560 ;
        RECT 1257.340 1594.360 1258.490 1594.500 ;
        RECT 1257.340 1593.880 1257.480 1594.360 ;
        RECT 1258.170 1594.300 1258.490 1594.360 ;
        RECT 1257.250 1593.620 1257.570 1593.880 ;
        RECT 1255.870 1393.900 1256.190 1393.960 ;
        RECT 1257.250 1393.900 1257.570 1393.960 ;
        RECT 1255.870 1393.760 1257.570 1393.900 ;
        RECT 1255.870 1393.700 1256.190 1393.760 ;
        RECT 1257.250 1393.700 1257.570 1393.760 ;
        RECT 1257.250 1369.420 1257.570 1369.480 ;
        RECT 1257.055 1369.280 1257.570 1369.420 ;
        RECT 1257.250 1369.220 1257.570 1369.280 ;
        RECT 1257.250 1304.480 1257.570 1304.540 ;
        RECT 1257.055 1304.340 1257.570 1304.480 ;
        RECT 1257.250 1304.280 1257.570 1304.340 ;
        RECT 1257.250 1297.000 1257.570 1297.060 ;
        RECT 1257.055 1296.860 1257.570 1297.000 ;
        RECT 1257.250 1296.800 1257.570 1296.860 ;
        RECT 1257.265 1255.520 1257.555 1255.565 ;
        RECT 1257.710 1255.520 1258.030 1255.580 ;
        RECT 1257.265 1255.380 1258.030 1255.520 ;
        RECT 1257.265 1255.335 1257.555 1255.380 ;
        RECT 1257.710 1255.320 1258.030 1255.380 ;
        RECT 1257.250 1207.580 1257.570 1207.640 ;
        RECT 1257.055 1207.440 1257.570 1207.580 ;
        RECT 1257.250 1207.380 1257.570 1207.440 ;
        RECT 1257.250 1200.780 1257.570 1200.840 ;
        RECT 1257.055 1200.640 1257.570 1200.780 ;
        RECT 1257.250 1200.580 1257.570 1200.640 ;
        RECT 1257.250 1200.100 1257.570 1200.160 ;
        RECT 1257.055 1199.960 1257.570 1200.100 ;
        RECT 1257.250 1199.900 1257.570 1199.960 ;
        RECT 1257.250 1152.500 1257.570 1152.560 ;
        RECT 1257.055 1152.360 1257.570 1152.500 ;
        RECT 1257.250 1152.300 1257.570 1152.360 ;
        RECT 1255.870 1121.220 1256.190 1121.280 ;
        RECT 1257.250 1121.220 1257.570 1121.280 ;
        RECT 1255.870 1121.080 1257.570 1121.220 ;
        RECT 1255.870 1121.020 1256.190 1121.080 ;
        RECT 1257.250 1121.020 1257.570 1121.080 ;
        RECT 1256.790 1048.800 1257.110 1048.860 ;
        RECT 1258.630 1048.800 1258.950 1048.860 ;
        RECT 1256.790 1048.660 1258.950 1048.800 ;
        RECT 1256.790 1048.600 1257.110 1048.660 ;
        RECT 1258.630 1048.600 1258.950 1048.660 ;
        RECT 1257.250 959.380 1257.570 959.440 ;
        RECT 1257.710 959.380 1258.030 959.440 ;
        RECT 1257.250 959.240 1258.030 959.380 ;
        RECT 1257.250 959.180 1257.570 959.240 ;
        RECT 1257.710 959.180 1258.030 959.240 ;
        RECT 1256.790 862.480 1257.110 862.540 ;
        RECT 1257.250 862.480 1257.570 862.540 ;
        RECT 1256.790 862.340 1257.570 862.480 ;
        RECT 1256.790 862.280 1257.110 862.340 ;
        RECT 1257.250 862.280 1257.570 862.340 ;
        RECT 1256.790 855.340 1257.110 855.400 ;
        RECT 1256.595 855.200 1257.110 855.340 ;
        RECT 1256.790 855.140 1257.110 855.200 ;
        RECT 1256.805 807.400 1257.095 807.445 ;
        RECT 1257.250 807.400 1257.570 807.460 ;
        RECT 1256.805 807.260 1257.570 807.400 ;
        RECT 1256.805 807.215 1257.095 807.260 ;
        RECT 1257.250 807.200 1257.570 807.260 ;
        RECT 1255.870 759.120 1256.190 759.180 ;
        RECT 1256.790 759.120 1257.110 759.180 ;
        RECT 1255.870 758.980 1257.110 759.120 ;
        RECT 1255.870 758.920 1256.190 758.980 ;
        RECT 1256.790 758.920 1257.110 758.980 ;
        RECT 1256.790 717.640 1257.110 717.700 ;
        RECT 1257.725 717.640 1258.015 717.685 ;
        RECT 1256.790 717.500 1258.015 717.640 ;
        RECT 1256.790 717.440 1257.110 717.500 ;
        RECT 1257.725 717.455 1258.015 717.500 ;
        RECT 1257.710 676.160 1258.030 676.220 ;
        RECT 1257.515 676.020 1258.030 676.160 ;
        RECT 1257.710 675.960 1258.030 676.020 ;
        RECT 1257.265 669.360 1257.555 669.405 ;
        RECT 1257.710 669.360 1258.030 669.420 ;
        RECT 1257.265 669.220 1258.030 669.360 ;
        RECT 1257.265 669.175 1257.555 669.220 ;
        RECT 1257.710 669.160 1258.030 669.220 ;
        RECT 1257.250 621.080 1257.570 621.140 ;
        RECT 1257.055 620.940 1257.570 621.080 ;
        RECT 1257.250 620.880 1257.570 620.940 ;
        RECT 1257.250 524.180 1257.570 524.240 ;
        RECT 1257.055 524.040 1257.570 524.180 ;
        RECT 1257.250 523.980 1257.570 524.040 ;
        RECT 1257.250 476.580 1257.570 476.640 ;
        RECT 1257.055 476.440 1257.570 476.580 ;
        RECT 1257.250 476.380 1257.570 476.440 ;
        RECT 1255.870 475.900 1256.190 475.960 ;
        RECT 1257.250 475.900 1257.570 475.960 ;
        RECT 1255.870 475.760 1257.570 475.900 ;
        RECT 1255.870 475.700 1256.190 475.760 ;
        RECT 1257.250 475.700 1257.570 475.760 ;
        RECT 1256.790 234.500 1257.110 234.560 ;
        RECT 1257.250 234.500 1257.570 234.560 ;
        RECT 1256.790 234.360 1257.570 234.500 ;
        RECT 1256.790 234.300 1257.110 234.360 ;
        RECT 1257.250 234.300 1257.570 234.360 ;
        RECT 1256.805 137.940 1257.095 137.985 ;
        RECT 1257.250 137.940 1257.570 138.000 ;
        RECT 1256.805 137.800 1257.570 137.940 ;
        RECT 1256.805 137.755 1257.095 137.800 ;
        RECT 1257.250 137.740 1257.570 137.800 ;
        RECT 1256.805 89.815 1257.095 90.045 ;
        RECT 1256.880 89.660 1257.020 89.815 ;
        RECT 1257.710 89.660 1258.030 89.720 ;
        RECT 1256.880 89.520 1258.030 89.660 ;
        RECT 1257.710 89.460 1258.030 89.520 ;
        RECT 294.010 30.840 294.330 30.900 ;
        RECT 1256.330 30.840 1256.650 30.900 ;
        RECT 294.010 30.700 1256.650 30.840 ;
        RECT 294.010 30.640 294.330 30.700 ;
        RECT 1256.330 30.640 1256.650 30.700 ;
      LAYER via ;
        RECT 1257.280 1641.900 1257.540 1642.160 ;
        RECT 1258.200 1641.900 1258.460 1642.160 ;
        RECT 1258.200 1594.300 1258.460 1594.560 ;
        RECT 1257.280 1593.620 1257.540 1593.880 ;
        RECT 1255.900 1393.700 1256.160 1393.960 ;
        RECT 1257.280 1393.700 1257.540 1393.960 ;
        RECT 1257.280 1369.220 1257.540 1369.480 ;
        RECT 1257.280 1304.280 1257.540 1304.540 ;
        RECT 1257.280 1296.800 1257.540 1297.060 ;
        RECT 1257.740 1255.320 1258.000 1255.580 ;
        RECT 1257.280 1207.380 1257.540 1207.640 ;
        RECT 1257.280 1200.580 1257.540 1200.840 ;
        RECT 1257.280 1199.900 1257.540 1200.160 ;
        RECT 1257.280 1152.300 1257.540 1152.560 ;
        RECT 1255.900 1121.020 1256.160 1121.280 ;
        RECT 1257.280 1121.020 1257.540 1121.280 ;
        RECT 1256.820 1048.600 1257.080 1048.860 ;
        RECT 1258.660 1048.600 1258.920 1048.860 ;
        RECT 1257.280 959.180 1257.540 959.440 ;
        RECT 1257.740 959.180 1258.000 959.440 ;
        RECT 1256.820 862.280 1257.080 862.540 ;
        RECT 1257.280 862.280 1257.540 862.540 ;
        RECT 1256.820 855.140 1257.080 855.400 ;
        RECT 1257.280 807.200 1257.540 807.460 ;
        RECT 1255.900 758.920 1256.160 759.180 ;
        RECT 1256.820 758.920 1257.080 759.180 ;
        RECT 1256.820 717.440 1257.080 717.700 ;
        RECT 1257.740 675.960 1258.000 676.220 ;
        RECT 1257.740 669.160 1258.000 669.420 ;
        RECT 1257.280 620.880 1257.540 621.140 ;
        RECT 1257.280 523.980 1257.540 524.240 ;
        RECT 1257.280 476.380 1257.540 476.640 ;
        RECT 1255.900 475.700 1256.160 475.960 ;
        RECT 1257.280 475.700 1257.540 475.960 ;
        RECT 1256.820 234.300 1257.080 234.560 ;
        RECT 1257.280 234.300 1257.540 234.560 ;
        RECT 1257.280 137.740 1257.540 138.000 ;
        RECT 1257.740 89.460 1258.000 89.720 ;
        RECT 294.040 30.640 294.300 30.900 ;
        RECT 1256.360 30.640 1256.620 30.900 ;
      LAYER met2 ;
        RECT 1259.965 1700.410 1260.245 1704.000 ;
        RECT 1258.260 1700.270 1260.245 1700.410 ;
        RECT 1258.260 1677.970 1258.400 1700.270 ;
        RECT 1259.965 1700.000 1260.245 1700.270 ;
        RECT 1257.340 1677.830 1258.400 1677.970 ;
        RECT 1257.340 1642.190 1257.480 1677.830 ;
        RECT 1257.280 1641.870 1257.540 1642.190 ;
        RECT 1258.200 1641.870 1258.460 1642.190 ;
        RECT 1258.260 1594.590 1258.400 1641.870 ;
        RECT 1258.200 1594.270 1258.460 1594.590 ;
        RECT 1257.280 1593.590 1257.540 1593.910 ;
        RECT 1255.890 1441.755 1256.170 1442.125 ;
        RECT 1256.810 1442.010 1257.090 1442.125 ;
        RECT 1257.340 1442.010 1257.480 1593.590 ;
        RECT 1256.810 1441.870 1257.480 1442.010 ;
        RECT 1256.810 1441.755 1257.090 1441.870 ;
        RECT 1255.960 1393.990 1256.100 1441.755 ;
        RECT 1255.900 1393.670 1256.160 1393.990 ;
        RECT 1257.280 1393.670 1257.540 1393.990 ;
        RECT 1257.340 1369.510 1257.480 1393.670 ;
        RECT 1257.280 1369.190 1257.540 1369.510 ;
        RECT 1257.280 1304.250 1257.540 1304.570 ;
        RECT 1257.340 1297.090 1257.480 1304.250 ;
        RECT 1257.280 1296.770 1257.540 1297.090 ;
        RECT 1257.740 1255.290 1258.000 1255.610 ;
        RECT 1257.800 1248.890 1257.940 1255.290 ;
        RECT 1257.340 1248.750 1257.940 1248.890 ;
        RECT 1257.340 1207.670 1257.480 1248.750 ;
        RECT 1257.280 1207.350 1257.540 1207.670 ;
        RECT 1257.280 1200.550 1257.540 1200.870 ;
        RECT 1257.340 1200.190 1257.480 1200.550 ;
        RECT 1257.280 1199.870 1257.540 1200.190 ;
        RECT 1257.280 1152.270 1257.540 1152.590 ;
        RECT 1257.340 1121.310 1257.480 1152.270 ;
        RECT 1255.900 1120.990 1256.160 1121.310 ;
        RECT 1257.280 1120.990 1257.540 1121.310 ;
        RECT 1255.960 1097.365 1256.100 1120.990 ;
        RECT 1255.890 1096.995 1256.170 1097.365 ;
        RECT 1256.810 1096.995 1257.090 1097.365 ;
        RECT 1256.880 1048.890 1257.020 1096.995 ;
        RECT 1256.820 1048.570 1257.080 1048.890 ;
        RECT 1258.660 1048.570 1258.920 1048.890 ;
        RECT 1258.720 1000.805 1258.860 1048.570 ;
        RECT 1257.730 1000.435 1258.010 1000.805 ;
        RECT 1258.650 1000.435 1258.930 1000.805 ;
        RECT 1257.800 959.470 1257.940 1000.435 ;
        RECT 1257.280 959.150 1257.540 959.470 ;
        RECT 1257.740 959.150 1258.000 959.470 ;
        RECT 1257.340 911.725 1257.480 959.150 ;
        RECT 1257.270 911.355 1257.550 911.725 ;
        RECT 1258.190 909.995 1258.470 910.365 ;
        RECT 1258.260 862.765 1258.400 909.995 ;
        RECT 1256.820 862.250 1257.080 862.570 ;
        RECT 1257.270 862.395 1257.550 862.765 ;
        RECT 1258.190 862.395 1258.470 862.765 ;
        RECT 1257.280 862.250 1257.540 862.395 ;
        RECT 1256.880 855.430 1257.020 862.250 ;
        RECT 1256.820 855.110 1257.080 855.430 ;
        RECT 1257.280 807.170 1257.540 807.490 ;
        RECT 1257.340 806.890 1257.480 807.170 ;
        RECT 1256.880 806.750 1257.480 806.890 ;
        RECT 1256.880 759.210 1257.020 806.750 ;
        RECT 1255.900 758.890 1256.160 759.210 ;
        RECT 1256.820 758.890 1257.080 759.210 ;
        RECT 1255.960 717.925 1256.100 758.890 ;
        RECT 1255.890 717.555 1256.170 717.925 ;
        RECT 1256.810 717.555 1257.090 717.925 ;
        RECT 1256.820 717.410 1257.080 717.555 ;
        RECT 1257.740 675.930 1258.000 676.250 ;
        RECT 1257.800 669.450 1257.940 675.930 ;
        RECT 1257.740 669.130 1258.000 669.450 ;
        RECT 1257.280 620.850 1257.540 621.170 ;
        RECT 1257.340 572.290 1257.480 620.850 ;
        RECT 1256.880 572.150 1257.480 572.290 ;
        RECT 1256.880 525.485 1257.020 572.150 ;
        RECT 1256.810 525.115 1257.090 525.485 ;
        RECT 1257.270 524.435 1257.550 524.805 ;
        RECT 1257.340 524.270 1257.480 524.435 ;
        RECT 1257.280 523.950 1257.540 524.270 ;
        RECT 1257.280 476.350 1257.540 476.670 ;
        RECT 1257.340 475.990 1257.480 476.350 ;
        RECT 1255.900 475.670 1256.160 475.990 ;
        RECT 1257.280 475.670 1257.540 475.990 ;
        RECT 1255.960 428.245 1256.100 475.670 ;
        RECT 1255.890 427.875 1256.170 428.245 ;
        RECT 1256.810 427.875 1257.090 428.245 ;
        RECT 1256.880 396.850 1257.020 427.875 ;
        RECT 1256.880 396.710 1257.480 396.850 ;
        RECT 1257.340 284.085 1257.480 396.710 ;
        RECT 1257.270 283.715 1257.550 284.085 ;
        RECT 1257.270 282.355 1257.550 282.725 ;
        RECT 1257.340 234.590 1257.480 282.355 ;
        RECT 1256.820 234.270 1257.080 234.590 ;
        RECT 1257.280 234.270 1257.540 234.590 ;
        RECT 1256.880 186.730 1257.020 234.270 ;
        RECT 1256.880 186.590 1257.480 186.730 ;
        RECT 1257.340 138.030 1257.480 186.590 ;
        RECT 1257.280 137.710 1257.540 138.030 ;
        RECT 1257.740 89.430 1258.000 89.750 ;
        RECT 1257.800 42.005 1257.940 89.430 ;
        RECT 1256.810 41.635 1257.090 42.005 ;
        RECT 1257.730 41.635 1258.010 42.005 ;
        RECT 1256.880 41.210 1257.020 41.635 ;
        RECT 1256.420 41.070 1257.020 41.210 ;
        RECT 1256.420 30.930 1256.560 41.070 ;
        RECT 294.040 30.610 294.300 30.930 ;
        RECT 1256.360 30.610 1256.620 30.930 ;
        RECT 294.100 2.400 294.240 30.610 ;
        RECT 293.890 -4.800 294.450 2.400 ;
      LAYER via2 ;
        RECT 1255.890 1441.800 1256.170 1442.080 ;
        RECT 1256.810 1441.800 1257.090 1442.080 ;
        RECT 1255.890 1097.040 1256.170 1097.320 ;
        RECT 1256.810 1097.040 1257.090 1097.320 ;
        RECT 1257.730 1000.480 1258.010 1000.760 ;
        RECT 1258.650 1000.480 1258.930 1000.760 ;
        RECT 1257.270 911.400 1257.550 911.680 ;
        RECT 1258.190 910.040 1258.470 910.320 ;
        RECT 1257.270 862.440 1257.550 862.720 ;
        RECT 1258.190 862.440 1258.470 862.720 ;
        RECT 1255.890 717.600 1256.170 717.880 ;
        RECT 1256.810 717.600 1257.090 717.880 ;
        RECT 1256.810 525.160 1257.090 525.440 ;
        RECT 1257.270 524.480 1257.550 524.760 ;
        RECT 1255.890 427.920 1256.170 428.200 ;
        RECT 1256.810 427.920 1257.090 428.200 ;
        RECT 1257.270 283.760 1257.550 284.040 ;
        RECT 1257.270 282.400 1257.550 282.680 ;
        RECT 1256.810 41.680 1257.090 41.960 ;
        RECT 1257.730 41.680 1258.010 41.960 ;
      LAYER met3 ;
        RECT 1255.865 1442.090 1256.195 1442.105 ;
        RECT 1256.785 1442.090 1257.115 1442.105 ;
        RECT 1255.865 1441.790 1257.115 1442.090 ;
        RECT 1255.865 1441.775 1256.195 1441.790 ;
        RECT 1256.785 1441.775 1257.115 1441.790 ;
        RECT 1255.865 1097.330 1256.195 1097.345 ;
        RECT 1256.785 1097.330 1257.115 1097.345 ;
        RECT 1255.865 1097.030 1257.115 1097.330 ;
        RECT 1255.865 1097.015 1256.195 1097.030 ;
        RECT 1256.785 1097.015 1257.115 1097.030 ;
        RECT 1257.705 1000.770 1258.035 1000.785 ;
        RECT 1258.625 1000.770 1258.955 1000.785 ;
        RECT 1257.705 1000.470 1258.955 1000.770 ;
        RECT 1257.705 1000.455 1258.035 1000.470 ;
        RECT 1258.625 1000.455 1258.955 1000.470 ;
        RECT 1257.245 911.690 1257.575 911.705 ;
        RECT 1257.030 911.375 1257.575 911.690 ;
        RECT 1257.030 910.330 1257.330 911.375 ;
        RECT 1258.165 910.330 1258.495 910.345 ;
        RECT 1257.030 910.030 1258.495 910.330 ;
        RECT 1258.165 910.015 1258.495 910.030 ;
        RECT 1257.245 862.730 1257.575 862.745 ;
        RECT 1258.165 862.730 1258.495 862.745 ;
        RECT 1257.245 862.430 1258.495 862.730 ;
        RECT 1257.245 862.415 1257.575 862.430 ;
        RECT 1258.165 862.415 1258.495 862.430 ;
        RECT 1255.865 717.890 1256.195 717.905 ;
        RECT 1256.785 717.890 1257.115 717.905 ;
        RECT 1255.865 717.590 1257.115 717.890 ;
        RECT 1255.865 717.575 1256.195 717.590 ;
        RECT 1256.785 717.575 1257.115 717.590 ;
        RECT 1256.785 525.450 1257.115 525.465 ;
        RECT 1256.785 525.150 1258.250 525.450 ;
        RECT 1256.785 525.135 1257.115 525.150 ;
        RECT 1257.245 524.770 1257.575 524.785 ;
        RECT 1257.950 524.770 1258.250 525.150 ;
        RECT 1257.245 524.470 1258.250 524.770 ;
        RECT 1257.245 524.455 1257.575 524.470 ;
        RECT 1255.865 428.210 1256.195 428.225 ;
        RECT 1256.785 428.210 1257.115 428.225 ;
        RECT 1255.865 427.910 1257.115 428.210 ;
        RECT 1255.865 427.895 1256.195 427.910 ;
        RECT 1256.785 427.895 1257.115 427.910 ;
        RECT 1257.245 284.050 1257.575 284.065 ;
        RECT 1257.030 283.735 1257.575 284.050 ;
        RECT 1257.030 282.705 1257.330 283.735 ;
        RECT 1257.030 282.390 1257.575 282.705 ;
        RECT 1257.245 282.375 1257.575 282.390 ;
        RECT 1256.785 41.970 1257.115 41.985 ;
        RECT 1257.705 41.970 1258.035 41.985 ;
        RECT 1256.785 41.670 1258.035 41.970 ;
        RECT 1256.785 41.655 1257.115 41.670 ;
        RECT 1257.705 41.655 1258.035 41.670 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1263.765 48.365 1263.935 113.815 ;
      LAYER mcon ;
        RECT 1263.765 113.645 1263.935 113.815 ;
      LAYER met1 ;
        RECT 1264.150 618.020 1264.470 618.080 ;
        RECT 1263.780 617.880 1264.470 618.020 ;
        RECT 1263.780 617.740 1263.920 617.880 ;
        RECT 1264.150 617.820 1264.470 617.880 ;
        RECT 1263.690 617.480 1264.010 617.740 ;
        RECT 1263.690 337.860 1264.010 337.920 ;
        RECT 1264.150 337.860 1264.470 337.920 ;
        RECT 1263.690 337.720 1264.470 337.860 ;
        RECT 1263.690 337.660 1264.010 337.720 ;
        RECT 1264.150 337.660 1264.470 337.720 ;
        RECT 1263.690 265.580 1264.010 265.840 ;
        RECT 1263.780 265.440 1263.920 265.580 ;
        RECT 1264.150 265.440 1264.470 265.500 ;
        RECT 1263.780 265.300 1264.470 265.440 ;
        RECT 1264.150 265.240 1264.470 265.300 ;
        RECT 1263.705 113.800 1263.995 113.845 ;
        RECT 1264.150 113.800 1264.470 113.860 ;
        RECT 1263.705 113.660 1264.470 113.800 ;
        RECT 1263.705 113.615 1263.995 113.660 ;
        RECT 1264.150 113.600 1264.470 113.660 ;
        RECT 1263.690 48.520 1264.010 48.580 ;
        RECT 1263.495 48.380 1264.010 48.520 ;
        RECT 1263.690 48.320 1264.010 48.380 ;
        RECT 311.950 31.180 312.270 31.240 ;
        RECT 1263.690 31.180 1264.010 31.240 ;
        RECT 311.950 31.040 1264.010 31.180 ;
        RECT 311.950 30.980 312.270 31.040 ;
        RECT 1263.690 30.980 1264.010 31.040 ;
      LAYER via ;
        RECT 1264.180 617.820 1264.440 618.080 ;
        RECT 1263.720 617.480 1263.980 617.740 ;
        RECT 1263.720 337.660 1263.980 337.920 ;
        RECT 1264.180 337.660 1264.440 337.920 ;
        RECT 1263.720 265.580 1263.980 265.840 ;
        RECT 1264.180 265.240 1264.440 265.500 ;
        RECT 1264.180 113.600 1264.440 113.860 ;
        RECT 1263.720 48.320 1263.980 48.580 ;
        RECT 311.980 30.980 312.240 31.240 ;
        RECT 1263.720 30.980 1263.980 31.240 ;
      LAYER met2 ;
        RECT 1266.405 1700.410 1266.685 1704.000 ;
        RECT 1264.700 1700.270 1266.685 1700.410 ;
        RECT 1264.700 1558.970 1264.840 1700.270 ;
        RECT 1266.405 1700.000 1266.685 1700.270 ;
        RECT 1264.240 1558.830 1264.840 1558.970 ;
        RECT 1264.240 1486.890 1264.380 1558.830 ;
        RECT 1263.780 1486.750 1264.380 1486.890 ;
        RECT 1263.780 1438.610 1263.920 1486.750 ;
        RECT 1263.780 1438.470 1264.380 1438.610 ;
        RECT 1264.240 1388.970 1264.380 1438.470 ;
        RECT 1263.780 1388.830 1264.380 1388.970 ;
        RECT 1263.780 1352.930 1263.920 1388.830 ;
        RECT 1263.780 1352.790 1264.380 1352.930 ;
        RECT 1264.240 1292.410 1264.380 1352.790 ;
        RECT 1263.780 1292.270 1264.380 1292.410 ;
        RECT 1263.780 1256.370 1263.920 1292.270 ;
        RECT 1263.780 1256.230 1264.380 1256.370 ;
        RECT 1264.240 1197.210 1264.380 1256.230 ;
        RECT 1263.780 1197.070 1264.380 1197.210 ;
        RECT 1263.780 1148.930 1263.920 1197.070 ;
        RECT 1263.780 1148.790 1264.380 1148.930 ;
        RECT 1264.240 1089.770 1264.380 1148.790 ;
        RECT 1263.780 1089.630 1264.380 1089.770 ;
        RECT 1263.780 1053.730 1263.920 1089.630 ;
        RECT 1263.780 1053.590 1264.380 1053.730 ;
        RECT 1264.240 993.210 1264.380 1053.590 ;
        RECT 1263.780 993.070 1264.380 993.210 ;
        RECT 1263.780 957.170 1263.920 993.070 ;
        RECT 1263.780 957.030 1264.380 957.170 ;
        RECT 1264.240 862.650 1264.380 957.030 ;
        RECT 1263.780 862.510 1264.380 862.650 ;
        RECT 1263.780 859.250 1263.920 862.510 ;
        RECT 1263.780 859.110 1264.380 859.250 ;
        RECT 1264.240 810.970 1264.380 859.110 ;
        RECT 1263.780 810.830 1264.380 810.970 ;
        RECT 1263.780 762.690 1263.920 810.830 ;
        RECT 1263.780 762.550 1264.380 762.690 ;
        RECT 1264.240 618.110 1264.380 762.550 ;
        RECT 1264.180 617.790 1264.440 618.110 ;
        RECT 1263.720 617.450 1263.980 617.770 ;
        RECT 1263.780 569.570 1263.920 617.450 ;
        RECT 1263.780 569.430 1264.380 569.570 ;
        RECT 1264.240 521.290 1264.380 569.430 ;
        RECT 1263.780 521.150 1264.380 521.290 ;
        RECT 1263.780 473.010 1263.920 521.150 ;
        RECT 1263.780 472.870 1264.380 473.010 ;
        RECT 1264.240 337.950 1264.380 472.870 ;
        RECT 1263.720 337.630 1263.980 337.950 ;
        RECT 1264.180 337.630 1264.440 337.950 ;
        RECT 1263.780 265.870 1263.920 337.630 ;
        RECT 1263.720 265.550 1263.980 265.870 ;
        RECT 1264.180 265.210 1264.440 265.530 ;
        RECT 1264.240 113.890 1264.380 265.210 ;
        RECT 1264.180 113.570 1264.440 113.890 ;
        RECT 1263.720 48.290 1263.980 48.610 ;
        RECT 1263.780 31.270 1263.920 48.290 ;
        RECT 311.980 30.950 312.240 31.270 ;
        RECT 1263.720 30.950 1263.980 31.270 ;
        RECT 312.040 2.400 312.180 30.950 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 31.520 330.210 31.580 ;
        RECT 1270.130 31.520 1270.450 31.580 ;
        RECT 329.890 31.380 1270.450 31.520 ;
        RECT 329.890 31.320 330.210 31.380 ;
        RECT 1270.130 31.320 1270.450 31.380 ;
      LAYER via ;
        RECT 329.920 31.320 330.180 31.580 ;
        RECT 1270.160 31.320 1270.420 31.580 ;
      LAYER met2 ;
        RECT 1273.305 1700.410 1273.585 1704.000 ;
        RECT 1271.600 1700.270 1273.585 1700.410 ;
        RECT 1271.600 1678.140 1271.740 1700.270 ;
        RECT 1273.305 1700.000 1273.585 1700.270 ;
        RECT 1270.220 1678.000 1271.740 1678.140 ;
        RECT 1270.220 31.610 1270.360 1678.000 ;
        RECT 329.920 31.290 330.180 31.610 ;
        RECT 1270.160 31.290 1270.420 31.610 ;
        RECT 329.980 2.400 330.120 31.290 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1278.025 1304.325 1278.195 1352.095 ;
        RECT 1278.025 1256.045 1278.195 1303.815 ;
        RECT 1278.025 931.345 1278.195 959.055 ;
        RECT 1278.025 862.665 1278.195 910.775 ;
        RECT 1278.025 524.365 1278.195 572.475 ;
        RECT 1278.485 469.285 1278.655 493.595 ;
        RECT 1278.485 421.005 1278.655 468.775 ;
        RECT 1278.025 323.425 1278.195 331.075 ;
        RECT 1278.025 228.225 1278.195 275.995 ;
      LAYER mcon ;
        RECT 1278.025 1351.925 1278.195 1352.095 ;
        RECT 1278.025 1303.645 1278.195 1303.815 ;
        RECT 1278.025 958.885 1278.195 959.055 ;
        RECT 1278.025 910.605 1278.195 910.775 ;
        RECT 1278.025 572.305 1278.195 572.475 ;
        RECT 1278.485 493.425 1278.655 493.595 ;
        RECT 1278.485 468.605 1278.655 468.775 ;
        RECT 1278.025 330.905 1278.195 331.075 ;
        RECT 1278.025 275.825 1278.195 275.995 ;
      LAYER met1 ;
        RECT 1278.410 1607.900 1278.730 1608.160 ;
        RECT 1278.500 1607.140 1278.640 1607.900 ;
        RECT 1278.410 1606.880 1278.730 1607.140 ;
        RECT 1277.490 1393.900 1277.810 1393.960 ;
        RECT 1279.330 1393.900 1279.650 1393.960 ;
        RECT 1277.490 1393.760 1279.650 1393.900 ;
        RECT 1277.490 1393.700 1277.810 1393.760 ;
        RECT 1279.330 1393.700 1279.650 1393.760 ;
        RECT 1277.950 1352.760 1278.270 1352.820 ;
        RECT 1279.330 1352.760 1279.650 1352.820 ;
        RECT 1277.950 1352.620 1279.650 1352.760 ;
        RECT 1277.950 1352.560 1278.270 1352.620 ;
        RECT 1279.330 1352.560 1279.650 1352.620 ;
        RECT 1277.950 1352.080 1278.270 1352.140 ;
        RECT 1277.755 1351.940 1278.270 1352.080 ;
        RECT 1277.950 1351.880 1278.270 1351.940 ;
        RECT 1277.965 1304.480 1278.255 1304.525 ;
        RECT 1278.410 1304.480 1278.730 1304.540 ;
        RECT 1277.965 1304.340 1278.730 1304.480 ;
        RECT 1277.965 1304.295 1278.255 1304.340 ;
        RECT 1278.410 1304.280 1278.730 1304.340 ;
        RECT 1277.965 1303.800 1278.255 1303.845 ;
        RECT 1278.410 1303.800 1278.730 1303.860 ;
        RECT 1277.965 1303.660 1278.730 1303.800 ;
        RECT 1277.965 1303.615 1278.255 1303.660 ;
        RECT 1278.410 1303.600 1278.730 1303.660 ;
        RECT 1277.950 1256.200 1278.270 1256.260 ;
        RECT 1277.755 1256.060 1278.270 1256.200 ;
        RECT 1277.950 1256.000 1278.270 1256.060 ;
        RECT 1278.870 1207.580 1279.190 1207.640 ;
        RECT 1279.330 1207.580 1279.650 1207.640 ;
        RECT 1278.870 1207.440 1279.650 1207.580 ;
        RECT 1278.870 1207.380 1279.190 1207.440 ;
        RECT 1279.330 1207.380 1279.650 1207.440 ;
        RECT 1278.870 1152.500 1279.190 1152.560 ;
        RECT 1279.330 1152.500 1279.650 1152.560 ;
        RECT 1278.870 1152.360 1279.650 1152.500 ;
        RECT 1278.870 1152.300 1279.190 1152.360 ;
        RECT 1279.330 1152.300 1279.650 1152.360 ;
        RECT 1277.950 1014.800 1278.270 1014.860 ;
        RECT 1278.410 1014.800 1278.730 1014.860 ;
        RECT 1277.950 1014.660 1278.730 1014.800 ;
        RECT 1277.950 1014.600 1278.270 1014.660 ;
        RECT 1278.410 1014.600 1278.730 1014.660 ;
        RECT 1277.950 959.040 1278.270 959.100 ;
        RECT 1277.755 958.900 1278.270 959.040 ;
        RECT 1277.950 958.840 1278.270 958.900 ;
        RECT 1277.950 931.500 1278.270 931.560 ;
        RECT 1277.755 931.360 1278.270 931.500 ;
        RECT 1277.950 931.300 1278.270 931.360 ;
        RECT 1277.965 910.760 1278.255 910.805 ;
        RECT 1278.410 910.760 1278.730 910.820 ;
        RECT 1277.965 910.620 1278.730 910.760 ;
        RECT 1277.965 910.575 1278.255 910.620 ;
        RECT 1278.410 910.560 1278.730 910.620 ;
        RECT 1277.950 862.820 1278.270 862.880 ;
        RECT 1277.755 862.680 1278.270 862.820 ;
        RECT 1277.950 862.620 1278.270 862.680 ;
        RECT 1277.950 821.140 1278.270 821.400 ;
        RECT 1278.040 820.660 1278.180 821.140 ;
        RECT 1278.410 820.660 1278.730 820.720 ;
        RECT 1278.040 820.520 1278.730 820.660 ;
        RECT 1278.410 820.460 1278.730 820.520 ;
        RECT 1277.950 773.400 1278.270 773.460 ;
        RECT 1278.410 773.400 1278.730 773.460 ;
        RECT 1277.950 773.260 1278.730 773.400 ;
        RECT 1277.950 773.200 1278.270 773.260 ;
        RECT 1278.410 773.200 1278.730 773.260 ;
        RECT 1276.570 765.920 1276.890 765.980 ;
        RECT 1277.950 765.920 1278.270 765.980 ;
        RECT 1276.570 765.780 1278.270 765.920 ;
        RECT 1276.570 765.720 1276.890 765.780 ;
        RECT 1277.950 765.720 1278.270 765.780 ;
        RECT 1277.490 652.360 1277.810 652.420 ;
        RECT 1278.870 652.360 1279.190 652.420 ;
        RECT 1277.490 652.220 1279.190 652.360 ;
        RECT 1277.490 652.160 1277.810 652.220 ;
        RECT 1278.870 652.160 1279.190 652.220 ;
        RECT 1277.950 572.460 1278.270 572.520 ;
        RECT 1277.755 572.320 1278.270 572.460 ;
        RECT 1277.950 572.260 1278.270 572.320 ;
        RECT 1277.950 524.520 1278.270 524.580 ;
        RECT 1277.755 524.380 1278.270 524.520 ;
        RECT 1277.950 524.320 1278.270 524.380 ;
        RECT 1277.950 493.580 1278.270 493.640 ;
        RECT 1278.425 493.580 1278.715 493.625 ;
        RECT 1277.950 493.440 1278.715 493.580 ;
        RECT 1277.950 493.380 1278.270 493.440 ;
        RECT 1278.425 493.395 1278.715 493.440 ;
        RECT 1278.410 469.440 1278.730 469.500 ;
        RECT 1278.410 469.300 1278.925 469.440 ;
        RECT 1278.410 469.240 1278.730 469.300 ;
        RECT 1278.410 468.760 1278.730 468.820 ;
        RECT 1278.215 468.620 1278.730 468.760 ;
        RECT 1278.410 468.560 1278.730 468.620 ;
        RECT 1278.425 421.160 1278.715 421.205 ;
        RECT 1278.870 421.160 1279.190 421.220 ;
        RECT 1278.425 421.020 1279.190 421.160 ;
        RECT 1278.425 420.975 1278.715 421.020 ;
        RECT 1278.870 420.960 1279.190 421.020 ;
        RECT 1277.950 387.840 1278.270 387.900 ;
        RECT 1278.870 387.840 1279.190 387.900 ;
        RECT 1277.950 387.700 1279.190 387.840 ;
        RECT 1277.950 387.640 1278.270 387.700 ;
        RECT 1278.870 387.640 1279.190 387.700 ;
        RECT 1277.950 331.060 1278.270 331.120 ;
        RECT 1277.755 330.920 1278.270 331.060 ;
        RECT 1277.950 330.860 1278.270 330.920 ;
        RECT 1277.965 323.580 1278.255 323.625 ;
        RECT 1278.870 323.580 1279.190 323.640 ;
        RECT 1277.965 323.440 1279.190 323.580 ;
        RECT 1277.965 323.395 1278.255 323.440 ;
        RECT 1278.870 323.380 1279.190 323.440 ;
        RECT 1277.965 275.980 1278.255 276.025 ;
        RECT 1278.870 275.980 1279.190 276.040 ;
        RECT 1277.965 275.840 1279.190 275.980 ;
        RECT 1277.965 275.795 1278.255 275.840 ;
        RECT 1278.870 275.780 1279.190 275.840 ;
        RECT 1277.950 228.380 1278.270 228.440 ;
        RECT 1277.755 228.240 1278.270 228.380 ;
        RECT 1277.950 228.180 1278.270 228.240 ;
        RECT 1277.950 227.700 1278.270 227.760 ;
        RECT 1278.410 227.700 1278.730 227.760 ;
        RECT 1277.950 227.560 1278.730 227.700 ;
        RECT 1277.950 227.500 1278.270 227.560 ;
        RECT 1278.410 227.500 1278.730 227.560 ;
        RECT 1276.570 113.800 1276.890 113.860 ;
        RECT 1278.410 113.800 1278.730 113.860 ;
        RECT 1276.570 113.660 1278.730 113.800 ;
        RECT 1276.570 113.600 1276.890 113.660 ;
        RECT 1278.410 113.600 1278.730 113.660 ;
        RECT 347.370 31.860 347.690 31.920 ;
        RECT 1277.030 31.860 1277.350 31.920 ;
        RECT 347.370 31.720 1277.350 31.860 ;
        RECT 347.370 31.660 347.690 31.720 ;
        RECT 1277.030 31.660 1277.350 31.720 ;
      LAYER via ;
        RECT 1278.440 1607.900 1278.700 1608.160 ;
        RECT 1278.440 1606.880 1278.700 1607.140 ;
        RECT 1277.520 1393.700 1277.780 1393.960 ;
        RECT 1279.360 1393.700 1279.620 1393.960 ;
        RECT 1277.980 1352.560 1278.240 1352.820 ;
        RECT 1279.360 1352.560 1279.620 1352.820 ;
        RECT 1277.980 1351.880 1278.240 1352.140 ;
        RECT 1278.440 1304.280 1278.700 1304.540 ;
        RECT 1278.440 1303.600 1278.700 1303.860 ;
        RECT 1277.980 1256.000 1278.240 1256.260 ;
        RECT 1278.900 1207.380 1279.160 1207.640 ;
        RECT 1279.360 1207.380 1279.620 1207.640 ;
        RECT 1278.900 1152.300 1279.160 1152.560 ;
        RECT 1279.360 1152.300 1279.620 1152.560 ;
        RECT 1277.980 1014.600 1278.240 1014.860 ;
        RECT 1278.440 1014.600 1278.700 1014.860 ;
        RECT 1277.980 958.840 1278.240 959.100 ;
        RECT 1277.980 931.300 1278.240 931.560 ;
        RECT 1278.440 910.560 1278.700 910.820 ;
        RECT 1277.980 862.620 1278.240 862.880 ;
        RECT 1277.980 821.140 1278.240 821.400 ;
        RECT 1278.440 820.460 1278.700 820.720 ;
        RECT 1277.980 773.200 1278.240 773.460 ;
        RECT 1278.440 773.200 1278.700 773.460 ;
        RECT 1276.600 765.720 1276.860 765.980 ;
        RECT 1277.980 765.720 1278.240 765.980 ;
        RECT 1277.520 652.160 1277.780 652.420 ;
        RECT 1278.900 652.160 1279.160 652.420 ;
        RECT 1277.980 572.260 1278.240 572.520 ;
        RECT 1277.980 524.320 1278.240 524.580 ;
        RECT 1277.980 493.380 1278.240 493.640 ;
        RECT 1278.440 469.240 1278.700 469.500 ;
        RECT 1278.440 468.560 1278.700 468.820 ;
        RECT 1278.900 420.960 1279.160 421.220 ;
        RECT 1277.980 387.640 1278.240 387.900 ;
        RECT 1278.900 387.640 1279.160 387.900 ;
        RECT 1277.980 330.860 1278.240 331.120 ;
        RECT 1278.900 323.380 1279.160 323.640 ;
        RECT 1278.900 275.780 1279.160 276.040 ;
        RECT 1277.980 228.180 1278.240 228.440 ;
        RECT 1277.980 227.500 1278.240 227.760 ;
        RECT 1278.440 227.500 1278.700 227.760 ;
        RECT 1276.600 113.600 1276.860 113.860 ;
        RECT 1278.440 113.600 1278.700 113.860 ;
        RECT 347.400 31.660 347.660 31.920 ;
        RECT 1277.060 31.660 1277.320 31.920 ;
      LAYER met2 ;
        RECT 1280.205 1700.410 1280.485 1704.000 ;
        RECT 1279.420 1700.270 1280.485 1700.410 ;
        RECT 1279.420 1656.210 1279.560 1700.270 ;
        RECT 1280.205 1700.000 1280.485 1700.270 ;
        RECT 1278.040 1656.070 1279.560 1656.210 ;
        RECT 1278.040 1655.530 1278.180 1656.070 ;
        RECT 1278.040 1655.390 1278.640 1655.530 ;
        RECT 1278.500 1608.190 1278.640 1655.390 ;
        RECT 1278.440 1607.870 1278.700 1608.190 ;
        RECT 1278.440 1606.850 1278.700 1607.170 ;
        RECT 1278.500 1463.090 1278.640 1606.850 ;
        RECT 1278.040 1462.950 1278.640 1463.090 ;
        RECT 1278.040 1442.010 1278.180 1462.950 ;
        RECT 1277.580 1441.870 1278.180 1442.010 ;
        RECT 1277.580 1393.990 1277.720 1441.870 ;
        RECT 1277.520 1393.670 1277.780 1393.990 ;
        RECT 1279.360 1393.670 1279.620 1393.990 ;
        RECT 1279.420 1352.850 1279.560 1393.670 ;
        RECT 1277.980 1352.530 1278.240 1352.850 ;
        RECT 1279.360 1352.530 1279.620 1352.850 ;
        RECT 1278.040 1352.170 1278.180 1352.530 ;
        RECT 1277.980 1351.850 1278.240 1352.170 ;
        RECT 1278.440 1304.250 1278.700 1304.570 ;
        RECT 1278.500 1303.890 1278.640 1304.250 ;
        RECT 1278.440 1303.570 1278.700 1303.890 ;
        RECT 1277.980 1255.970 1278.240 1256.290 ;
        RECT 1278.040 1255.805 1278.180 1255.970 ;
        RECT 1277.970 1255.435 1278.250 1255.805 ;
        RECT 1278.890 1255.435 1279.170 1255.805 ;
        RECT 1278.960 1207.670 1279.100 1255.435 ;
        RECT 1278.900 1207.350 1279.160 1207.670 ;
        RECT 1279.360 1207.350 1279.620 1207.670 ;
        RECT 1279.420 1152.590 1279.560 1207.350 ;
        RECT 1278.900 1152.270 1279.160 1152.590 ;
        RECT 1279.360 1152.270 1279.620 1152.590 ;
        RECT 1278.960 1104.050 1279.100 1152.270 ;
        RECT 1278.040 1103.910 1279.100 1104.050 ;
        RECT 1278.040 1014.890 1278.180 1103.910 ;
        RECT 1277.980 1014.570 1278.240 1014.890 ;
        RECT 1278.440 1014.570 1278.700 1014.890 ;
        RECT 1278.500 960.005 1278.640 1014.570 ;
        RECT 1278.430 959.635 1278.710 960.005 ;
        RECT 1277.970 958.955 1278.250 959.325 ;
        RECT 1277.980 958.810 1278.240 958.955 ;
        RECT 1277.980 931.270 1278.240 931.590 ;
        RECT 1278.040 910.930 1278.180 931.270 ;
        RECT 1278.040 910.850 1278.640 910.930 ;
        RECT 1278.040 910.790 1278.700 910.850 ;
        RECT 1278.440 910.530 1278.700 910.790 ;
        RECT 1277.980 862.590 1278.240 862.910 ;
        RECT 1278.040 821.430 1278.180 862.590 ;
        RECT 1277.980 821.110 1278.240 821.430 ;
        RECT 1278.440 820.430 1278.700 820.750 ;
        RECT 1278.500 773.490 1278.640 820.430 ;
        RECT 1277.980 773.170 1278.240 773.490 ;
        RECT 1278.440 773.170 1278.700 773.490 ;
        RECT 1278.040 766.010 1278.180 773.170 ;
        RECT 1276.600 765.690 1276.860 766.010 ;
        RECT 1277.980 765.690 1278.240 766.010 ;
        RECT 1276.660 717.925 1276.800 765.690 ;
        RECT 1276.590 717.555 1276.870 717.925 ;
        RECT 1277.510 717.555 1277.790 717.925 ;
        RECT 1277.580 652.450 1277.720 717.555 ;
        RECT 1277.520 652.130 1277.780 652.450 ;
        RECT 1278.900 652.130 1279.160 652.450 ;
        RECT 1278.960 580.450 1279.100 652.130 ;
        RECT 1278.500 580.310 1279.100 580.450 ;
        RECT 1278.500 579.770 1278.640 580.310 ;
        RECT 1278.040 579.630 1278.640 579.770 ;
        RECT 1278.040 572.550 1278.180 579.630 ;
        RECT 1277.980 572.230 1278.240 572.550 ;
        RECT 1277.980 524.290 1278.240 524.610 ;
        RECT 1278.040 493.670 1278.180 524.290 ;
        RECT 1277.980 493.350 1278.240 493.670 ;
        RECT 1278.440 469.210 1278.700 469.530 ;
        RECT 1278.500 468.850 1278.640 469.210 ;
        RECT 1278.440 468.530 1278.700 468.850 ;
        RECT 1278.900 420.930 1279.160 421.250 ;
        RECT 1278.960 387.930 1279.100 420.930 ;
        RECT 1277.980 387.610 1278.240 387.930 ;
        RECT 1278.900 387.610 1279.160 387.930 ;
        RECT 1278.040 331.150 1278.180 387.610 ;
        RECT 1277.980 330.830 1278.240 331.150 ;
        RECT 1278.900 323.350 1279.160 323.670 ;
        RECT 1278.960 276.070 1279.100 323.350 ;
        RECT 1278.900 275.750 1279.160 276.070 ;
        RECT 1277.980 228.150 1278.240 228.470 ;
        RECT 1278.040 227.790 1278.180 228.150 ;
        RECT 1277.980 227.470 1278.240 227.790 ;
        RECT 1278.440 227.470 1278.700 227.790 ;
        RECT 1278.500 113.890 1278.640 227.470 ;
        RECT 1276.600 113.570 1276.860 113.890 ;
        RECT 1278.440 113.570 1278.700 113.890 ;
        RECT 1276.660 61.610 1276.800 113.570 ;
        RECT 1276.660 61.470 1277.260 61.610 ;
        RECT 1277.120 31.950 1277.260 61.470 ;
        RECT 347.400 31.630 347.660 31.950 ;
        RECT 1277.060 31.630 1277.320 31.950 ;
        RECT 347.460 2.400 347.600 31.630 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 1277.970 1255.480 1278.250 1255.760 ;
        RECT 1278.890 1255.480 1279.170 1255.760 ;
        RECT 1278.430 959.680 1278.710 959.960 ;
        RECT 1277.970 959.000 1278.250 959.280 ;
        RECT 1276.590 717.600 1276.870 717.880 ;
        RECT 1277.510 717.600 1277.790 717.880 ;
      LAYER met3 ;
        RECT 1277.945 1255.770 1278.275 1255.785 ;
        RECT 1278.865 1255.770 1279.195 1255.785 ;
        RECT 1277.945 1255.470 1279.195 1255.770 ;
        RECT 1277.945 1255.455 1278.275 1255.470 ;
        RECT 1278.865 1255.455 1279.195 1255.470 ;
        RECT 1278.405 959.970 1278.735 959.985 ;
        RECT 1277.270 959.670 1278.735 959.970 ;
        RECT 1277.270 959.290 1277.570 959.670 ;
        RECT 1278.405 959.655 1278.735 959.670 ;
        RECT 1277.945 959.290 1278.275 959.305 ;
        RECT 1277.270 958.990 1278.275 959.290 ;
        RECT 1277.945 958.975 1278.275 958.990 ;
        RECT 1276.565 717.890 1276.895 717.905 ;
        RECT 1277.485 717.890 1277.815 717.905 ;
        RECT 1276.565 717.590 1277.815 717.890 ;
        RECT 1276.565 717.575 1276.895 717.590 ;
        RECT 1277.485 717.575 1277.815 717.590 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 32.200 365.630 32.260 ;
        RECT 1284.850 32.200 1285.170 32.260 ;
        RECT 365.310 32.060 1285.170 32.200 ;
        RECT 365.310 32.000 365.630 32.060 ;
        RECT 1284.850 32.000 1285.170 32.060 ;
      LAYER via ;
        RECT 365.340 32.000 365.600 32.260 ;
        RECT 1284.880 32.000 1285.140 32.260 ;
      LAYER met2 ;
        RECT 1286.645 1700.410 1286.925 1704.000 ;
        RECT 1284.940 1700.270 1286.925 1700.410 ;
        RECT 1284.940 32.290 1285.080 1700.270 ;
        RECT 1286.645 1700.000 1286.925 1700.270 ;
        RECT 365.340 31.970 365.600 32.290 ;
        RECT 1284.880 31.970 1285.140 32.290 ;
        RECT 365.400 2.400 365.540 31.970 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 32.540 383.570 32.600 ;
        RECT 1291.750 32.540 1292.070 32.600 ;
        RECT 383.250 32.400 1292.070 32.540 ;
        RECT 383.250 32.340 383.570 32.400 ;
        RECT 1291.750 32.340 1292.070 32.400 ;
      LAYER via ;
        RECT 383.280 32.340 383.540 32.600 ;
        RECT 1291.780 32.340 1292.040 32.600 ;
      LAYER met2 ;
        RECT 1293.545 1700.410 1293.825 1704.000 ;
        RECT 1291.840 1700.270 1293.825 1700.410 ;
        RECT 1291.840 32.630 1291.980 1700.270 ;
        RECT 1293.545 1700.000 1293.825 1700.270 ;
        RECT 383.280 32.310 383.540 32.630 ;
        RECT 1291.780 32.310 1292.040 32.630 ;
        RECT 383.340 2.400 383.480 32.310 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 40.360 401.510 40.420 ;
        RECT 1298.650 40.360 1298.970 40.420 ;
        RECT 401.190 40.220 1298.970 40.360 ;
        RECT 401.190 40.160 401.510 40.220 ;
        RECT 1298.650 40.160 1298.970 40.220 ;
      LAYER via ;
        RECT 401.220 40.160 401.480 40.420 ;
        RECT 1298.680 40.160 1298.940 40.420 ;
      LAYER met2 ;
        RECT 1299.985 1700.410 1300.265 1704.000 ;
        RECT 1298.740 1700.270 1300.265 1700.410 ;
        RECT 1298.740 40.450 1298.880 1700.270 ;
        RECT 1299.985 1700.000 1300.265 1700.270 ;
        RECT 401.220 40.130 401.480 40.450 ;
        RECT 1298.680 40.130 1298.940 40.450 ;
        RECT 401.280 2.400 401.420 40.130 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1167.625 1642.285 1167.795 1672.375 ;
        RECT 1167.165 655.605 1167.335 662.575 ;
        RECT 1167.165 607.325 1167.335 627.555 ;
      LAYER mcon ;
        RECT 1167.625 1672.205 1167.795 1672.375 ;
        RECT 1167.165 662.405 1167.335 662.575 ;
        RECT 1167.165 627.385 1167.335 627.555 ;
      LAYER met1 ;
        RECT 1167.565 1672.360 1167.855 1672.405 ;
        RECT 1170.310 1672.360 1170.630 1672.420 ;
        RECT 1167.565 1672.220 1170.630 1672.360 ;
        RECT 1167.565 1672.175 1167.855 1672.220 ;
        RECT 1170.310 1672.160 1170.630 1672.220 ;
        RECT 1167.550 1642.440 1167.870 1642.500 ;
        RECT 1167.355 1642.300 1167.870 1642.440 ;
        RECT 1167.550 1642.240 1167.870 1642.300 ;
        RECT 1166.630 1511.200 1166.950 1511.260 ;
        RECT 1167.550 1511.200 1167.870 1511.260 ;
        RECT 1166.630 1511.060 1167.870 1511.200 ;
        RECT 1166.630 1511.000 1166.950 1511.060 ;
        RECT 1167.550 1511.000 1167.870 1511.060 ;
        RECT 1166.630 1414.640 1166.950 1414.700 ;
        RECT 1167.550 1414.640 1167.870 1414.700 ;
        RECT 1166.630 1414.500 1167.870 1414.640 ;
        RECT 1166.630 1414.440 1166.950 1414.500 ;
        RECT 1167.550 1414.440 1167.870 1414.500 ;
        RECT 1166.630 1318.080 1166.950 1318.140 ;
        RECT 1167.550 1318.080 1167.870 1318.140 ;
        RECT 1166.630 1317.940 1167.870 1318.080 ;
        RECT 1166.630 1317.880 1166.950 1317.940 ;
        RECT 1167.550 1317.880 1167.870 1317.940 ;
        RECT 1166.630 1221.520 1166.950 1221.580 ;
        RECT 1167.550 1221.520 1167.870 1221.580 ;
        RECT 1166.630 1221.380 1167.870 1221.520 ;
        RECT 1166.630 1221.320 1166.950 1221.380 ;
        RECT 1167.550 1221.320 1167.870 1221.380 ;
        RECT 1166.630 1124.960 1166.950 1125.020 ;
        RECT 1167.550 1124.960 1167.870 1125.020 ;
        RECT 1166.630 1124.820 1167.870 1124.960 ;
        RECT 1166.630 1124.760 1166.950 1124.820 ;
        RECT 1167.550 1124.760 1167.870 1124.820 ;
        RECT 1166.630 1028.400 1166.950 1028.460 ;
        RECT 1167.550 1028.400 1167.870 1028.460 ;
        RECT 1166.630 1028.260 1167.870 1028.400 ;
        RECT 1166.630 1028.200 1166.950 1028.260 ;
        RECT 1167.550 1028.200 1167.870 1028.260 ;
        RECT 1166.630 931.840 1166.950 931.900 ;
        RECT 1167.550 931.840 1167.870 931.900 ;
        RECT 1166.630 931.700 1167.870 931.840 ;
        RECT 1166.630 931.640 1166.950 931.700 ;
        RECT 1167.550 931.640 1167.870 931.700 ;
        RECT 1166.630 835.280 1166.950 835.340 ;
        RECT 1167.550 835.280 1167.870 835.340 ;
        RECT 1166.630 835.140 1167.870 835.280 ;
        RECT 1166.630 835.080 1166.950 835.140 ;
        RECT 1167.550 835.080 1167.870 835.140 ;
        RECT 1166.630 738.380 1166.950 738.440 ;
        RECT 1167.550 738.380 1167.870 738.440 ;
        RECT 1166.630 738.240 1167.870 738.380 ;
        RECT 1166.630 738.180 1166.950 738.240 ;
        RECT 1167.550 738.180 1167.870 738.240 ;
        RECT 1167.090 662.560 1167.410 662.620 ;
        RECT 1166.895 662.420 1167.410 662.560 ;
        RECT 1167.090 662.360 1167.410 662.420 ;
        RECT 1167.090 655.760 1167.410 655.820 ;
        RECT 1166.895 655.620 1167.410 655.760 ;
        RECT 1167.090 655.560 1167.410 655.620 ;
        RECT 1167.090 627.540 1167.410 627.600 ;
        RECT 1166.895 627.400 1167.410 627.540 ;
        RECT 1167.090 627.340 1167.410 627.400 ;
        RECT 1167.090 607.480 1167.410 607.540 ;
        RECT 1166.895 607.340 1167.410 607.480 ;
        RECT 1167.090 607.280 1167.410 607.340 ;
        RECT 1166.630 448.700 1166.950 448.760 ;
        RECT 1167.550 448.700 1167.870 448.760 ;
        RECT 1166.630 448.560 1167.870 448.700 ;
        RECT 1166.630 448.500 1166.950 448.560 ;
        RECT 1167.550 448.500 1167.870 448.560 ;
        RECT 1167.090 386.480 1167.410 386.540 ;
        RECT 1167.550 386.480 1167.870 386.540 ;
        RECT 1167.090 386.340 1167.870 386.480 ;
        RECT 1167.090 386.280 1167.410 386.340 ;
        RECT 1167.550 386.280 1167.870 386.340 ;
        RECT 1167.090 324.600 1167.410 324.660 ;
        RECT 1167.550 324.600 1167.870 324.660 ;
        RECT 1167.090 324.460 1167.870 324.600 ;
        RECT 1167.090 324.400 1167.410 324.460 ;
        RECT 1167.550 324.400 1167.870 324.460 ;
        RECT 62.170 25.400 62.490 25.460 ;
        RECT 1166.170 25.400 1166.490 25.460 ;
        RECT 62.170 25.260 1166.490 25.400 ;
        RECT 62.170 25.200 62.490 25.260 ;
        RECT 1166.170 25.200 1166.490 25.260 ;
      LAYER via ;
        RECT 1170.340 1672.160 1170.600 1672.420 ;
        RECT 1167.580 1642.240 1167.840 1642.500 ;
        RECT 1166.660 1511.000 1166.920 1511.260 ;
        RECT 1167.580 1511.000 1167.840 1511.260 ;
        RECT 1166.660 1414.440 1166.920 1414.700 ;
        RECT 1167.580 1414.440 1167.840 1414.700 ;
        RECT 1166.660 1317.880 1166.920 1318.140 ;
        RECT 1167.580 1317.880 1167.840 1318.140 ;
        RECT 1166.660 1221.320 1166.920 1221.580 ;
        RECT 1167.580 1221.320 1167.840 1221.580 ;
        RECT 1166.660 1124.760 1166.920 1125.020 ;
        RECT 1167.580 1124.760 1167.840 1125.020 ;
        RECT 1166.660 1028.200 1166.920 1028.460 ;
        RECT 1167.580 1028.200 1167.840 1028.460 ;
        RECT 1166.660 931.640 1166.920 931.900 ;
        RECT 1167.580 931.640 1167.840 931.900 ;
        RECT 1166.660 835.080 1166.920 835.340 ;
        RECT 1167.580 835.080 1167.840 835.340 ;
        RECT 1166.660 738.180 1166.920 738.440 ;
        RECT 1167.580 738.180 1167.840 738.440 ;
        RECT 1167.120 662.360 1167.380 662.620 ;
        RECT 1167.120 655.560 1167.380 655.820 ;
        RECT 1167.120 627.340 1167.380 627.600 ;
        RECT 1167.120 607.280 1167.380 607.540 ;
        RECT 1166.660 448.500 1166.920 448.760 ;
        RECT 1167.580 448.500 1167.840 448.760 ;
        RECT 1167.120 386.280 1167.380 386.540 ;
        RECT 1167.580 386.280 1167.840 386.540 ;
        RECT 1167.120 324.400 1167.380 324.660 ;
        RECT 1167.580 324.400 1167.840 324.660 ;
        RECT 62.200 25.200 62.460 25.460 ;
        RECT 1166.200 25.200 1166.460 25.460 ;
      LAYER met2 ;
        RECT 1172.105 1700.410 1172.385 1704.000 ;
        RECT 1170.400 1700.270 1172.385 1700.410 ;
        RECT 1170.400 1672.450 1170.540 1700.270 ;
        RECT 1172.105 1700.000 1172.385 1700.270 ;
        RECT 1170.340 1672.130 1170.600 1672.450 ;
        RECT 1167.580 1642.210 1167.840 1642.530 ;
        RECT 1167.640 1511.290 1167.780 1642.210 ;
        RECT 1166.660 1510.970 1166.920 1511.290 ;
        RECT 1167.580 1510.970 1167.840 1511.290 ;
        RECT 1166.720 1510.690 1166.860 1510.970 ;
        RECT 1166.720 1510.550 1167.320 1510.690 ;
        RECT 1167.180 1463.090 1167.320 1510.550 ;
        RECT 1167.180 1462.950 1167.780 1463.090 ;
        RECT 1167.640 1414.730 1167.780 1462.950 ;
        RECT 1166.660 1414.410 1166.920 1414.730 ;
        RECT 1167.580 1414.410 1167.840 1414.730 ;
        RECT 1166.720 1414.130 1166.860 1414.410 ;
        RECT 1166.720 1413.990 1167.320 1414.130 ;
        RECT 1167.180 1366.530 1167.320 1413.990 ;
        RECT 1167.180 1366.390 1167.780 1366.530 ;
        RECT 1167.640 1318.170 1167.780 1366.390 ;
        RECT 1166.660 1317.850 1166.920 1318.170 ;
        RECT 1167.580 1317.850 1167.840 1318.170 ;
        RECT 1166.720 1317.570 1166.860 1317.850 ;
        RECT 1166.720 1317.430 1167.320 1317.570 ;
        RECT 1167.180 1269.970 1167.320 1317.430 ;
        RECT 1167.180 1269.830 1167.780 1269.970 ;
        RECT 1167.640 1221.610 1167.780 1269.830 ;
        RECT 1166.660 1221.290 1166.920 1221.610 ;
        RECT 1167.580 1221.290 1167.840 1221.610 ;
        RECT 1166.720 1221.010 1166.860 1221.290 ;
        RECT 1166.720 1220.870 1167.320 1221.010 ;
        RECT 1167.180 1173.410 1167.320 1220.870 ;
        RECT 1167.180 1173.270 1167.780 1173.410 ;
        RECT 1167.640 1125.050 1167.780 1173.270 ;
        RECT 1166.660 1124.730 1166.920 1125.050 ;
        RECT 1167.580 1124.730 1167.840 1125.050 ;
        RECT 1166.720 1124.450 1166.860 1124.730 ;
        RECT 1166.720 1124.310 1167.320 1124.450 ;
        RECT 1167.180 1076.850 1167.320 1124.310 ;
        RECT 1167.180 1076.710 1167.780 1076.850 ;
        RECT 1167.640 1028.490 1167.780 1076.710 ;
        RECT 1166.660 1028.170 1166.920 1028.490 ;
        RECT 1167.580 1028.170 1167.840 1028.490 ;
        RECT 1166.720 1027.890 1166.860 1028.170 ;
        RECT 1166.720 1027.750 1167.320 1027.890 ;
        RECT 1167.180 980.290 1167.320 1027.750 ;
        RECT 1167.180 980.150 1167.780 980.290 ;
        RECT 1167.640 931.930 1167.780 980.150 ;
        RECT 1166.660 931.610 1166.920 931.930 ;
        RECT 1167.580 931.610 1167.840 931.930 ;
        RECT 1166.720 931.330 1166.860 931.610 ;
        RECT 1166.720 931.190 1167.320 931.330 ;
        RECT 1167.180 917.730 1167.320 931.190 ;
        RECT 1167.180 917.590 1167.780 917.730 ;
        RECT 1167.640 835.370 1167.780 917.590 ;
        RECT 1166.660 835.050 1166.920 835.370 ;
        RECT 1167.580 835.050 1167.840 835.370 ;
        RECT 1166.720 834.770 1166.860 835.050 ;
        RECT 1166.720 834.630 1167.320 834.770 ;
        RECT 1167.180 796.690 1167.320 834.630 ;
        RECT 1167.180 796.550 1167.780 796.690 ;
        RECT 1167.640 738.470 1167.780 796.550 ;
        RECT 1166.660 738.210 1166.920 738.470 ;
        RECT 1166.660 738.150 1167.320 738.210 ;
        RECT 1167.580 738.150 1167.840 738.470 ;
        RECT 1166.720 738.070 1167.320 738.150 ;
        RECT 1167.180 662.650 1167.320 738.070 ;
        RECT 1167.120 662.330 1167.380 662.650 ;
        RECT 1167.120 655.530 1167.380 655.850 ;
        RECT 1167.180 627.630 1167.320 655.530 ;
        RECT 1167.120 627.310 1167.380 627.630 ;
        RECT 1167.120 607.250 1167.380 607.570 ;
        RECT 1167.180 594.050 1167.320 607.250 ;
        RECT 1167.180 593.910 1167.780 594.050 ;
        RECT 1167.640 524.690 1167.780 593.910 ;
        RECT 1167.180 524.550 1167.780 524.690 ;
        RECT 1167.180 500.210 1167.320 524.550 ;
        RECT 1167.180 500.070 1167.780 500.210 ;
        RECT 1167.640 448.790 1167.780 500.070 ;
        RECT 1166.660 448.530 1166.920 448.790 ;
        RECT 1166.660 448.470 1167.320 448.530 ;
        RECT 1167.580 448.470 1167.840 448.790 ;
        RECT 1166.720 448.390 1167.320 448.470 ;
        RECT 1167.180 386.570 1167.320 448.390 ;
        RECT 1167.120 386.250 1167.380 386.570 ;
        RECT 1167.580 386.250 1167.840 386.570 ;
        RECT 1167.640 324.690 1167.780 386.250 ;
        RECT 1167.120 324.370 1167.380 324.690 ;
        RECT 1167.580 324.370 1167.840 324.690 ;
        RECT 1167.180 303.690 1167.320 324.370 ;
        RECT 1167.180 303.550 1167.780 303.690 ;
        RECT 1167.640 255.410 1167.780 303.550 ;
        RECT 1166.720 255.270 1167.780 255.410 ;
        RECT 1166.720 254.730 1166.860 255.270 ;
        RECT 1166.720 254.590 1167.320 254.730 ;
        RECT 1167.180 158.850 1167.320 254.590 ;
        RECT 1166.720 158.710 1167.320 158.850 ;
        RECT 1166.720 62.290 1166.860 158.710 ;
        RECT 1166.260 62.150 1166.860 62.290 ;
        RECT 1166.260 25.490 1166.400 62.150 ;
        RECT 62.200 25.170 62.460 25.490 ;
        RECT 1166.200 25.170 1166.460 25.490 ;
        RECT 62.260 2.400 62.400 25.170 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 40.700 419.450 40.760 ;
        RECT 1305.090 40.700 1305.410 40.760 ;
        RECT 419.130 40.560 1305.410 40.700 ;
        RECT 419.130 40.500 419.450 40.560 ;
        RECT 1305.090 40.500 1305.410 40.560 ;
      LAYER via ;
        RECT 419.160 40.500 419.420 40.760 ;
        RECT 1305.120 40.500 1305.380 40.760 ;
      LAYER met2 ;
        RECT 1306.885 1700.410 1307.165 1704.000 ;
        RECT 1305.180 1700.270 1307.165 1700.410 ;
        RECT 1305.180 40.790 1305.320 1700.270 ;
        RECT 1306.885 1700.000 1307.165 1700.270 ;
        RECT 419.160 40.470 419.420 40.790 ;
        RECT 1305.120 40.470 1305.380 40.790 ;
        RECT 419.220 2.400 419.360 40.470 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.990 1394.580 1312.310 1394.640 ;
        RECT 1311.620 1394.440 1312.310 1394.580 ;
        RECT 1311.620 1393.900 1311.760 1394.440 ;
        RECT 1311.990 1394.380 1312.310 1394.440 ;
        RECT 1311.990 1393.900 1312.310 1393.960 ;
        RECT 1311.620 1393.760 1312.310 1393.900 ;
        RECT 1311.990 1393.700 1312.310 1393.760 ;
        RECT 436.610 41.040 436.930 41.100 ;
        RECT 1311.990 41.040 1312.310 41.100 ;
        RECT 436.610 40.900 1312.310 41.040 ;
        RECT 436.610 40.840 436.930 40.900 ;
        RECT 1311.990 40.840 1312.310 40.900 ;
      LAYER via ;
        RECT 1312.020 1394.380 1312.280 1394.640 ;
        RECT 1312.020 1393.700 1312.280 1393.960 ;
        RECT 436.640 40.840 436.900 41.100 ;
        RECT 1312.020 40.840 1312.280 41.100 ;
      LAYER met2 ;
        RECT 1313.785 1700.410 1314.065 1704.000 ;
        RECT 1312.080 1700.270 1314.065 1700.410 ;
        RECT 1312.080 1394.670 1312.220 1700.270 ;
        RECT 1313.785 1700.000 1314.065 1700.270 ;
        RECT 1312.020 1394.350 1312.280 1394.670 ;
        RECT 1312.020 1393.670 1312.280 1393.990 ;
        RECT 1312.080 41.130 1312.220 1393.670 ;
        RECT 436.640 40.810 436.900 41.130 ;
        RECT 1312.020 40.810 1312.280 41.130 ;
        RECT 436.700 2.400 436.840 40.810 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.010 53.280 455.330 53.340 ;
        RECT 1318.890 53.280 1319.210 53.340 ;
        RECT 455.010 53.140 1319.210 53.280 ;
        RECT 455.010 53.080 455.330 53.140 ;
        RECT 1318.890 53.080 1319.210 53.140 ;
      LAYER via ;
        RECT 455.040 53.080 455.300 53.340 ;
        RECT 1318.920 53.080 1319.180 53.340 ;
      LAYER met2 ;
        RECT 1320.225 1700.410 1320.505 1704.000 ;
        RECT 1318.980 1700.270 1320.505 1700.410 ;
        RECT 1318.980 53.370 1319.120 1700.270 ;
        RECT 1320.225 1700.000 1320.505 1700.270 ;
        RECT 455.040 53.050 455.300 53.370 ;
        RECT 1318.920 53.050 1319.180 53.370 ;
        RECT 455.100 17.410 455.240 53.050 ;
        RECT 454.640 17.270 455.240 17.410 ;
        RECT 454.640 2.400 454.780 17.270 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.710 53.620 476.030 53.680 ;
        RECT 1325.790 53.620 1326.110 53.680 ;
        RECT 475.710 53.480 1326.110 53.620 ;
        RECT 475.710 53.420 476.030 53.480 ;
        RECT 1325.790 53.420 1326.110 53.480 ;
        RECT 472.490 15.540 472.810 15.600 ;
        RECT 475.710 15.540 476.030 15.600 ;
        RECT 472.490 15.400 476.030 15.540 ;
        RECT 472.490 15.340 472.810 15.400 ;
        RECT 475.710 15.340 476.030 15.400 ;
      LAYER via ;
        RECT 475.740 53.420 476.000 53.680 ;
        RECT 1325.820 53.420 1326.080 53.680 ;
        RECT 472.520 15.340 472.780 15.600 ;
        RECT 475.740 15.340 476.000 15.600 ;
      LAYER met2 ;
        RECT 1327.125 1700.410 1327.405 1704.000 ;
        RECT 1325.880 1700.270 1327.405 1700.410 ;
        RECT 1325.880 53.710 1326.020 1700.270 ;
        RECT 1327.125 1700.000 1327.405 1700.270 ;
        RECT 475.740 53.390 476.000 53.710 ;
        RECT 1325.820 53.390 1326.080 53.710 ;
        RECT 475.800 15.630 475.940 53.390 ;
        RECT 472.520 15.310 472.780 15.630 ;
        RECT 475.740 15.310 476.000 15.630 ;
        RECT 472.580 2.400 472.720 15.310 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 53.960 496.270 54.020 ;
        RECT 1332.690 53.960 1333.010 54.020 ;
        RECT 495.950 53.820 1333.010 53.960 ;
        RECT 495.950 53.760 496.270 53.820 ;
        RECT 1332.690 53.760 1333.010 53.820 ;
        RECT 490.430 15.540 490.750 15.600 ;
        RECT 495.950 15.540 496.270 15.600 ;
        RECT 490.430 15.400 496.270 15.540 ;
        RECT 490.430 15.340 490.750 15.400 ;
        RECT 495.950 15.340 496.270 15.400 ;
      LAYER via ;
        RECT 495.980 53.760 496.240 54.020 ;
        RECT 1332.720 53.760 1332.980 54.020 ;
        RECT 490.460 15.340 490.720 15.600 ;
        RECT 495.980 15.340 496.240 15.600 ;
      LAYER met2 ;
        RECT 1334.025 1700.410 1334.305 1704.000 ;
        RECT 1332.780 1700.270 1334.305 1700.410 ;
        RECT 1332.780 54.050 1332.920 1700.270 ;
        RECT 1334.025 1700.000 1334.305 1700.270 ;
        RECT 495.980 53.730 496.240 54.050 ;
        RECT 1332.720 53.730 1332.980 54.050 ;
        RECT 496.040 15.630 496.180 53.730 ;
        RECT 490.460 15.310 490.720 15.630 ;
        RECT 495.980 15.310 496.240 15.630 ;
        RECT 490.520 2.400 490.660 15.310 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 54.300 510.530 54.360 ;
        RECT 1339.590 54.300 1339.910 54.360 ;
        RECT 510.210 54.160 1339.910 54.300 ;
        RECT 510.210 54.100 510.530 54.160 ;
        RECT 1339.590 54.100 1339.910 54.160 ;
        RECT 507.910 15.540 508.230 15.600 ;
        RECT 510.210 15.540 510.530 15.600 ;
        RECT 507.910 15.400 510.530 15.540 ;
        RECT 507.910 15.340 508.230 15.400 ;
        RECT 510.210 15.340 510.530 15.400 ;
      LAYER via ;
        RECT 510.240 54.100 510.500 54.360 ;
        RECT 1339.620 54.100 1339.880 54.360 ;
        RECT 507.940 15.340 508.200 15.600 ;
        RECT 510.240 15.340 510.500 15.600 ;
      LAYER met2 ;
        RECT 1340.465 1700.410 1340.745 1704.000 ;
        RECT 1339.680 1700.270 1340.745 1700.410 ;
        RECT 1339.680 54.390 1339.820 1700.270 ;
        RECT 1340.465 1700.000 1340.745 1700.270 ;
        RECT 510.240 54.070 510.500 54.390 ;
        RECT 1339.620 54.070 1339.880 54.390 ;
        RECT 510.300 15.630 510.440 54.070 ;
        RECT 507.940 15.310 508.200 15.630 ;
        RECT 510.240 15.310 510.500 15.630 ;
        RECT 508.000 2.400 508.140 15.310 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.910 54.640 531.230 54.700 ;
        RECT 1346.490 54.640 1346.810 54.700 ;
        RECT 530.910 54.500 1346.810 54.640 ;
        RECT 530.910 54.440 531.230 54.500 ;
        RECT 1346.490 54.440 1346.810 54.500 ;
        RECT 525.850 15.540 526.170 15.600 ;
        RECT 530.910 15.540 531.230 15.600 ;
        RECT 525.850 15.400 531.230 15.540 ;
        RECT 525.850 15.340 526.170 15.400 ;
        RECT 530.910 15.340 531.230 15.400 ;
      LAYER via ;
        RECT 530.940 54.440 531.200 54.700 ;
        RECT 1346.520 54.440 1346.780 54.700 ;
        RECT 525.880 15.340 526.140 15.600 ;
        RECT 530.940 15.340 531.200 15.600 ;
      LAYER met2 ;
        RECT 1347.365 1700.410 1347.645 1704.000 ;
        RECT 1346.580 1700.270 1347.645 1700.410 ;
        RECT 1346.580 54.730 1346.720 1700.270 ;
        RECT 1347.365 1700.000 1347.645 1700.270 ;
        RECT 530.940 54.410 531.200 54.730 ;
        RECT 1346.520 54.410 1346.780 54.730 ;
        RECT 531.000 15.630 531.140 54.410 ;
        RECT 525.880 15.310 526.140 15.630 ;
        RECT 530.940 15.310 531.200 15.630 ;
        RECT 525.940 2.400 526.080 15.310 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 544.710 54.980 545.030 55.040 ;
        RECT 1353.390 54.980 1353.710 55.040 ;
        RECT 544.710 54.840 1353.710 54.980 ;
        RECT 544.710 54.780 545.030 54.840 ;
        RECT 1353.390 54.780 1353.710 54.840 ;
      LAYER via ;
        RECT 544.740 54.780 545.000 55.040 ;
        RECT 1353.420 54.780 1353.680 55.040 ;
      LAYER met2 ;
        RECT 1354.265 1700.410 1354.545 1704.000 ;
        RECT 1353.480 1700.270 1354.545 1700.410 ;
        RECT 1353.480 55.070 1353.620 1700.270 ;
        RECT 1354.265 1700.000 1354.545 1700.270 ;
        RECT 544.740 54.750 545.000 55.070 ;
        RECT 1353.420 54.750 1353.680 55.070 ;
        RECT 544.800 16.730 544.940 54.750 ;
        RECT 543.880 16.590 544.940 16.730 ;
        RECT 543.880 2.400 544.020 16.590 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 51.240 565.730 51.300 ;
        RECT 1360.290 51.240 1360.610 51.300 ;
        RECT 565.410 51.100 1360.610 51.240 ;
        RECT 565.410 51.040 565.730 51.100 ;
        RECT 1360.290 51.040 1360.610 51.100 ;
        RECT 561.730 14.860 562.050 14.920 ;
        RECT 565.410 14.860 565.730 14.920 ;
        RECT 561.730 14.720 565.730 14.860 ;
        RECT 561.730 14.660 562.050 14.720 ;
        RECT 565.410 14.660 565.730 14.720 ;
      LAYER via ;
        RECT 565.440 51.040 565.700 51.300 ;
        RECT 1360.320 51.040 1360.580 51.300 ;
        RECT 561.760 14.660 562.020 14.920 ;
        RECT 565.440 14.660 565.700 14.920 ;
      LAYER met2 ;
        RECT 1360.705 1700.410 1360.985 1704.000 ;
        RECT 1360.380 1700.270 1360.985 1700.410 ;
        RECT 1360.380 51.330 1360.520 1700.270 ;
        RECT 1360.705 1700.000 1360.985 1700.270 ;
        RECT 565.440 51.010 565.700 51.330 ;
        RECT 1360.320 51.010 1360.580 51.330 ;
        RECT 565.500 14.950 565.640 51.010 ;
        RECT 561.760 14.630 562.020 14.950 ;
        RECT 565.440 14.630 565.700 14.950 ;
        RECT 561.820 2.400 561.960 14.630 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1367.650 1677.120 1367.970 1677.180 ;
        RECT 1367.280 1676.980 1367.970 1677.120 ;
        RECT 1367.280 1676.160 1367.420 1676.980 ;
        RECT 1367.650 1676.920 1367.970 1676.980 ;
        RECT 1367.190 1675.900 1367.510 1676.160 ;
        RECT 585.650 50.900 585.970 50.960 ;
        RECT 1367.190 50.900 1367.510 50.960 ;
        RECT 585.650 50.760 1367.510 50.900 ;
        RECT 585.650 50.700 585.970 50.760 ;
        RECT 1367.190 50.700 1367.510 50.760 ;
        RECT 579.670 14.860 579.990 14.920 ;
        RECT 584.730 14.860 585.050 14.920 ;
        RECT 579.670 14.720 585.050 14.860 ;
        RECT 579.670 14.660 579.990 14.720 ;
        RECT 584.730 14.660 585.050 14.720 ;
      LAYER via ;
        RECT 1367.680 1676.920 1367.940 1677.180 ;
        RECT 1367.220 1675.900 1367.480 1676.160 ;
        RECT 585.680 50.700 585.940 50.960 ;
        RECT 1367.220 50.700 1367.480 50.960 ;
        RECT 579.700 14.660 579.960 14.920 ;
        RECT 584.760 14.660 585.020 14.920 ;
      LAYER met2 ;
        RECT 1367.605 1700.000 1367.885 1704.000 ;
        RECT 1367.740 1677.210 1367.880 1700.000 ;
        RECT 1367.680 1676.890 1367.940 1677.210 ;
        RECT 1367.220 1675.870 1367.480 1676.190 ;
        RECT 1367.280 50.990 1367.420 1675.870 ;
        RECT 585.680 50.670 585.940 50.990 ;
        RECT 1367.220 50.670 1367.480 50.990 ;
        RECT 585.740 18.090 585.880 50.670 ;
        RECT 584.820 17.950 585.880 18.090 ;
        RECT 584.820 14.950 584.960 17.950 ;
        RECT 579.700 14.630 579.960 14.950 ;
        RECT 584.760 14.630 585.020 14.950 ;
        RECT 579.760 2.400 579.900 14.630 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 38.320 86.410 38.380 ;
        RECT 1180.890 38.320 1181.210 38.380 ;
        RECT 86.090 38.180 1181.210 38.320 ;
        RECT 86.090 38.120 86.410 38.180 ;
        RECT 1180.890 38.120 1181.210 38.180 ;
      LAYER via ;
        RECT 86.120 38.120 86.380 38.380 ;
        RECT 1180.920 38.120 1181.180 38.380 ;
      LAYER met2 ;
        RECT 1181.305 1700.410 1181.585 1704.000 ;
        RECT 1180.980 1700.270 1181.585 1700.410 ;
        RECT 1180.980 38.410 1181.120 1700.270 ;
        RECT 1181.305 1700.000 1181.585 1700.270 ;
        RECT 86.120 38.090 86.380 38.410 ;
        RECT 1180.920 38.090 1181.180 38.410 ;
        RECT 86.180 2.400 86.320 38.090 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 50.560 600.230 50.620 ;
        RECT 1374.090 50.560 1374.410 50.620 ;
        RECT 599.910 50.420 1374.410 50.560 ;
        RECT 599.910 50.360 600.230 50.420 ;
        RECT 1374.090 50.360 1374.410 50.420 ;
        RECT 597.150 14.860 597.470 14.920 ;
        RECT 599.910 14.860 600.230 14.920 ;
        RECT 597.150 14.720 600.230 14.860 ;
        RECT 597.150 14.660 597.470 14.720 ;
        RECT 599.910 14.660 600.230 14.720 ;
      LAYER via ;
        RECT 599.940 50.360 600.200 50.620 ;
        RECT 1374.120 50.360 1374.380 50.620 ;
        RECT 597.180 14.660 597.440 14.920 ;
        RECT 599.940 14.660 600.200 14.920 ;
      LAYER met2 ;
        RECT 1374.045 1700.000 1374.325 1704.000 ;
        RECT 1374.180 50.650 1374.320 1700.000 ;
        RECT 599.940 50.330 600.200 50.650 ;
        RECT 1374.120 50.330 1374.380 50.650 ;
        RECT 600.000 14.950 600.140 50.330 ;
        RECT 597.180 14.630 597.440 14.950 ;
        RECT 599.940 14.630 600.200 14.950 ;
        RECT 597.240 2.400 597.380 14.630 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 50.220 620.930 50.280 ;
        RECT 1380.990 50.220 1381.310 50.280 ;
        RECT 620.610 50.080 1381.310 50.220 ;
        RECT 620.610 50.020 620.930 50.080 ;
        RECT 1380.990 50.020 1381.310 50.080 ;
      LAYER via ;
        RECT 620.640 50.020 620.900 50.280 ;
        RECT 1381.020 50.020 1381.280 50.280 ;
      LAYER met2 ;
        RECT 1380.945 1700.000 1381.225 1704.000 ;
        RECT 1381.080 50.310 1381.220 1700.000 ;
        RECT 620.640 49.990 620.900 50.310 ;
        RECT 1381.020 49.990 1381.280 50.310 ;
        RECT 620.700 17.410 620.840 49.990 ;
        RECT 615.180 17.270 620.840 17.410 ;
        RECT 615.180 2.400 615.320 17.270 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 38.660 109.870 38.720 ;
        RECT 1188.250 38.660 1188.570 38.720 ;
        RECT 109.550 38.520 1188.570 38.660 ;
        RECT 109.550 38.460 109.870 38.520 ;
        RECT 1188.250 38.460 1188.570 38.520 ;
      LAYER via ;
        RECT 109.580 38.460 109.840 38.720 ;
        RECT 1188.280 38.460 1188.540 38.720 ;
      LAYER met2 ;
        RECT 1190.045 1700.410 1190.325 1704.000 ;
        RECT 1188.340 1700.270 1190.325 1700.410 ;
        RECT 1188.340 38.750 1188.480 1700.270 ;
        RECT 1190.045 1700.000 1190.325 1700.270 ;
        RECT 109.580 38.430 109.840 38.750 ;
        RECT 1188.280 38.430 1188.540 38.750 ;
        RECT 109.640 2.400 109.780 38.430 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1195.685 1594.005 1195.855 1683.595 ;
        RECT 1196.605 1338.665 1196.775 1370.455 ;
        RECT 1195.685 1200.625 1195.855 1249.415 ;
        RECT 1195.685 1013.965 1195.855 1055.615 ;
        RECT 1195.685 869.125 1195.855 910.775 ;
        RECT 1195.225 758.965 1195.395 773.415 ;
        RECT 1195.685 662.405 1195.855 710.515 ;
        RECT 1195.225 255.085 1195.395 289.595 ;
        RECT 1194.765 41.565 1194.935 131.155 ;
      LAYER mcon ;
        RECT 1195.685 1683.425 1195.855 1683.595 ;
        RECT 1196.605 1370.285 1196.775 1370.455 ;
        RECT 1195.685 1249.245 1195.855 1249.415 ;
        RECT 1195.685 1055.445 1195.855 1055.615 ;
        RECT 1195.685 910.605 1195.855 910.775 ;
        RECT 1195.225 773.245 1195.395 773.415 ;
        RECT 1195.685 710.345 1195.855 710.515 ;
        RECT 1195.225 289.425 1195.395 289.595 ;
        RECT 1194.765 130.985 1194.935 131.155 ;
      LAYER met1 ;
        RECT 1195.610 1690.720 1195.930 1690.780 ;
        RECT 1199.290 1690.720 1199.610 1690.780 ;
        RECT 1195.610 1690.580 1199.610 1690.720 ;
        RECT 1195.610 1690.520 1195.930 1690.580 ;
        RECT 1199.290 1690.520 1199.610 1690.580 ;
        RECT 1195.610 1683.580 1195.930 1683.640 ;
        RECT 1195.415 1683.440 1195.930 1683.580 ;
        RECT 1195.610 1683.380 1195.930 1683.440 ;
        RECT 1195.610 1594.160 1195.930 1594.220 ;
        RECT 1195.415 1594.020 1195.930 1594.160 ;
        RECT 1195.610 1593.960 1195.930 1594.020 ;
        RECT 1195.150 1490.460 1195.470 1490.520 ;
        RECT 1195.610 1490.460 1195.930 1490.520 ;
        RECT 1195.150 1490.320 1195.930 1490.460 ;
        RECT 1195.150 1490.260 1195.470 1490.320 ;
        RECT 1195.610 1490.260 1195.930 1490.320 ;
        RECT 1195.610 1393.900 1195.930 1393.960 ;
        RECT 1196.530 1393.900 1196.850 1393.960 ;
        RECT 1195.610 1393.760 1196.850 1393.900 ;
        RECT 1195.610 1393.700 1195.930 1393.760 ;
        RECT 1196.530 1393.700 1196.850 1393.760 ;
        RECT 1195.610 1370.440 1195.930 1370.500 ;
        RECT 1196.545 1370.440 1196.835 1370.485 ;
        RECT 1195.610 1370.300 1196.835 1370.440 ;
        RECT 1195.610 1370.240 1195.930 1370.300 ;
        RECT 1196.545 1370.255 1196.835 1370.300 ;
        RECT 1196.530 1338.820 1196.850 1338.880 ;
        RECT 1196.530 1338.680 1197.045 1338.820 ;
        RECT 1196.530 1338.620 1196.850 1338.680 ;
        RECT 1195.610 1297.340 1195.930 1297.400 ;
        RECT 1196.530 1297.340 1196.850 1297.400 ;
        RECT 1195.610 1297.200 1196.850 1297.340 ;
        RECT 1195.610 1297.140 1195.930 1297.200 ;
        RECT 1196.530 1297.140 1196.850 1297.200 ;
        RECT 1195.625 1249.400 1195.915 1249.445 ;
        RECT 1196.070 1249.400 1196.390 1249.460 ;
        RECT 1195.625 1249.260 1196.390 1249.400 ;
        RECT 1195.625 1249.215 1195.915 1249.260 ;
        RECT 1196.070 1249.200 1196.390 1249.260 ;
        RECT 1195.610 1200.780 1195.930 1200.840 ;
        RECT 1195.415 1200.640 1195.930 1200.780 ;
        RECT 1195.610 1200.580 1195.930 1200.640 ;
        RECT 1195.610 1104.220 1195.930 1104.280 ;
        RECT 1196.070 1104.220 1196.390 1104.280 ;
        RECT 1195.610 1104.080 1196.390 1104.220 ;
        RECT 1195.610 1104.020 1195.930 1104.080 ;
        RECT 1196.070 1104.020 1196.390 1104.080 ;
        RECT 1195.150 1056.280 1195.470 1056.340 ;
        RECT 1195.610 1056.280 1195.930 1056.340 ;
        RECT 1195.150 1056.140 1195.930 1056.280 ;
        RECT 1195.150 1056.080 1195.470 1056.140 ;
        RECT 1195.610 1056.080 1195.930 1056.140 ;
        RECT 1195.610 1055.600 1195.930 1055.660 ;
        RECT 1195.415 1055.460 1195.930 1055.600 ;
        RECT 1195.610 1055.400 1195.930 1055.460 ;
        RECT 1195.610 1014.120 1195.930 1014.180 ;
        RECT 1195.415 1013.980 1195.930 1014.120 ;
        RECT 1195.610 1013.920 1195.930 1013.980 ;
        RECT 1195.610 965.980 1195.930 966.240 ;
        RECT 1195.700 965.840 1195.840 965.980 ;
        RECT 1196.070 965.840 1196.390 965.900 ;
        RECT 1195.700 965.700 1196.390 965.840 ;
        RECT 1196.070 965.640 1196.390 965.700 ;
        RECT 1195.610 917.900 1195.930 917.960 ;
        RECT 1196.070 917.900 1196.390 917.960 ;
        RECT 1195.610 917.760 1196.390 917.900 ;
        RECT 1195.610 917.700 1195.930 917.760 ;
        RECT 1196.070 917.700 1196.390 917.760 ;
        RECT 1195.610 910.760 1195.930 910.820 ;
        RECT 1195.415 910.620 1195.930 910.760 ;
        RECT 1195.610 910.560 1195.930 910.620 ;
        RECT 1195.610 869.280 1195.930 869.340 ;
        RECT 1195.415 869.140 1195.930 869.280 ;
        RECT 1195.610 869.080 1195.930 869.140 ;
        RECT 1195.610 845.480 1195.930 845.540 ;
        RECT 1196.530 845.480 1196.850 845.540 ;
        RECT 1195.610 845.340 1196.850 845.480 ;
        RECT 1195.610 845.280 1195.930 845.340 ;
        RECT 1196.530 845.280 1196.850 845.340 ;
        RECT 1195.165 773.400 1195.455 773.445 ;
        RECT 1195.610 773.400 1195.930 773.460 ;
        RECT 1195.165 773.260 1195.930 773.400 ;
        RECT 1195.165 773.215 1195.455 773.260 ;
        RECT 1195.610 773.200 1195.930 773.260 ;
        RECT 1195.150 759.120 1195.470 759.180 ;
        RECT 1194.955 758.980 1195.470 759.120 ;
        RECT 1195.150 758.920 1195.470 758.980 ;
        RECT 1195.150 717.640 1195.470 717.700 ;
        RECT 1195.610 717.640 1195.930 717.700 ;
        RECT 1195.150 717.500 1195.930 717.640 ;
        RECT 1195.150 717.440 1195.470 717.500 ;
        RECT 1195.610 717.440 1195.930 717.500 ;
        RECT 1195.610 710.500 1195.930 710.560 ;
        RECT 1195.415 710.360 1195.930 710.500 ;
        RECT 1195.610 710.300 1195.930 710.360 ;
        RECT 1195.610 662.560 1195.930 662.620 ;
        RECT 1195.415 662.420 1195.930 662.560 ;
        RECT 1195.610 662.360 1195.930 662.420 ;
        RECT 1195.610 545.400 1195.930 545.660 ;
        RECT 1194.690 544.580 1195.010 544.640 ;
        RECT 1195.700 544.580 1195.840 545.400 ;
        RECT 1194.690 544.440 1195.840 544.580 ;
        RECT 1194.690 544.380 1195.010 544.440 ;
        RECT 1194.690 500.380 1195.010 500.440 ;
        RECT 1195.610 500.380 1195.930 500.440 ;
        RECT 1194.690 500.240 1195.930 500.380 ;
        RECT 1194.690 500.180 1195.010 500.240 ;
        RECT 1195.610 500.180 1195.930 500.240 ;
        RECT 1195.165 289.580 1195.455 289.625 ;
        RECT 1195.610 289.580 1195.930 289.640 ;
        RECT 1195.165 289.440 1195.930 289.580 ;
        RECT 1195.165 289.395 1195.455 289.440 ;
        RECT 1195.610 289.380 1195.930 289.440 ;
        RECT 1195.150 255.240 1195.470 255.300 ;
        RECT 1194.955 255.100 1195.470 255.240 ;
        RECT 1195.150 255.040 1195.470 255.100 ;
        RECT 1195.150 241.300 1195.470 241.360 ;
        RECT 1195.610 241.300 1195.930 241.360 ;
        RECT 1195.150 241.160 1195.930 241.300 ;
        RECT 1195.150 241.100 1195.470 241.160 ;
        RECT 1195.610 241.100 1195.930 241.160 ;
        RECT 1194.705 131.140 1194.995 131.185 ;
        RECT 1195.610 131.140 1195.930 131.200 ;
        RECT 1194.705 131.000 1195.930 131.140 ;
        RECT 1194.705 130.955 1194.995 131.000 ;
        RECT 1195.610 130.940 1195.930 131.000 ;
        RECT 1194.705 41.720 1194.995 41.765 ;
        RECT 1195.150 41.720 1195.470 41.780 ;
        RECT 1194.705 41.580 1195.470 41.720 ;
        RECT 1194.705 41.535 1194.995 41.580 ;
        RECT 1195.150 41.520 1195.470 41.580 ;
        RECT 133.470 39.000 133.790 39.060 ;
        RECT 1195.150 39.000 1195.470 39.060 ;
        RECT 133.470 38.860 1195.470 39.000 ;
        RECT 133.470 38.800 133.790 38.860 ;
        RECT 1195.150 38.800 1195.470 38.860 ;
      LAYER via ;
        RECT 1195.640 1690.520 1195.900 1690.780 ;
        RECT 1199.320 1690.520 1199.580 1690.780 ;
        RECT 1195.640 1683.380 1195.900 1683.640 ;
        RECT 1195.640 1593.960 1195.900 1594.220 ;
        RECT 1195.180 1490.260 1195.440 1490.520 ;
        RECT 1195.640 1490.260 1195.900 1490.520 ;
        RECT 1195.640 1393.700 1195.900 1393.960 ;
        RECT 1196.560 1393.700 1196.820 1393.960 ;
        RECT 1195.640 1370.240 1195.900 1370.500 ;
        RECT 1196.560 1338.620 1196.820 1338.880 ;
        RECT 1195.640 1297.140 1195.900 1297.400 ;
        RECT 1196.560 1297.140 1196.820 1297.400 ;
        RECT 1196.100 1249.200 1196.360 1249.460 ;
        RECT 1195.640 1200.580 1195.900 1200.840 ;
        RECT 1195.640 1104.020 1195.900 1104.280 ;
        RECT 1196.100 1104.020 1196.360 1104.280 ;
        RECT 1195.180 1056.080 1195.440 1056.340 ;
        RECT 1195.640 1056.080 1195.900 1056.340 ;
        RECT 1195.640 1055.400 1195.900 1055.660 ;
        RECT 1195.640 1013.920 1195.900 1014.180 ;
        RECT 1195.640 965.980 1195.900 966.240 ;
        RECT 1196.100 965.640 1196.360 965.900 ;
        RECT 1195.640 917.700 1195.900 917.960 ;
        RECT 1196.100 917.700 1196.360 917.960 ;
        RECT 1195.640 910.560 1195.900 910.820 ;
        RECT 1195.640 869.080 1195.900 869.340 ;
        RECT 1195.640 845.280 1195.900 845.540 ;
        RECT 1196.560 845.280 1196.820 845.540 ;
        RECT 1195.640 773.200 1195.900 773.460 ;
        RECT 1195.180 758.920 1195.440 759.180 ;
        RECT 1195.180 717.440 1195.440 717.700 ;
        RECT 1195.640 717.440 1195.900 717.700 ;
        RECT 1195.640 710.300 1195.900 710.560 ;
        RECT 1195.640 662.360 1195.900 662.620 ;
        RECT 1195.640 545.400 1195.900 545.660 ;
        RECT 1194.720 544.380 1194.980 544.640 ;
        RECT 1194.720 500.180 1194.980 500.440 ;
        RECT 1195.640 500.180 1195.900 500.440 ;
        RECT 1195.640 289.380 1195.900 289.640 ;
        RECT 1195.180 255.040 1195.440 255.300 ;
        RECT 1195.180 241.100 1195.440 241.360 ;
        RECT 1195.640 241.100 1195.900 241.360 ;
        RECT 1195.640 130.940 1195.900 131.200 ;
        RECT 1195.180 41.520 1195.440 41.780 ;
        RECT 133.500 38.800 133.760 39.060 ;
        RECT 1195.180 38.800 1195.440 39.060 ;
      LAYER met2 ;
        RECT 1199.245 1700.000 1199.525 1704.000 ;
        RECT 1199.380 1690.810 1199.520 1700.000 ;
        RECT 1195.640 1690.490 1195.900 1690.810 ;
        RECT 1199.320 1690.490 1199.580 1690.810 ;
        RECT 1195.700 1683.670 1195.840 1690.490 ;
        RECT 1195.640 1683.350 1195.900 1683.670 ;
        RECT 1195.640 1593.930 1195.900 1594.250 ;
        RECT 1195.700 1490.550 1195.840 1593.930 ;
        RECT 1195.180 1490.230 1195.440 1490.550 ;
        RECT 1195.640 1490.230 1195.900 1490.550 ;
        RECT 1195.240 1483.605 1195.380 1490.230 ;
        RECT 1195.170 1483.235 1195.450 1483.605 ;
        RECT 1196.550 1483.235 1196.830 1483.605 ;
        RECT 1196.620 1393.990 1196.760 1483.235 ;
        RECT 1195.640 1393.670 1195.900 1393.990 ;
        RECT 1196.560 1393.670 1196.820 1393.990 ;
        RECT 1195.700 1370.530 1195.840 1393.670 ;
        RECT 1195.640 1370.210 1195.900 1370.530 ;
        RECT 1196.560 1338.590 1196.820 1338.910 ;
        RECT 1195.700 1297.430 1195.840 1297.585 ;
        RECT 1196.620 1297.430 1196.760 1338.590 ;
        RECT 1195.640 1297.170 1195.900 1297.430 ;
        RECT 1195.640 1297.110 1196.300 1297.170 ;
        RECT 1196.560 1297.110 1196.820 1297.430 ;
        RECT 1195.700 1297.030 1196.300 1297.110 ;
        RECT 1196.160 1249.490 1196.300 1297.030 ;
        RECT 1196.100 1249.170 1196.360 1249.490 ;
        RECT 1195.640 1200.725 1195.900 1200.870 ;
        RECT 1195.630 1200.355 1195.910 1200.725 ;
        RECT 1196.090 1199.675 1196.370 1200.045 ;
        RECT 1196.160 1104.310 1196.300 1199.675 ;
        RECT 1195.640 1104.165 1195.900 1104.310 ;
        RECT 1195.630 1103.795 1195.910 1104.165 ;
        RECT 1196.100 1103.990 1196.360 1104.310 ;
        RECT 1195.170 1103.115 1195.450 1103.485 ;
        RECT 1195.240 1056.370 1195.380 1103.115 ;
        RECT 1195.180 1056.050 1195.440 1056.370 ;
        RECT 1195.640 1056.050 1195.900 1056.370 ;
        RECT 1195.700 1055.690 1195.840 1056.050 ;
        RECT 1195.640 1055.370 1195.900 1055.690 ;
        RECT 1195.640 1013.890 1195.900 1014.210 ;
        RECT 1195.700 966.270 1195.840 1013.890 ;
        RECT 1195.640 965.950 1195.900 966.270 ;
        RECT 1196.100 965.610 1196.360 965.930 ;
        RECT 1196.160 917.990 1196.300 965.610 ;
        RECT 1195.640 917.670 1195.900 917.990 ;
        RECT 1196.100 917.670 1196.360 917.990 ;
        RECT 1195.700 910.850 1195.840 917.670 ;
        RECT 1195.640 910.530 1195.900 910.850 ;
        RECT 1195.640 869.050 1195.900 869.370 ;
        RECT 1195.700 845.570 1195.840 869.050 ;
        RECT 1195.640 845.250 1195.900 845.570 ;
        RECT 1196.560 845.250 1196.820 845.570 ;
        RECT 1196.620 821.285 1196.760 845.250 ;
        RECT 1195.630 820.915 1195.910 821.285 ;
        RECT 1196.550 820.915 1196.830 821.285 ;
        RECT 1195.700 773.490 1195.840 820.915 ;
        RECT 1195.640 773.170 1195.900 773.490 ;
        RECT 1195.180 758.890 1195.440 759.210 ;
        RECT 1195.240 717.730 1195.380 758.890 ;
        RECT 1195.180 717.410 1195.440 717.730 ;
        RECT 1195.640 717.410 1195.900 717.730 ;
        RECT 1195.700 710.590 1195.840 717.410 ;
        RECT 1195.640 710.270 1195.900 710.590 ;
        RECT 1195.640 662.330 1195.900 662.650 ;
        RECT 1195.700 545.690 1195.840 662.330 ;
        RECT 1195.640 545.370 1195.900 545.690 ;
        RECT 1194.720 544.350 1194.980 544.670 ;
        RECT 1194.780 500.470 1194.920 544.350 ;
        RECT 1194.720 500.150 1194.980 500.470 ;
        RECT 1195.640 500.150 1195.900 500.470 ;
        RECT 1195.700 289.670 1195.840 500.150 ;
        RECT 1195.640 289.350 1195.900 289.670 ;
        RECT 1195.180 255.010 1195.440 255.330 ;
        RECT 1195.240 241.390 1195.380 255.010 ;
        RECT 1195.180 241.070 1195.440 241.390 ;
        RECT 1195.640 241.070 1195.900 241.390 ;
        RECT 1195.700 131.230 1195.840 241.070 ;
        RECT 1195.640 130.910 1195.900 131.230 ;
        RECT 1195.180 41.490 1195.440 41.810 ;
        RECT 1195.240 39.090 1195.380 41.490 ;
        RECT 133.500 38.770 133.760 39.090 ;
        RECT 1195.180 38.770 1195.440 39.090 ;
        RECT 133.560 2.400 133.700 38.770 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 1195.170 1483.280 1195.450 1483.560 ;
        RECT 1196.550 1483.280 1196.830 1483.560 ;
        RECT 1195.630 1200.400 1195.910 1200.680 ;
        RECT 1196.090 1199.720 1196.370 1200.000 ;
        RECT 1195.630 1103.840 1195.910 1104.120 ;
        RECT 1195.170 1103.160 1195.450 1103.440 ;
        RECT 1195.630 820.960 1195.910 821.240 ;
        RECT 1196.550 820.960 1196.830 821.240 ;
      LAYER met3 ;
        RECT 1195.145 1483.570 1195.475 1483.585 ;
        RECT 1196.525 1483.570 1196.855 1483.585 ;
        RECT 1195.145 1483.270 1196.855 1483.570 ;
        RECT 1195.145 1483.255 1195.475 1483.270 ;
        RECT 1196.525 1483.255 1196.855 1483.270 ;
        RECT 1195.605 1200.690 1195.935 1200.705 ;
        RECT 1195.390 1200.375 1195.935 1200.690 ;
        RECT 1195.390 1200.010 1195.690 1200.375 ;
        RECT 1196.065 1200.010 1196.395 1200.025 ;
        RECT 1195.390 1199.710 1196.395 1200.010 ;
        RECT 1196.065 1199.695 1196.395 1199.710 ;
        RECT 1195.605 1104.130 1195.935 1104.145 ;
        RECT 1195.390 1103.815 1195.935 1104.130 ;
        RECT 1195.390 1103.465 1195.690 1103.815 ;
        RECT 1195.145 1103.150 1195.690 1103.465 ;
        RECT 1195.145 1103.135 1195.475 1103.150 ;
        RECT 1195.605 821.250 1195.935 821.265 ;
        RECT 1196.525 821.250 1196.855 821.265 ;
        RECT 1195.605 820.950 1196.855 821.250 ;
        RECT 1195.605 820.935 1195.935 820.950 ;
        RECT 1196.525 820.935 1196.855 820.950 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1202.125 1442.025 1202.295 1490.475 ;
        RECT 1202.125 965.685 1202.295 1007.335 ;
        RECT 1202.125 766.445 1202.295 773.075 ;
        RECT 1201.665 717.825 1201.835 765.935 ;
        RECT 1201.665 662.405 1201.835 710.515 ;
        RECT 1201.665 524.365 1201.835 613.955 ;
        RECT 1202.585 421.005 1202.755 469.115 ;
        RECT 1202.585 331.585 1202.755 379.355 ;
        RECT 1201.665 276.165 1201.835 324.275 ;
        RECT 1201.205 41.565 1201.375 89.675 ;
      LAYER mcon ;
        RECT 1202.125 1490.305 1202.295 1490.475 ;
        RECT 1202.125 1007.165 1202.295 1007.335 ;
        RECT 1202.125 772.905 1202.295 773.075 ;
        RECT 1201.665 765.765 1201.835 765.935 ;
        RECT 1201.665 710.345 1201.835 710.515 ;
        RECT 1201.665 613.785 1201.835 613.955 ;
        RECT 1202.585 468.945 1202.755 469.115 ;
        RECT 1202.585 379.185 1202.755 379.355 ;
        RECT 1201.665 324.105 1201.835 324.275 ;
        RECT 1201.205 89.505 1201.375 89.675 ;
      LAYER met1 ;
        RECT 1202.050 1635.640 1202.370 1635.700 ;
        RECT 1204.350 1635.640 1204.670 1635.700 ;
        RECT 1202.050 1635.500 1204.670 1635.640 ;
        RECT 1202.050 1635.440 1202.370 1635.500 ;
        RECT 1204.350 1635.440 1204.670 1635.500 ;
        RECT 1202.050 1490.460 1202.370 1490.520 ;
        RECT 1201.855 1490.320 1202.370 1490.460 ;
        RECT 1202.050 1490.260 1202.370 1490.320 ;
        RECT 1202.050 1442.180 1202.370 1442.240 ;
        RECT 1201.855 1442.040 1202.370 1442.180 ;
        RECT 1202.050 1441.980 1202.370 1442.040 ;
        RECT 1201.130 1345.620 1201.450 1345.680 ;
        RECT 1202.050 1345.620 1202.370 1345.680 ;
        RECT 1201.130 1345.480 1202.370 1345.620 ;
        RECT 1201.130 1345.420 1201.450 1345.480 ;
        RECT 1202.050 1345.420 1202.370 1345.480 ;
        RECT 1201.130 1249.060 1201.450 1249.120 ;
        RECT 1202.050 1249.060 1202.370 1249.120 ;
        RECT 1201.130 1248.920 1202.370 1249.060 ;
        RECT 1201.130 1248.860 1201.450 1248.920 ;
        RECT 1202.050 1248.860 1202.370 1248.920 ;
        RECT 1201.130 1152.500 1201.450 1152.560 ;
        RECT 1202.050 1152.500 1202.370 1152.560 ;
        RECT 1201.130 1152.360 1202.370 1152.500 ;
        RECT 1201.130 1152.300 1201.450 1152.360 ;
        RECT 1202.050 1152.300 1202.370 1152.360 ;
        RECT 1202.050 1007.320 1202.370 1007.380 ;
        RECT 1201.855 1007.180 1202.370 1007.320 ;
        RECT 1202.050 1007.120 1202.370 1007.180 ;
        RECT 1202.065 965.840 1202.355 965.885 ;
        RECT 1202.510 965.840 1202.830 965.900 ;
        RECT 1202.065 965.700 1202.830 965.840 ;
        RECT 1202.065 965.655 1202.355 965.700 ;
        RECT 1202.510 965.640 1202.830 965.700 ;
        RECT 1202.050 869.620 1202.370 869.680 ;
        RECT 1202.510 869.620 1202.830 869.680 ;
        RECT 1202.050 869.480 1202.830 869.620 ;
        RECT 1202.050 869.420 1202.370 869.480 ;
        RECT 1202.510 869.420 1202.830 869.480 ;
        RECT 1202.065 773.060 1202.355 773.105 ;
        RECT 1202.510 773.060 1202.830 773.120 ;
        RECT 1202.065 772.920 1202.830 773.060 ;
        RECT 1202.065 772.875 1202.355 772.920 ;
        RECT 1202.510 772.860 1202.830 772.920 ;
        RECT 1202.050 766.600 1202.370 766.660 ;
        RECT 1201.855 766.460 1202.370 766.600 ;
        RECT 1202.050 766.400 1202.370 766.460 ;
        RECT 1201.605 765.920 1201.895 765.965 ;
        RECT 1202.050 765.920 1202.370 765.980 ;
        RECT 1201.605 765.780 1202.370 765.920 ;
        RECT 1201.605 765.735 1201.895 765.780 ;
        RECT 1202.050 765.720 1202.370 765.780 ;
        RECT 1201.590 717.980 1201.910 718.040 ;
        RECT 1201.395 717.840 1201.910 717.980 ;
        RECT 1201.590 717.780 1201.910 717.840 ;
        RECT 1201.590 710.500 1201.910 710.560 ;
        RECT 1201.395 710.360 1201.910 710.500 ;
        RECT 1201.590 710.300 1201.910 710.360 ;
        RECT 1201.605 662.560 1201.895 662.605 ;
        RECT 1202.050 662.560 1202.370 662.620 ;
        RECT 1201.605 662.420 1202.370 662.560 ;
        RECT 1201.605 662.375 1201.895 662.420 ;
        RECT 1202.050 662.360 1202.370 662.420 ;
        RECT 1201.605 613.940 1201.895 613.985 ;
        RECT 1202.050 613.940 1202.370 614.000 ;
        RECT 1201.605 613.800 1202.370 613.940 ;
        RECT 1201.605 613.755 1201.895 613.800 ;
        RECT 1202.050 613.740 1202.370 613.800 ;
        RECT 1201.590 524.520 1201.910 524.580 ;
        RECT 1201.395 524.380 1201.910 524.520 ;
        RECT 1201.590 524.320 1201.910 524.380 ;
        RECT 1202.050 475.900 1202.370 475.960 ;
        RECT 1202.510 475.900 1202.830 475.960 ;
        RECT 1202.050 475.760 1202.830 475.900 ;
        RECT 1202.050 475.700 1202.370 475.760 ;
        RECT 1202.510 475.700 1202.830 475.760 ;
        RECT 1202.510 469.100 1202.830 469.160 ;
        RECT 1202.315 468.960 1202.830 469.100 ;
        RECT 1202.510 468.900 1202.830 468.960 ;
        RECT 1202.050 421.160 1202.370 421.220 ;
        RECT 1202.525 421.160 1202.815 421.205 ;
        RECT 1202.050 421.020 1202.815 421.160 ;
        RECT 1202.050 420.960 1202.370 421.020 ;
        RECT 1202.525 420.975 1202.815 421.020 ;
        RECT 1202.050 379.340 1202.370 379.400 ;
        RECT 1202.525 379.340 1202.815 379.385 ;
        RECT 1202.050 379.200 1202.815 379.340 ;
        RECT 1202.050 379.140 1202.370 379.200 ;
        RECT 1202.525 379.155 1202.815 379.200 ;
        RECT 1202.050 331.740 1202.370 331.800 ;
        RECT 1202.525 331.740 1202.815 331.785 ;
        RECT 1202.050 331.600 1202.815 331.740 ;
        RECT 1202.050 331.540 1202.370 331.600 ;
        RECT 1202.525 331.555 1202.815 331.600 ;
        RECT 1201.605 324.260 1201.895 324.305 ;
        RECT 1202.050 324.260 1202.370 324.320 ;
        RECT 1201.605 324.120 1202.370 324.260 ;
        RECT 1201.605 324.075 1201.895 324.120 ;
        RECT 1202.050 324.060 1202.370 324.120 ;
        RECT 1201.590 276.320 1201.910 276.380 ;
        RECT 1201.395 276.180 1201.910 276.320 ;
        RECT 1201.590 276.120 1201.910 276.180 ;
        RECT 1201.590 241.640 1201.910 241.700 ;
        RECT 1202.050 241.640 1202.370 241.700 ;
        RECT 1201.590 241.500 1202.370 241.640 ;
        RECT 1201.590 241.440 1201.910 241.500 ;
        RECT 1202.050 241.440 1202.370 241.500 ;
        RECT 1201.145 89.660 1201.435 89.705 ;
        RECT 1201.590 89.660 1201.910 89.720 ;
        RECT 1201.145 89.520 1201.910 89.660 ;
        RECT 1201.145 89.475 1201.435 89.520 ;
        RECT 1201.590 89.460 1201.910 89.520 ;
        RECT 1201.130 41.720 1201.450 41.780 ;
        RECT 1200.935 41.580 1201.450 41.720 ;
        RECT 1201.130 41.520 1201.450 41.580 ;
        RECT 151.410 39.340 151.730 39.400 ;
        RECT 1201.130 39.340 1201.450 39.400 ;
        RECT 151.410 39.200 1201.450 39.340 ;
        RECT 151.410 39.140 151.730 39.200 ;
        RECT 1201.130 39.140 1201.450 39.200 ;
      LAYER via ;
        RECT 1202.080 1635.440 1202.340 1635.700 ;
        RECT 1204.380 1635.440 1204.640 1635.700 ;
        RECT 1202.080 1490.260 1202.340 1490.520 ;
        RECT 1202.080 1441.980 1202.340 1442.240 ;
        RECT 1201.160 1345.420 1201.420 1345.680 ;
        RECT 1202.080 1345.420 1202.340 1345.680 ;
        RECT 1201.160 1248.860 1201.420 1249.120 ;
        RECT 1202.080 1248.860 1202.340 1249.120 ;
        RECT 1201.160 1152.300 1201.420 1152.560 ;
        RECT 1202.080 1152.300 1202.340 1152.560 ;
        RECT 1202.080 1007.120 1202.340 1007.380 ;
        RECT 1202.540 965.640 1202.800 965.900 ;
        RECT 1202.080 869.420 1202.340 869.680 ;
        RECT 1202.540 869.420 1202.800 869.680 ;
        RECT 1202.540 772.860 1202.800 773.120 ;
        RECT 1202.080 766.400 1202.340 766.660 ;
        RECT 1202.080 765.720 1202.340 765.980 ;
        RECT 1201.620 717.780 1201.880 718.040 ;
        RECT 1201.620 710.300 1201.880 710.560 ;
        RECT 1202.080 662.360 1202.340 662.620 ;
        RECT 1202.080 613.740 1202.340 614.000 ;
        RECT 1201.620 524.320 1201.880 524.580 ;
        RECT 1202.080 475.700 1202.340 475.960 ;
        RECT 1202.540 475.700 1202.800 475.960 ;
        RECT 1202.540 468.900 1202.800 469.160 ;
        RECT 1202.080 420.960 1202.340 421.220 ;
        RECT 1202.080 379.140 1202.340 379.400 ;
        RECT 1202.080 331.540 1202.340 331.800 ;
        RECT 1202.080 324.060 1202.340 324.320 ;
        RECT 1201.620 276.120 1201.880 276.380 ;
        RECT 1201.620 241.440 1201.880 241.700 ;
        RECT 1202.080 241.440 1202.340 241.700 ;
        RECT 1201.620 89.460 1201.880 89.720 ;
        RECT 1201.160 41.520 1201.420 41.780 ;
        RECT 151.440 39.140 151.700 39.400 ;
        RECT 1201.160 39.140 1201.420 39.400 ;
      LAYER met2 ;
        RECT 1205.685 1700.410 1205.965 1704.000 ;
        RECT 1204.440 1700.270 1205.965 1700.410 ;
        RECT 1204.440 1635.730 1204.580 1700.270 ;
        RECT 1205.685 1700.000 1205.965 1700.270 ;
        RECT 1202.080 1635.410 1202.340 1635.730 ;
        RECT 1204.380 1635.410 1204.640 1635.730 ;
        RECT 1202.140 1490.550 1202.280 1635.410 ;
        RECT 1202.080 1490.230 1202.340 1490.550 ;
        RECT 1202.080 1441.950 1202.340 1442.270 ;
        RECT 1202.140 1393.845 1202.280 1441.950 ;
        RECT 1201.150 1393.475 1201.430 1393.845 ;
        RECT 1202.070 1393.475 1202.350 1393.845 ;
        RECT 1201.220 1345.710 1201.360 1393.475 ;
        RECT 1201.160 1345.390 1201.420 1345.710 ;
        RECT 1202.080 1345.390 1202.340 1345.710 ;
        RECT 1202.140 1297.285 1202.280 1345.390 ;
        RECT 1201.150 1296.915 1201.430 1297.285 ;
        RECT 1202.070 1296.915 1202.350 1297.285 ;
        RECT 1201.220 1249.150 1201.360 1296.915 ;
        RECT 1201.160 1248.830 1201.420 1249.150 ;
        RECT 1202.080 1248.830 1202.340 1249.150 ;
        RECT 1202.140 1200.725 1202.280 1248.830 ;
        RECT 1201.150 1200.355 1201.430 1200.725 ;
        RECT 1202.070 1200.355 1202.350 1200.725 ;
        RECT 1201.220 1152.590 1201.360 1200.355 ;
        RECT 1201.160 1152.270 1201.420 1152.590 ;
        RECT 1202.080 1152.270 1202.340 1152.590 ;
        RECT 1202.140 1104.165 1202.280 1152.270 ;
        RECT 1201.150 1103.795 1201.430 1104.165 ;
        RECT 1202.070 1103.795 1202.350 1104.165 ;
        RECT 1201.220 1055.885 1201.360 1103.795 ;
        RECT 1201.150 1055.515 1201.430 1055.885 ;
        RECT 1202.070 1055.515 1202.350 1055.885 ;
        RECT 1202.140 1007.410 1202.280 1055.515 ;
        RECT 1202.080 1007.090 1202.340 1007.410 ;
        RECT 1202.540 965.610 1202.800 965.930 ;
        RECT 1202.600 869.710 1202.740 965.610 ;
        RECT 1202.080 869.565 1202.340 869.710 ;
        RECT 1202.070 869.195 1202.350 869.565 ;
        RECT 1202.540 869.390 1202.800 869.710 ;
        RECT 1202.990 869.195 1203.270 869.565 ;
        RECT 1203.060 821.170 1203.200 869.195 ;
        RECT 1202.600 821.030 1203.200 821.170 ;
        RECT 1202.600 773.150 1202.740 821.030 ;
        RECT 1202.540 772.830 1202.800 773.150 ;
        RECT 1202.080 766.370 1202.340 766.690 ;
        RECT 1202.140 766.010 1202.280 766.370 ;
        RECT 1202.080 765.690 1202.340 766.010 ;
        RECT 1201.620 717.750 1201.880 718.070 ;
        RECT 1201.680 710.590 1201.820 717.750 ;
        RECT 1201.620 710.270 1201.880 710.590 ;
        RECT 1202.080 662.330 1202.340 662.650 ;
        RECT 1202.140 614.030 1202.280 662.330 ;
        RECT 1202.080 613.710 1202.340 614.030 ;
        RECT 1201.620 524.290 1201.880 524.610 ;
        RECT 1201.680 524.010 1201.820 524.290 ;
        RECT 1201.680 523.870 1202.740 524.010 ;
        RECT 1202.600 496.130 1202.740 523.870 ;
        RECT 1202.140 495.990 1202.740 496.130 ;
        RECT 1202.140 475.990 1202.280 495.990 ;
        RECT 1202.080 475.670 1202.340 475.990 ;
        RECT 1202.540 475.670 1202.800 475.990 ;
        RECT 1202.600 469.190 1202.740 475.670 ;
        RECT 1202.540 468.870 1202.800 469.190 ;
        RECT 1202.080 420.930 1202.340 421.250 ;
        RECT 1202.140 379.430 1202.280 420.930 ;
        RECT 1202.080 379.110 1202.340 379.430 ;
        RECT 1202.080 331.510 1202.340 331.830 ;
        RECT 1202.140 324.350 1202.280 331.510 ;
        RECT 1202.080 324.030 1202.340 324.350 ;
        RECT 1201.620 276.090 1201.880 276.410 ;
        RECT 1201.680 241.730 1201.820 276.090 ;
        RECT 1201.620 241.410 1201.880 241.730 ;
        RECT 1202.080 241.410 1202.340 241.730 ;
        RECT 1202.140 90.965 1202.280 241.410 ;
        RECT 1202.070 90.595 1202.350 90.965 ;
        RECT 1201.610 89.915 1201.890 90.285 ;
        RECT 1201.680 89.750 1201.820 89.915 ;
        RECT 1201.620 89.430 1201.880 89.750 ;
        RECT 1201.160 41.490 1201.420 41.810 ;
        RECT 1201.220 39.430 1201.360 41.490 ;
        RECT 151.440 39.110 151.700 39.430 ;
        RECT 1201.160 39.110 1201.420 39.430 ;
        RECT 151.500 2.400 151.640 39.110 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1201.150 1393.520 1201.430 1393.800 ;
        RECT 1202.070 1393.520 1202.350 1393.800 ;
        RECT 1201.150 1296.960 1201.430 1297.240 ;
        RECT 1202.070 1296.960 1202.350 1297.240 ;
        RECT 1201.150 1200.400 1201.430 1200.680 ;
        RECT 1202.070 1200.400 1202.350 1200.680 ;
        RECT 1201.150 1103.840 1201.430 1104.120 ;
        RECT 1202.070 1103.840 1202.350 1104.120 ;
        RECT 1201.150 1055.560 1201.430 1055.840 ;
        RECT 1202.070 1055.560 1202.350 1055.840 ;
        RECT 1202.070 869.240 1202.350 869.520 ;
        RECT 1202.990 869.240 1203.270 869.520 ;
        RECT 1202.070 90.640 1202.350 90.920 ;
        RECT 1201.610 89.960 1201.890 90.240 ;
      LAYER met3 ;
        RECT 1201.125 1393.810 1201.455 1393.825 ;
        RECT 1202.045 1393.810 1202.375 1393.825 ;
        RECT 1201.125 1393.510 1202.375 1393.810 ;
        RECT 1201.125 1393.495 1201.455 1393.510 ;
        RECT 1202.045 1393.495 1202.375 1393.510 ;
        RECT 1201.125 1297.250 1201.455 1297.265 ;
        RECT 1202.045 1297.250 1202.375 1297.265 ;
        RECT 1201.125 1296.950 1202.375 1297.250 ;
        RECT 1201.125 1296.935 1201.455 1296.950 ;
        RECT 1202.045 1296.935 1202.375 1296.950 ;
        RECT 1201.125 1200.690 1201.455 1200.705 ;
        RECT 1202.045 1200.690 1202.375 1200.705 ;
        RECT 1201.125 1200.390 1202.375 1200.690 ;
        RECT 1201.125 1200.375 1201.455 1200.390 ;
        RECT 1202.045 1200.375 1202.375 1200.390 ;
        RECT 1201.125 1104.130 1201.455 1104.145 ;
        RECT 1202.045 1104.130 1202.375 1104.145 ;
        RECT 1201.125 1103.830 1202.375 1104.130 ;
        RECT 1201.125 1103.815 1201.455 1103.830 ;
        RECT 1202.045 1103.815 1202.375 1103.830 ;
        RECT 1201.125 1055.850 1201.455 1055.865 ;
        RECT 1202.045 1055.850 1202.375 1055.865 ;
        RECT 1201.125 1055.550 1202.375 1055.850 ;
        RECT 1201.125 1055.535 1201.455 1055.550 ;
        RECT 1202.045 1055.535 1202.375 1055.550 ;
        RECT 1202.045 869.530 1202.375 869.545 ;
        RECT 1202.965 869.530 1203.295 869.545 ;
        RECT 1202.045 869.230 1203.295 869.530 ;
        RECT 1202.045 869.215 1202.375 869.230 ;
        RECT 1202.965 869.215 1203.295 869.230 ;
        RECT 1202.045 90.930 1202.375 90.945 ;
        RECT 1200.910 90.630 1202.375 90.930 ;
        RECT 1200.910 90.250 1201.210 90.630 ;
        RECT 1202.045 90.615 1202.375 90.630 ;
        RECT 1201.585 90.250 1201.915 90.265 ;
        RECT 1200.910 89.950 1201.915 90.250 ;
        RECT 1201.585 89.935 1201.915 89.950 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1209.485 1442.025 1209.655 1490.475 ;
        RECT 1209.025 869.465 1209.195 894.115 ;
        RECT 1209.485 766.105 1209.655 814.215 ;
        RECT 1209.485 628.065 1209.655 676.175 ;
        RECT 1209.485 572.645 1209.655 620.755 ;
        RECT 1209.025 476.085 1209.195 524.195 ;
        RECT 1209.025 144.925 1209.195 220.575 ;
        RECT 1208.105 41.565 1208.275 89.675 ;
      LAYER mcon ;
        RECT 1209.485 1490.305 1209.655 1490.475 ;
        RECT 1209.025 893.945 1209.195 894.115 ;
        RECT 1209.485 814.045 1209.655 814.215 ;
        RECT 1209.485 676.005 1209.655 676.175 ;
        RECT 1209.485 620.585 1209.655 620.755 ;
        RECT 1209.025 524.025 1209.195 524.195 ;
        RECT 1209.025 220.405 1209.195 220.575 ;
        RECT 1208.105 89.505 1208.275 89.675 ;
      LAYER met1 ;
        RECT 1209.410 1635.640 1209.730 1635.700 ;
        RECT 1210.790 1635.640 1211.110 1635.700 ;
        RECT 1209.410 1635.500 1211.110 1635.640 ;
        RECT 1209.410 1635.440 1209.730 1635.500 ;
        RECT 1210.790 1635.440 1211.110 1635.500 ;
        RECT 1209.410 1490.460 1209.730 1490.520 ;
        RECT 1209.215 1490.320 1209.730 1490.460 ;
        RECT 1209.410 1490.260 1209.730 1490.320 ;
        RECT 1209.410 1442.180 1209.730 1442.240 ;
        RECT 1209.215 1442.040 1209.730 1442.180 ;
        RECT 1209.410 1441.980 1209.730 1442.040 ;
        RECT 1209.410 1345.620 1209.730 1345.680 ;
        RECT 1210.330 1345.620 1210.650 1345.680 ;
        RECT 1209.410 1345.480 1210.650 1345.620 ;
        RECT 1209.410 1345.420 1209.730 1345.480 ;
        RECT 1210.330 1345.420 1210.650 1345.480 ;
        RECT 1209.410 1249.060 1209.730 1249.120 ;
        RECT 1210.330 1249.060 1210.650 1249.120 ;
        RECT 1209.410 1248.920 1210.650 1249.060 ;
        RECT 1209.410 1248.860 1209.730 1248.920 ;
        RECT 1210.330 1248.860 1210.650 1248.920 ;
        RECT 1209.410 1152.500 1209.730 1152.560 ;
        RECT 1210.330 1152.500 1210.650 1152.560 ;
        RECT 1209.410 1152.360 1210.650 1152.500 ;
        RECT 1209.410 1152.300 1209.730 1152.360 ;
        RECT 1210.330 1152.300 1210.650 1152.360 ;
        RECT 1209.410 918.240 1209.730 918.300 ;
        RECT 1209.040 918.100 1209.730 918.240 ;
        RECT 1209.040 917.960 1209.180 918.100 ;
        RECT 1209.410 918.040 1209.730 918.100 ;
        RECT 1208.950 917.700 1209.270 917.960 ;
        RECT 1208.950 894.100 1209.270 894.160 ;
        RECT 1208.755 893.960 1209.270 894.100 ;
        RECT 1208.950 893.900 1209.270 893.960 ;
        RECT 1208.950 869.620 1209.270 869.680 ;
        RECT 1208.755 869.480 1209.270 869.620 ;
        RECT 1208.950 869.420 1209.270 869.480 ;
        RECT 1209.410 814.200 1209.730 814.260 ;
        RECT 1209.215 814.060 1209.730 814.200 ;
        RECT 1209.410 814.000 1209.730 814.060 ;
        RECT 1209.410 766.260 1209.730 766.320 ;
        RECT 1209.215 766.120 1209.730 766.260 ;
        RECT 1209.410 766.060 1209.730 766.120 ;
        RECT 1208.950 724.440 1209.270 724.500 ;
        RECT 1209.870 724.440 1210.190 724.500 ;
        RECT 1208.950 724.300 1210.190 724.440 ;
        RECT 1208.950 724.240 1209.270 724.300 ;
        RECT 1209.870 724.240 1210.190 724.300 ;
        RECT 1209.410 676.160 1209.730 676.220 ;
        RECT 1209.215 676.020 1209.730 676.160 ;
        RECT 1209.410 675.960 1209.730 676.020 ;
        RECT 1209.410 628.220 1209.730 628.280 ;
        RECT 1209.215 628.080 1209.730 628.220 ;
        RECT 1209.410 628.020 1209.730 628.080 ;
        RECT 1209.410 620.740 1209.730 620.800 ;
        RECT 1209.215 620.600 1209.730 620.740 ;
        RECT 1209.410 620.540 1209.730 620.600 ;
        RECT 1209.410 572.800 1209.730 572.860 ;
        RECT 1209.215 572.660 1209.730 572.800 ;
        RECT 1209.410 572.600 1209.730 572.660 ;
        RECT 1208.030 555.460 1208.350 555.520 ;
        RECT 1209.410 555.460 1209.730 555.520 ;
        RECT 1208.030 555.320 1209.730 555.460 ;
        RECT 1208.030 555.260 1208.350 555.320 ;
        RECT 1209.410 555.260 1209.730 555.320 ;
        RECT 1208.950 524.180 1209.270 524.240 ;
        RECT 1208.755 524.040 1209.270 524.180 ;
        RECT 1208.950 523.980 1209.270 524.040 ;
        RECT 1208.965 476.240 1209.255 476.285 ;
        RECT 1209.410 476.240 1209.730 476.300 ;
        RECT 1208.965 476.100 1209.730 476.240 ;
        RECT 1208.965 476.055 1209.255 476.100 ;
        RECT 1209.410 476.040 1209.730 476.100 ;
        RECT 1208.950 220.560 1209.270 220.620 ;
        RECT 1208.755 220.420 1209.270 220.560 ;
        RECT 1208.950 220.360 1209.270 220.420 ;
        RECT 1208.950 145.080 1209.270 145.140 ;
        RECT 1208.755 144.940 1209.270 145.080 ;
        RECT 1208.950 144.880 1209.270 144.940 ;
        RECT 1208.030 89.660 1208.350 89.720 ;
        RECT 1207.835 89.520 1208.350 89.660 ;
        RECT 1208.030 89.460 1208.350 89.520 ;
        RECT 1208.045 41.720 1208.335 41.765 ;
        RECT 1208.490 41.720 1208.810 41.780 ;
        RECT 1208.045 41.580 1208.810 41.720 ;
        RECT 1208.045 41.535 1208.335 41.580 ;
        RECT 1208.490 41.520 1208.810 41.580 ;
        RECT 169.350 39.680 169.670 39.740 ;
        RECT 1208.490 39.680 1208.810 39.740 ;
        RECT 169.350 39.540 1208.810 39.680 ;
        RECT 169.350 39.480 169.670 39.540 ;
        RECT 1208.490 39.480 1208.810 39.540 ;
      LAYER via ;
        RECT 1209.440 1635.440 1209.700 1635.700 ;
        RECT 1210.820 1635.440 1211.080 1635.700 ;
        RECT 1209.440 1490.260 1209.700 1490.520 ;
        RECT 1209.440 1441.980 1209.700 1442.240 ;
        RECT 1209.440 1345.420 1209.700 1345.680 ;
        RECT 1210.360 1345.420 1210.620 1345.680 ;
        RECT 1209.440 1248.860 1209.700 1249.120 ;
        RECT 1210.360 1248.860 1210.620 1249.120 ;
        RECT 1209.440 1152.300 1209.700 1152.560 ;
        RECT 1210.360 1152.300 1210.620 1152.560 ;
        RECT 1209.440 918.040 1209.700 918.300 ;
        RECT 1208.980 917.700 1209.240 917.960 ;
        RECT 1208.980 893.900 1209.240 894.160 ;
        RECT 1208.980 869.420 1209.240 869.680 ;
        RECT 1209.440 814.000 1209.700 814.260 ;
        RECT 1209.440 766.060 1209.700 766.320 ;
        RECT 1208.980 724.240 1209.240 724.500 ;
        RECT 1209.900 724.240 1210.160 724.500 ;
        RECT 1209.440 675.960 1209.700 676.220 ;
        RECT 1209.440 628.020 1209.700 628.280 ;
        RECT 1209.440 620.540 1209.700 620.800 ;
        RECT 1209.440 572.600 1209.700 572.860 ;
        RECT 1208.060 555.260 1208.320 555.520 ;
        RECT 1209.440 555.260 1209.700 555.520 ;
        RECT 1208.980 523.980 1209.240 524.240 ;
        RECT 1209.440 476.040 1209.700 476.300 ;
        RECT 1208.980 220.360 1209.240 220.620 ;
        RECT 1208.980 144.880 1209.240 145.140 ;
        RECT 1208.060 89.460 1208.320 89.720 ;
        RECT 1208.520 41.520 1208.780 41.780 ;
        RECT 169.380 39.480 169.640 39.740 ;
        RECT 1208.520 39.480 1208.780 39.740 ;
      LAYER met2 ;
        RECT 1212.585 1700.410 1212.865 1704.000 ;
        RECT 1210.880 1700.270 1212.865 1700.410 ;
        RECT 1210.880 1635.730 1211.020 1700.270 ;
        RECT 1212.585 1700.000 1212.865 1700.270 ;
        RECT 1209.440 1635.410 1209.700 1635.730 ;
        RECT 1210.820 1635.410 1211.080 1635.730 ;
        RECT 1209.500 1490.550 1209.640 1635.410 ;
        RECT 1209.440 1490.230 1209.700 1490.550 ;
        RECT 1209.440 1441.950 1209.700 1442.270 ;
        RECT 1209.500 1393.845 1209.640 1441.950 ;
        RECT 1209.430 1393.475 1209.710 1393.845 ;
        RECT 1210.350 1393.475 1210.630 1393.845 ;
        RECT 1210.420 1345.710 1210.560 1393.475 ;
        RECT 1209.440 1345.390 1209.700 1345.710 ;
        RECT 1210.360 1345.390 1210.620 1345.710 ;
        RECT 1209.500 1297.285 1209.640 1345.390 ;
        RECT 1209.430 1296.915 1209.710 1297.285 ;
        RECT 1210.350 1296.915 1210.630 1297.285 ;
        RECT 1210.420 1249.150 1210.560 1296.915 ;
        RECT 1209.440 1248.830 1209.700 1249.150 ;
        RECT 1210.360 1248.830 1210.620 1249.150 ;
        RECT 1209.500 1200.725 1209.640 1248.830 ;
        RECT 1209.430 1200.355 1209.710 1200.725 ;
        RECT 1210.350 1200.355 1210.630 1200.725 ;
        RECT 1210.420 1152.590 1210.560 1200.355 ;
        RECT 1209.440 1152.270 1209.700 1152.590 ;
        RECT 1210.360 1152.270 1210.620 1152.590 ;
        RECT 1209.500 1104.165 1209.640 1152.270 ;
        RECT 1209.430 1103.795 1209.710 1104.165 ;
        RECT 1210.350 1103.795 1210.630 1104.165 ;
        RECT 1210.420 1055.885 1210.560 1103.795 ;
        RECT 1209.430 1055.515 1209.710 1055.885 ;
        RECT 1210.350 1055.515 1210.630 1055.885 ;
        RECT 1209.500 918.330 1209.640 1055.515 ;
        RECT 1209.440 918.010 1209.700 918.330 ;
        RECT 1208.980 917.670 1209.240 917.990 ;
        RECT 1209.040 894.190 1209.180 917.670 ;
        RECT 1208.980 893.870 1209.240 894.190 ;
        RECT 1208.980 869.390 1209.240 869.710 ;
        RECT 1209.040 821.170 1209.180 869.390 ;
        RECT 1209.040 821.030 1209.640 821.170 ;
        RECT 1209.500 814.290 1209.640 821.030 ;
        RECT 1209.440 813.970 1209.700 814.290 ;
        RECT 1209.440 766.030 1209.700 766.350 ;
        RECT 1209.500 738.210 1209.640 766.030 ;
        RECT 1209.040 738.070 1209.640 738.210 ;
        RECT 1209.040 724.530 1209.180 738.070 ;
        RECT 1208.980 724.210 1209.240 724.530 ;
        RECT 1209.900 724.210 1210.160 724.530 ;
        RECT 1209.960 676.330 1210.100 724.210 ;
        RECT 1209.500 676.250 1210.100 676.330 ;
        RECT 1209.440 676.190 1210.100 676.250 ;
        RECT 1209.440 675.930 1209.700 676.190 ;
        RECT 1209.500 675.775 1209.640 675.930 ;
        RECT 1209.440 627.990 1209.700 628.310 ;
        RECT 1209.500 620.830 1209.640 627.990 ;
        RECT 1209.440 620.510 1209.700 620.830 ;
        RECT 1209.440 572.570 1209.700 572.890 ;
        RECT 1209.500 555.550 1209.640 572.570 ;
        RECT 1208.060 555.230 1208.320 555.550 ;
        RECT 1209.440 555.230 1209.700 555.550 ;
        RECT 1208.120 531.605 1208.260 555.230 ;
        RECT 1208.050 531.235 1208.330 531.605 ;
        RECT 1208.970 531.235 1209.250 531.605 ;
        RECT 1209.040 524.270 1209.180 531.235 ;
        RECT 1208.980 523.950 1209.240 524.270 ;
        RECT 1209.440 476.010 1209.700 476.330 ;
        RECT 1209.500 289.410 1209.640 476.010 ;
        RECT 1209.040 289.270 1209.640 289.410 ;
        RECT 1209.040 252.010 1209.180 289.270 ;
        RECT 1209.040 251.870 1209.640 252.010 ;
        RECT 1209.500 228.210 1209.640 251.870 ;
        RECT 1209.040 228.070 1209.640 228.210 ;
        RECT 1209.040 220.650 1209.180 228.070 ;
        RECT 1208.980 220.330 1209.240 220.650 ;
        RECT 1208.980 144.850 1209.240 145.170 ;
        RECT 1209.040 90.965 1209.180 144.850 ;
        RECT 1208.970 90.595 1209.250 90.965 ;
        RECT 1208.050 89.915 1208.330 90.285 ;
        RECT 1208.120 89.750 1208.260 89.915 ;
        RECT 1208.060 89.430 1208.320 89.750 ;
        RECT 1208.520 41.490 1208.780 41.810 ;
        RECT 1208.580 39.770 1208.720 41.490 ;
        RECT 169.380 39.450 169.640 39.770 ;
        RECT 1208.520 39.450 1208.780 39.770 ;
        RECT 169.440 2.400 169.580 39.450 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 1209.430 1393.520 1209.710 1393.800 ;
        RECT 1210.350 1393.520 1210.630 1393.800 ;
        RECT 1209.430 1296.960 1209.710 1297.240 ;
        RECT 1210.350 1296.960 1210.630 1297.240 ;
        RECT 1209.430 1200.400 1209.710 1200.680 ;
        RECT 1210.350 1200.400 1210.630 1200.680 ;
        RECT 1209.430 1103.840 1209.710 1104.120 ;
        RECT 1210.350 1103.840 1210.630 1104.120 ;
        RECT 1209.430 1055.560 1209.710 1055.840 ;
        RECT 1210.350 1055.560 1210.630 1055.840 ;
        RECT 1208.050 531.280 1208.330 531.560 ;
        RECT 1208.970 531.280 1209.250 531.560 ;
        RECT 1208.970 90.640 1209.250 90.920 ;
        RECT 1208.050 89.960 1208.330 90.240 ;
      LAYER met3 ;
        RECT 1209.405 1393.810 1209.735 1393.825 ;
        RECT 1210.325 1393.810 1210.655 1393.825 ;
        RECT 1209.405 1393.510 1210.655 1393.810 ;
        RECT 1209.405 1393.495 1209.735 1393.510 ;
        RECT 1210.325 1393.495 1210.655 1393.510 ;
        RECT 1209.405 1297.250 1209.735 1297.265 ;
        RECT 1210.325 1297.250 1210.655 1297.265 ;
        RECT 1209.405 1296.950 1210.655 1297.250 ;
        RECT 1209.405 1296.935 1209.735 1296.950 ;
        RECT 1210.325 1296.935 1210.655 1296.950 ;
        RECT 1209.405 1200.690 1209.735 1200.705 ;
        RECT 1210.325 1200.690 1210.655 1200.705 ;
        RECT 1209.405 1200.390 1210.655 1200.690 ;
        RECT 1209.405 1200.375 1209.735 1200.390 ;
        RECT 1210.325 1200.375 1210.655 1200.390 ;
        RECT 1209.405 1104.130 1209.735 1104.145 ;
        RECT 1210.325 1104.130 1210.655 1104.145 ;
        RECT 1209.405 1103.830 1210.655 1104.130 ;
        RECT 1209.405 1103.815 1209.735 1103.830 ;
        RECT 1210.325 1103.815 1210.655 1103.830 ;
        RECT 1209.405 1055.850 1209.735 1055.865 ;
        RECT 1210.325 1055.850 1210.655 1055.865 ;
        RECT 1209.405 1055.550 1210.655 1055.850 ;
        RECT 1209.405 1055.535 1209.735 1055.550 ;
        RECT 1210.325 1055.535 1210.655 1055.550 ;
        RECT 1208.025 531.570 1208.355 531.585 ;
        RECT 1208.945 531.570 1209.275 531.585 ;
        RECT 1208.025 531.270 1209.275 531.570 ;
        RECT 1208.025 531.255 1208.355 531.270 ;
        RECT 1208.945 531.255 1209.275 531.270 ;
        RECT 1208.945 90.930 1209.275 90.945 ;
        RECT 1208.040 90.630 1209.275 90.930 ;
        RECT 1208.040 90.265 1208.340 90.630 ;
        RECT 1208.945 90.615 1209.275 90.630 ;
        RECT 1208.025 89.935 1208.355 90.265 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 40.020 187.150 40.080 ;
        RECT 1215.390 40.020 1215.710 40.080 ;
        RECT 186.830 39.880 1215.710 40.020 ;
        RECT 186.830 39.820 187.150 39.880 ;
        RECT 1215.390 39.820 1215.710 39.880 ;
      LAYER via ;
        RECT 186.860 39.820 187.120 40.080 ;
        RECT 1215.420 39.820 1215.680 40.080 ;
      LAYER met2 ;
        RECT 1219.485 1700.410 1219.765 1704.000 ;
        RECT 1217.780 1700.270 1219.765 1700.410 ;
        RECT 1217.780 1678.480 1217.920 1700.270 ;
        RECT 1219.485 1700.000 1219.765 1700.270 ;
        RECT 1215.480 1678.340 1217.920 1678.480 ;
        RECT 1215.480 40.110 1215.620 1678.340 ;
        RECT 186.860 39.790 187.120 40.110 ;
        RECT 1215.420 39.790 1215.680 40.110 ;
        RECT 186.920 2.400 187.060 39.790 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1222.365 427.805 1222.535 473.195 ;
      LAYER mcon ;
        RECT 1222.365 473.025 1222.535 473.195 ;
      LAYER met1 ;
        RECT 1222.290 1158.960 1222.610 1159.020 ;
        RECT 1222.750 1158.960 1223.070 1159.020 ;
        RECT 1222.290 1158.820 1223.070 1158.960 ;
        RECT 1222.290 1158.760 1222.610 1158.820 ;
        RECT 1222.750 1158.760 1223.070 1158.820 ;
        RECT 1222.290 473.180 1222.610 473.240 ;
        RECT 1222.095 473.040 1222.610 473.180 ;
        RECT 1222.290 472.980 1222.610 473.040 ;
        RECT 1222.290 427.960 1222.610 428.020 ;
        RECT 1222.095 427.820 1222.610 427.960 ;
        RECT 1222.290 427.760 1222.610 427.820 ;
        RECT 1222.290 386.480 1222.610 386.540 ;
        RECT 1222.750 386.480 1223.070 386.540 ;
        RECT 1222.290 386.340 1223.070 386.480 ;
        RECT 1222.290 386.280 1222.610 386.340 ;
        RECT 1222.750 386.280 1223.070 386.340 ;
        RECT 1222.290 379.340 1222.610 379.400 ;
        RECT 1222.750 379.340 1223.070 379.400 ;
        RECT 1222.290 379.200 1223.070 379.340 ;
        RECT 1222.290 379.140 1222.610 379.200 ;
        RECT 1222.750 379.140 1223.070 379.200 ;
        RECT 1222.750 97.140 1223.070 97.200 ;
        RECT 1222.380 97.000 1223.070 97.140 ;
        RECT 1222.380 96.860 1222.520 97.000 ;
        RECT 1222.750 96.940 1223.070 97.000 ;
        RECT 1222.290 96.600 1222.610 96.860 ;
        RECT 204.770 45.460 205.090 45.520 ;
        RECT 1222.290 45.460 1222.610 45.520 ;
        RECT 204.770 45.320 1222.610 45.460 ;
        RECT 204.770 45.260 205.090 45.320 ;
        RECT 1222.290 45.260 1222.610 45.320 ;
      LAYER via ;
        RECT 1222.320 1158.760 1222.580 1159.020 ;
        RECT 1222.780 1158.760 1223.040 1159.020 ;
        RECT 1222.320 472.980 1222.580 473.240 ;
        RECT 1222.320 427.760 1222.580 428.020 ;
        RECT 1222.320 386.280 1222.580 386.540 ;
        RECT 1222.780 386.280 1223.040 386.540 ;
        RECT 1222.320 379.140 1222.580 379.400 ;
        RECT 1222.780 379.140 1223.040 379.400 ;
        RECT 1222.780 96.940 1223.040 97.200 ;
        RECT 1222.320 96.600 1222.580 96.860 ;
        RECT 204.800 45.260 205.060 45.520 ;
        RECT 1222.320 45.260 1222.580 45.520 ;
      LAYER met2 ;
        RECT 1225.925 1700.410 1226.205 1704.000 ;
        RECT 1224.680 1700.270 1226.205 1700.410 ;
        RECT 1224.680 1658.930 1224.820 1700.270 ;
        RECT 1225.925 1700.000 1226.205 1700.270 ;
        RECT 1222.840 1658.790 1224.820 1658.930 ;
        RECT 1222.840 1583.450 1222.980 1658.790 ;
        RECT 1222.380 1583.310 1222.980 1583.450 ;
        RECT 1222.380 1535.170 1222.520 1583.310 ;
        RECT 1222.380 1535.030 1222.980 1535.170 ;
        RECT 1222.840 1486.890 1222.980 1535.030 ;
        RECT 1222.380 1486.750 1222.980 1486.890 ;
        RECT 1222.380 1438.610 1222.520 1486.750 ;
        RECT 1222.380 1438.470 1222.980 1438.610 ;
        RECT 1222.840 1388.970 1222.980 1438.470 ;
        RECT 1222.380 1388.830 1222.980 1388.970 ;
        RECT 1222.380 1352.930 1222.520 1388.830 ;
        RECT 1222.380 1352.790 1222.980 1352.930 ;
        RECT 1222.840 1292.410 1222.980 1352.790 ;
        RECT 1222.380 1292.270 1222.980 1292.410 ;
        RECT 1222.380 1256.370 1222.520 1292.270 ;
        RECT 1222.380 1256.230 1222.980 1256.370 ;
        RECT 1222.840 1197.210 1222.980 1256.230 ;
        RECT 1222.380 1197.070 1222.980 1197.210 ;
        RECT 1222.380 1159.050 1222.520 1197.070 ;
        RECT 1222.320 1158.730 1222.580 1159.050 ;
        RECT 1222.780 1158.730 1223.040 1159.050 ;
        RECT 1222.840 1089.770 1222.980 1158.730 ;
        RECT 1222.380 1089.630 1222.980 1089.770 ;
        RECT 1222.380 1053.730 1222.520 1089.630 ;
        RECT 1222.380 1053.590 1222.980 1053.730 ;
        RECT 1222.840 993.210 1222.980 1053.590 ;
        RECT 1222.380 993.070 1222.980 993.210 ;
        RECT 1222.380 957.170 1222.520 993.070 ;
        RECT 1222.380 957.030 1222.980 957.170 ;
        RECT 1222.840 810.970 1222.980 957.030 ;
        RECT 1222.380 810.830 1222.980 810.970 ;
        RECT 1222.380 762.690 1222.520 810.830 ;
        RECT 1222.380 762.550 1222.980 762.690 ;
        RECT 1222.840 617.850 1222.980 762.550 ;
        RECT 1222.380 617.710 1222.980 617.850 ;
        RECT 1222.380 569.570 1222.520 617.710 ;
        RECT 1222.380 569.430 1222.980 569.570 ;
        RECT 1222.840 521.290 1222.980 569.430 ;
        RECT 1222.380 521.150 1222.980 521.290 ;
        RECT 1222.380 473.270 1222.520 521.150 ;
        RECT 1222.320 472.950 1222.580 473.270 ;
        RECT 1222.320 427.730 1222.580 428.050 ;
        RECT 1222.380 386.570 1222.520 427.730 ;
        RECT 1222.320 386.250 1222.580 386.570 ;
        RECT 1222.780 386.250 1223.040 386.570 ;
        RECT 1222.840 379.430 1222.980 386.250 ;
        RECT 1222.320 379.110 1222.580 379.430 ;
        RECT 1222.780 379.110 1223.040 379.430 ;
        RECT 1222.380 279.210 1222.520 379.110 ;
        RECT 1222.380 279.070 1222.980 279.210 ;
        RECT 1222.840 97.230 1222.980 279.070 ;
        RECT 1222.780 96.910 1223.040 97.230 ;
        RECT 1222.320 96.570 1222.580 96.890 ;
        RECT 1222.380 45.550 1222.520 96.570 ;
        RECT 204.800 45.230 205.060 45.550 ;
        RECT 1222.320 45.230 1222.580 45.550 ;
        RECT 204.860 2.400 205.000 45.230 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1229.725 1304.325 1229.895 1352.435 ;
        RECT 1229.725 1207.425 1229.895 1255.875 ;
        RECT 1229.725 531.505 1229.895 579.615 ;
        RECT 1229.725 241.485 1229.895 289.595 ;
        RECT 1229.725 144.925 1229.895 193.035 ;
      LAYER mcon ;
        RECT 1229.725 1352.265 1229.895 1352.435 ;
        RECT 1229.725 1255.705 1229.895 1255.875 ;
        RECT 1229.725 579.445 1229.895 579.615 ;
        RECT 1229.725 289.425 1229.895 289.595 ;
        RECT 1229.725 192.865 1229.895 193.035 ;
      LAYER met1 ;
        RECT 1229.650 1635.640 1229.970 1635.700 ;
        RECT 1231.030 1635.640 1231.350 1635.700 ;
        RECT 1229.650 1635.500 1231.350 1635.640 ;
        RECT 1229.650 1635.440 1229.970 1635.500 ;
        RECT 1231.030 1635.440 1231.350 1635.500 ;
        RECT 1229.650 1352.420 1229.970 1352.480 ;
        RECT 1229.455 1352.280 1229.970 1352.420 ;
        RECT 1229.650 1352.220 1229.970 1352.280 ;
        RECT 1229.650 1304.480 1229.970 1304.540 ;
        RECT 1229.455 1304.340 1229.970 1304.480 ;
        RECT 1229.650 1304.280 1229.970 1304.340 ;
        RECT 1229.650 1255.860 1229.970 1255.920 ;
        RECT 1229.455 1255.720 1229.970 1255.860 ;
        RECT 1229.650 1255.660 1229.970 1255.720 ;
        RECT 1229.650 1207.580 1229.970 1207.640 ;
        RECT 1229.455 1207.440 1229.970 1207.580 ;
        RECT 1229.650 1207.380 1229.970 1207.440 ;
        RECT 1228.730 1111.020 1229.050 1111.080 ;
        RECT 1229.650 1111.020 1229.970 1111.080 ;
        RECT 1228.730 1110.880 1229.970 1111.020 ;
        RECT 1228.730 1110.820 1229.050 1110.880 ;
        RECT 1229.650 1110.820 1229.970 1110.880 ;
        RECT 1228.730 772.720 1229.050 772.780 ;
        RECT 1229.650 772.720 1229.970 772.780 ;
        RECT 1228.730 772.580 1229.970 772.720 ;
        RECT 1228.730 772.520 1229.050 772.580 ;
        RECT 1229.650 772.520 1229.970 772.580 ;
        RECT 1228.730 676.160 1229.050 676.220 ;
        RECT 1229.650 676.160 1229.970 676.220 ;
        RECT 1228.730 676.020 1229.970 676.160 ;
        RECT 1228.730 675.960 1229.050 676.020 ;
        RECT 1229.650 675.960 1229.970 676.020 ;
        RECT 1229.650 579.600 1229.970 579.660 ;
        RECT 1229.455 579.460 1229.970 579.600 ;
        RECT 1229.650 579.400 1229.970 579.460 ;
        RECT 1229.650 531.660 1229.970 531.720 ;
        RECT 1229.455 531.520 1229.970 531.660 ;
        RECT 1229.650 531.460 1229.970 531.520 ;
        RECT 1229.650 289.580 1229.970 289.640 ;
        RECT 1229.455 289.440 1229.970 289.580 ;
        RECT 1229.650 289.380 1229.970 289.440 ;
        RECT 1229.650 241.640 1229.970 241.700 ;
        RECT 1229.455 241.500 1229.970 241.640 ;
        RECT 1229.650 241.440 1229.970 241.500 ;
        RECT 1229.650 193.020 1229.970 193.080 ;
        RECT 1229.455 192.880 1229.970 193.020 ;
        RECT 1229.650 192.820 1229.970 192.880 ;
        RECT 1229.650 145.080 1229.970 145.140 ;
        RECT 1229.455 144.940 1229.970 145.080 ;
        RECT 1229.650 144.880 1229.970 144.940 ;
        RECT 1229.650 110.740 1229.970 110.800 ;
        RECT 1228.820 110.600 1229.970 110.740 ;
        RECT 1228.820 110.460 1228.960 110.600 ;
        RECT 1229.650 110.540 1229.970 110.600 ;
        RECT 1228.730 110.200 1229.050 110.460 ;
        RECT 222.710 45.800 223.030 45.860 ;
        RECT 1228.730 45.800 1229.050 45.860 ;
        RECT 222.710 45.660 1229.050 45.800 ;
        RECT 222.710 45.600 223.030 45.660 ;
        RECT 1228.730 45.600 1229.050 45.660 ;
      LAYER via ;
        RECT 1229.680 1635.440 1229.940 1635.700 ;
        RECT 1231.060 1635.440 1231.320 1635.700 ;
        RECT 1229.680 1352.220 1229.940 1352.480 ;
        RECT 1229.680 1304.280 1229.940 1304.540 ;
        RECT 1229.680 1255.660 1229.940 1255.920 ;
        RECT 1229.680 1207.380 1229.940 1207.640 ;
        RECT 1228.760 1110.820 1229.020 1111.080 ;
        RECT 1229.680 1110.820 1229.940 1111.080 ;
        RECT 1228.760 772.520 1229.020 772.780 ;
        RECT 1229.680 772.520 1229.940 772.780 ;
        RECT 1228.760 675.960 1229.020 676.220 ;
        RECT 1229.680 675.960 1229.940 676.220 ;
        RECT 1229.680 579.400 1229.940 579.660 ;
        RECT 1229.680 531.460 1229.940 531.720 ;
        RECT 1229.680 289.380 1229.940 289.640 ;
        RECT 1229.680 241.440 1229.940 241.700 ;
        RECT 1229.680 192.820 1229.940 193.080 ;
        RECT 1229.680 144.880 1229.940 145.140 ;
        RECT 1229.680 110.540 1229.940 110.800 ;
        RECT 1228.760 110.200 1229.020 110.460 ;
        RECT 222.740 45.600 223.000 45.860 ;
        RECT 1228.760 45.600 1229.020 45.860 ;
      LAYER met2 ;
        RECT 1232.825 1700.410 1233.105 1704.000 ;
        RECT 1231.120 1700.270 1233.105 1700.410 ;
        RECT 1231.120 1635.730 1231.260 1700.270 ;
        RECT 1232.825 1700.000 1233.105 1700.270 ;
        RECT 1229.680 1635.410 1229.940 1635.730 ;
        RECT 1231.060 1635.410 1231.320 1635.730 ;
        RECT 1229.740 1352.510 1229.880 1635.410 ;
        RECT 1229.680 1352.190 1229.940 1352.510 ;
        RECT 1229.680 1304.250 1229.940 1304.570 ;
        RECT 1229.740 1255.950 1229.880 1304.250 ;
        RECT 1229.680 1255.630 1229.940 1255.950 ;
        RECT 1229.680 1207.350 1229.940 1207.670 ;
        RECT 1229.740 1159.245 1229.880 1207.350 ;
        RECT 1228.750 1158.875 1229.030 1159.245 ;
        RECT 1229.670 1158.875 1229.950 1159.245 ;
        RECT 1228.820 1111.110 1228.960 1158.875 ;
        RECT 1228.760 1110.790 1229.020 1111.110 ;
        RECT 1229.680 1110.790 1229.940 1111.110 ;
        RECT 1229.740 772.810 1229.880 1110.790 ;
        RECT 1228.760 772.490 1229.020 772.810 ;
        RECT 1229.680 772.490 1229.940 772.810 ;
        RECT 1228.820 724.725 1228.960 772.490 ;
        RECT 1228.750 724.355 1229.030 724.725 ;
        RECT 1229.670 724.355 1229.950 724.725 ;
        RECT 1229.740 676.250 1229.880 724.355 ;
        RECT 1228.760 675.930 1229.020 676.250 ;
        RECT 1229.680 675.930 1229.940 676.250 ;
        RECT 1228.820 628.165 1228.960 675.930 ;
        RECT 1228.750 627.795 1229.030 628.165 ;
        RECT 1229.670 627.795 1229.950 628.165 ;
        RECT 1229.740 579.690 1229.880 627.795 ;
        RECT 1229.680 579.370 1229.940 579.690 ;
        RECT 1229.680 531.430 1229.940 531.750 ;
        RECT 1229.740 289.670 1229.880 531.430 ;
        RECT 1229.680 289.350 1229.940 289.670 ;
        RECT 1229.680 241.410 1229.940 241.730 ;
        RECT 1229.740 193.110 1229.880 241.410 ;
        RECT 1229.680 192.790 1229.940 193.110 ;
        RECT 1229.680 144.850 1229.940 145.170 ;
        RECT 1229.740 110.830 1229.880 144.850 ;
        RECT 1229.680 110.510 1229.940 110.830 ;
        RECT 1228.760 110.170 1229.020 110.490 ;
        RECT 1228.820 45.890 1228.960 110.170 ;
        RECT 222.740 45.570 223.000 45.890 ;
        RECT 1228.760 45.570 1229.020 45.890 ;
        RECT 222.800 2.400 222.940 45.570 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 1228.750 1158.920 1229.030 1159.200 ;
        RECT 1229.670 1158.920 1229.950 1159.200 ;
        RECT 1228.750 724.400 1229.030 724.680 ;
        RECT 1229.670 724.400 1229.950 724.680 ;
        RECT 1228.750 627.840 1229.030 628.120 ;
        RECT 1229.670 627.840 1229.950 628.120 ;
      LAYER met3 ;
        RECT 1228.725 1159.210 1229.055 1159.225 ;
        RECT 1229.645 1159.210 1229.975 1159.225 ;
        RECT 1228.725 1158.910 1229.975 1159.210 ;
        RECT 1228.725 1158.895 1229.055 1158.910 ;
        RECT 1229.645 1158.895 1229.975 1158.910 ;
        RECT 1228.725 724.690 1229.055 724.705 ;
        RECT 1229.645 724.690 1229.975 724.705 ;
        RECT 1228.725 724.390 1229.975 724.690 ;
        RECT 1228.725 724.375 1229.055 724.390 ;
        RECT 1229.645 724.375 1229.975 724.390 ;
        RECT 1228.725 628.130 1229.055 628.145 ;
        RECT 1229.645 628.130 1229.975 628.145 ;
        RECT 1228.725 627.830 1229.975 628.130 ;
        RECT 1228.725 627.815 1229.055 627.830 ;
        RECT 1229.645 627.815 1229.975 627.830 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.465 1700.410 1156.745 1704.000 ;
        RECT 1155.220 1700.270 1156.745 1700.410 ;
        RECT 1155.220 1678.650 1155.360 1700.270 ;
        RECT 1156.465 1700.000 1156.745 1700.270 ;
        RECT 1152.920 1678.510 1155.360 1678.650 ;
        RECT 1152.920 37.925 1153.060 1678.510 ;
        RECT 19.870 37.555 20.150 37.925 ;
        RECT 1152.850 37.555 1153.130 37.925 ;
        RECT 19.940 3.130 20.080 37.555 ;
        RECT 19.940 2.990 20.540 3.130 ;
        RECT 20.400 2.400 20.540 2.990 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 19.870 37.600 20.150 37.880 ;
        RECT 1152.850 37.600 1153.130 37.880 ;
      LAYER met3 ;
        RECT 19.845 37.890 20.175 37.905 ;
        RECT 1152.825 37.890 1153.155 37.905 ;
        RECT 19.845 37.590 1153.155 37.890 ;
        RECT 19.845 37.575 20.175 37.590 ;
        RECT 1152.825 37.575 1153.155 37.590 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1138.185 34.425 1138.355 37.995 ;
      LAYER mcon ;
        RECT 1138.185 37.825 1138.355 37.995 ;
      LAYER met1 ;
        RECT 1160.190 1678.480 1160.510 1678.540 ;
        RECT 1163.870 1678.480 1164.190 1678.540 ;
        RECT 1160.190 1678.340 1164.190 1678.480 ;
        RECT 1160.190 1678.280 1160.510 1678.340 ;
        RECT 1163.870 1678.280 1164.190 1678.340 ;
        RECT 44.230 37.980 44.550 38.040 ;
        RECT 1138.125 37.980 1138.415 38.025 ;
        RECT 44.230 37.840 1138.415 37.980 ;
        RECT 44.230 37.780 44.550 37.840 ;
        RECT 1138.125 37.795 1138.415 37.840 ;
        RECT 1138.125 34.580 1138.415 34.625 ;
        RECT 1160.190 34.580 1160.510 34.640 ;
        RECT 1138.125 34.440 1160.510 34.580 ;
        RECT 1138.125 34.395 1138.415 34.440 ;
        RECT 1160.190 34.380 1160.510 34.440 ;
      LAYER via ;
        RECT 1160.220 1678.280 1160.480 1678.540 ;
        RECT 1163.900 1678.280 1164.160 1678.540 ;
        RECT 44.260 37.780 44.520 38.040 ;
        RECT 1160.220 34.380 1160.480 34.640 ;
      LAYER met2 ;
        RECT 1165.665 1700.410 1165.945 1704.000 ;
        RECT 1163.960 1700.270 1165.945 1700.410 ;
        RECT 1163.960 1678.570 1164.100 1700.270 ;
        RECT 1165.665 1700.000 1165.945 1700.270 ;
        RECT 1160.220 1678.250 1160.480 1678.570 ;
        RECT 1163.900 1678.250 1164.160 1678.570 ;
        RECT 44.260 37.750 44.520 38.070 ;
        RECT 44.320 2.400 44.460 37.750 ;
        RECT 1160.280 34.670 1160.420 1678.250 ;
        RECT 1160.220 34.350 1160.480 34.670 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 51.580 246.950 51.640 ;
        RECT 1242.530 51.580 1242.850 51.640 ;
        RECT 246.630 51.440 1242.850 51.580 ;
        RECT 246.630 51.380 246.950 51.440 ;
        RECT 1242.530 51.380 1242.850 51.440 ;
      LAYER via ;
        RECT 246.660 51.380 246.920 51.640 ;
        RECT 1242.560 51.380 1242.820 51.640 ;
      LAYER met2 ;
        RECT 1242.025 1700.410 1242.305 1704.000 ;
        RECT 1242.025 1700.270 1242.760 1700.410 ;
        RECT 1242.025 1700.000 1242.305 1700.270 ;
        RECT 1242.620 51.670 1242.760 1700.270 ;
        RECT 246.660 51.350 246.920 51.670 ;
        RECT 1242.560 51.350 1242.820 51.670 ;
        RECT 246.720 2.400 246.860 51.350 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.990 1662.160 1243.310 1662.220 ;
        RECT 1246.670 1662.160 1246.990 1662.220 ;
        RECT 1242.990 1662.020 1246.990 1662.160 ;
        RECT 1242.990 1661.960 1243.310 1662.020 ;
        RECT 1246.670 1661.960 1246.990 1662.020 ;
        RECT 264.110 51.920 264.430 51.980 ;
        RECT 1242.990 51.920 1243.310 51.980 ;
        RECT 264.110 51.780 1243.310 51.920 ;
        RECT 264.110 51.720 264.430 51.780 ;
        RECT 1242.990 51.720 1243.310 51.780 ;
      LAYER via ;
        RECT 1243.020 1661.960 1243.280 1662.220 ;
        RECT 1246.700 1661.960 1246.960 1662.220 ;
        RECT 264.140 51.720 264.400 51.980 ;
        RECT 1243.020 51.720 1243.280 51.980 ;
      LAYER met2 ;
        RECT 1248.465 1700.410 1248.745 1704.000 ;
        RECT 1246.760 1700.270 1248.745 1700.410 ;
        RECT 1246.760 1662.250 1246.900 1700.270 ;
        RECT 1248.465 1700.000 1248.745 1700.270 ;
        RECT 1243.020 1661.930 1243.280 1662.250 ;
        RECT 1246.700 1661.930 1246.960 1662.250 ;
        RECT 1243.080 52.010 1243.220 1661.930 ;
        RECT 264.140 51.690 264.400 52.010 ;
        RECT 1243.020 51.690 1243.280 52.010 ;
        RECT 264.200 2.400 264.340 51.690 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1249.430 1678.140 1249.750 1678.200 ;
        RECT 1254.030 1678.140 1254.350 1678.200 ;
        RECT 1249.430 1678.000 1254.350 1678.140 ;
        RECT 1249.430 1677.940 1249.750 1678.000 ;
        RECT 1254.030 1677.940 1254.350 1678.000 ;
        RECT 282.050 52.260 282.370 52.320 ;
        RECT 1249.430 52.260 1249.750 52.320 ;
        RECT 282.050 52.120 1249.750 52.260 ;
        RECT 282.050 52.060 282.370 52.120 ;
        RECT 1249.430 52.060 1249.750 52.120 ;
      LAYER via ;
        RECT 1249.460 1677.940 1249.720 1678.200 ;
        RECT 1254.060 1677.940 1254.320 1678.200 ;
        RECT 282.080 52.060 282.340 52.320 ;
        RECT 1249.460 52.060 1249.720 52.320 ;
      LAYER met2 ;
        RECT 1255.365 1700.410 1255.645 1704.000 ;
        RECT 1254.120 1700.270 1255.645 1700.410 ;
        RECT 1254.120 1678.230 1254.260 1700.270 ;
        RECT 1255.365 1700.000 1255.645 1700.270 ;
        RECT 1249.460 1677.910 1249.720 1678.230 ;
        RECT 1254.060 1677.910 1254.320 1678.230 ;
        RECT 1249.520 52.350 1249.660 1677.910 ;
        RECT 282.080 52.030 282.340 52.350 ;
        RECT 1249.460 52.030 1249.720 52.350 ;
        RECT 282.140 2.400 282.280 52.030 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1256.330 1678.140 1256.650 1678.200 ;
        RECT 1260.470 1678.140 1260.790 1678.200 ;
        RECT 1256.330 1678.000 1260.790 1678.140 ;
        RECT 1256.330 1677.940 1256.650 1678.000 ;
        RECT 1260.470 1677.940 1260.790 1678.000 ;
        RECT 299.990 52.600 300.310 52.660 ;
        RECT 1256.330 52.600 1256.650 52.660 ;
        RECT 299.990 52.460 1256.650 52.600 ;
        RECT 299.990 52.400 300.310 52.460 ;
        RECT 1256.330 52.400 1256.650 52.460 ;
      LAYER via ;
        RECT 1256.360 1677.940 1256.620 1678.200 ;
        RECT 1260.500 1677.940 1260.760 1678.200 ;
        RECT 300.020 52.400 300.280 52.660 ;
        RECT 1256.360 52.400 1256.620 52.660 ;
      LAYER met2 ;
        RECT 1261.805 1700.410 1262.085 1704.000 ;
        RECT 1260.560 1700.270 1262.085 1700.410 ;
        RECT 1260.560 1678.230 1260.700 1700.270 ;
        RECT 1261.805 1700.000 1262.085 1700.270 ;
        RECT 1256.360 1677.910 1256.620 1678.230 ;
        RECT 1260.500 1677.910 1260.760 1678.230 ;
        RECT 1256.420 52.690 1256.560 1677.910 ;
        RECT 300.020 52.370 300.280 52.690 ;
        RECT 1256.360 52.370 1256.620 52.690 ;
        RECT 300.080 2.400 300.220 52.370 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1263.230 1678.140 1263.550 1678.200 ;
        RECT 1266.910 1678.140 1267.230 1678.200 ;
        RECT 1263.230 1678.000 1267.230 1678.140 ;
        RECT 1263.230 1677.940 1263.550 1678.000 ;
        RECT 1266.910 1677.940 1267.230 1678.000 ;
        RECT 317.930 52.940 318.250 53.000 ;
        RECT 1263.230 52.940 1263.550 53.000 ;
        RECT 317.930 52.800 1263.550 52.940 ;
        RECT 317.930 52.740 318.250 52.800 ;
        RECT 1263.230 52.740 1263.550 52.800 ;
      LAYER via ;
        RECT 1263.260 1677.940 1263.520 1678.200 ;
        RECT 1266.940 1677.940 1267.200 1678.200 ;
        RECT 317.960 52.740 318.220 53.000 ;
        RECT 1263.260 52.740 1263.520 53.000 ;
      LAYER met2 ;
        RECT 1268.705 1700.410 1268.985 1704.000 ;
        RECT 1267.000 1700.270 1268.985 1700.410 ;
        RECT 1267.000 1678.230 1267.140 1700.270 ;
        RECT 1268.705 1700.000 1268.985 1700.270 ;
        RECT 1263.260 1677.910 1263.520 1678.230 ;
        RECT 1266.940 1677.910 1267.200 1678.230 ;
        RECT 1263.320 53.030 1263.460 1677.910 ;
        RECT 317.960 52.710 318.220 53.030 ;
        RECT 1263.260 52.710 1263.520 53.030 ;
        RECT 318.020 2.400 318.160 52.710 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1271.125 1352.605 1271.295 1400.715 ;
        RECT 1271.125 1256.045 1271.295 1304.155 ;
        RECT 1271.125 579.785 1271.295 627.895 ;
        RECT 1270.665 234.685 1270.835 282.795 ;
        RECT 1270.665 48.365 1270.835 113.815 ;
      LAYER mcon ;
        RECT 1271.125 1400.545 1271.295 1400.715 ;
        RECT 1271.125 1303.985 1271.295 1304.155 ;
        RECT 1271.125 627.725 1271.295 627.895 ;
        RECT 1270.665 282.625 1270.835 282.795 ;
        RECT 1270.665 113.645 1270.835 113.815 ;
      LAYER met1 ;
        RECT 1271.050 1642.100 1271.370 1642.160 ;
        RECT 1271.510 1642.100 1271.830 1642.160 ;
        RECT 1271.050 1641.960 1271.830 1642.100 ;
        RECT 1271.050 1641.900 1271.370 1641.960 ;
        RECT 1271.510 1641.900 1271.830 1641.960 ;
        RECT 1270.590 1532.280 1270.910 1532.340 ;
        RECT 1271.510 1532.280 1271.830 1532.340 ;
        RECT 1270.590 1532.140 1271.830 1532.280 ;
        RECT 1270.590 1532.080 1270.910 1532.140 ;
        RECT 1271.510 1532.080 1271.830 1532.140 ;
        RECT 1269.670 1483.660 1269.990 1483.720 ;
        RECT 1271.050 1483.660 1271.370 1483.720 ;
        RECT 1269.670 1483.520 1271.370 1483.660 ;
        RECT 1269.670 1483.460 1269.990 1483.520 ;
        RECT 1271.050 1483.460 1271.370 1483.520 ;
        RECT 1271.050 1463.060 1271.370 1463.320 ;
        RECT 1271.140 1462.640 1271.280 1463.060 ;
        RECT 1271.050 1462.380 1271.370 1462.640 ;
        RECT 1271.050 1400.700 1271.370 1400.760 ;
        RECT 1270.855 1400.560 1271.370 1400.700 ;
        RECT 1271.050 1400.500 1271.370 1400.560 ;
        RECT 1271.050 1352.760 1271.370 1352.820 ;
        RECT 1270.855 1352.620 1271.370 1352.760 ;
        RECT 1271.050 1352.560 1271.370 1352.620 ;
        RECT 1271.050 1304.140 1271.370 1304.200 ;
        RECT 1270.855 1304.000 1271.370 1304.140 ;
        RECT 1271.050 1303.940 1271.370 1304.000 ;
        RECT 1271.050 1256.200 1271.370 1256.260 ;
        RECT 1270.855 1256.060 1271.370 1256.200 ;
        RECT 1271.050 1256.000 1271.370 1256.060 ;
        RECT 1271.050 1159.300 1271.370 1159.360 ;
        RECT 1271.970 1159.300 1272.290 1159.360 ;
        RECT 1271.050 1159.160 1272.290 1159.300 ;
        RECT 1271.050 1159.100 1271.370 1159.160 ;
        RECT 1271.970 1159.100 1272.290 1159.160 ;
        RECT 1271.050 1062.740 1271.370 1062.800 ;
        RECT 1271.970 1062.740 1272.290 1062.800 ;
        RECT 1271.050 1062.600 1272.290 1062.740 ;
        RECT 1271.050 1062.540 1271.370 1062.600 ;
        RECT 1271.970 1062.540 1272.290 1062.600 ;
        RECT 1271.050 983.180 1271.370 983.240 ;
        RECT 1271.970 983.180 1272.290 983.240 ;
        RECT 1271.050 983.040 1272.290 983.180 ;
        RECT 1271.050 982.980 1271.370 983.040 ;
        RECT 1271.970 982.980 1272.290 983.040 ;
        RECT 1271.050 821.000 1271.370 821.060 ;
        RECT 1271.970 821.000 1272.290 821.060 ;
        RECT 1271.050 820.860 1272.290 821.000 ;
        RECT 1271.050 820.800 1271.370 820.860 ;
        RECT 1271.970 820.800 1272.290 820.860 ;
        RECT 1271.050 724.440 1271.370 724.500 ;
        RECT 1271.970 724.440 1272.290 724.500 ;
        RECT 1271.050 724.300 1272.290 724.440 ;
        RECT 1271.050 724.240 1271.370 724.300 ;
        RECT 1271.970 724.240 1272.290 724.300 ;
        RECT 1271.050 627.880 1271.370 627.940 ;
        RECT 1270.855 627.740 1271.370 627.880 ;
        RECT 1271.050 627.680 1271.370 627.740 ;
        RECT 1271.050 579.940 1271.370 580.000 ;
        RECT 1270.855 579.800 1271.370 579.940 ;
        RECT 1271.050 579.740 1271.370 579.800 ;
        RECT 1271.050 400.220 1271.370 400.480 ;
        RECT 1271.140 399.800 1271.280 400.220 ;
        RECT 1271.050 399.540 1271.370 399.800 ;
        RECT 1270.590 282.780 1270.910 282.840 ;
        RECT 1270.395 282.640 1270.910 282.780 ;
        RECT 1270.590 282.580 1270.910 282.640 ;
        RECT 1270.590 234.840 1270.910 234.900 ;
        RECT 1270.395 234.700 1270.910 234.840 ;
        RECT 1270.590 234.640 1270.910 234.700 ;
        RECT 1270.590 186.560 1270.910 186.620 ;
        RECT 1271.050 186.560 1271.370 186.620 ;
        RECT 1270.590 186.420 1271.370 186.560 ;
        RECT 1270.590 186.360 1270.910 186.420 ;
        RECT 1271.050 186.360 1271.370 186.420 ;
        RECT 1269.670 162.080 1269.990 162.140 ;
        RECT 1271.050 162.080 1271.370 162.140 ;
        RECT 1269.670 161.940 1271.370 162.080 ;
        RECT 1269.670 161.880 1269.990 161.940 ;
        RECT 1271.050 161.880 1271.370 161.940 ;
        RECT 1269.670 113.800 1269.990 113.860 ;
        RECT 1270.605 113.800 1270.895 113.845 ;
        RECT 1269.670 113.660 1270.895 113.800 ;
        RECT 1269.670 113.600 1269.990 113.660 ;
        RECT 1270.605 113.615 1270.895 113.660 ;
        RECT 1270.590 48.520 1270.910 48.580 ;
        RECT 1270.395 48.380 1270.910 48.520 ;
        RECT 1270.590 48.320 1270.910 48.380 ;
        RECT 335.870 26.420 336.190 26.480 ;
        RECT 1270.590 26.420 1270.910 26.480 ;
        RECT 335.870 26.280 1270.910 26.420 ;
        RECT 335.870 26.220 336.190 26.280 ;
        RECT 1270.590 26.220 1270.910 26.280 ;
      LAYER via ;
        RECT 1271.080 1641.900 1271.340 1642.160 ;
        RECT 1271.540 1641.900 1271.800 1642.160 ;
        RECT 1270.620 1532.080 1270.880 1532.340 ;
        RECT 1271.540 1532.080 1271.800 1532.340 ;
        RECT 1269.700 1483.460 1269.960 1483.720 ;
        RECT 1271.080 1483.460 1271.340 1483.720 ;
        RECT 1271.080 1463.060 1271.340 1463.320 ;
        RECT 1271.080 1462.380 1271.340 1462.640 ;
        RECT 1271.080 1400.500 1271.340 1400.760 ;
        RECT 1271.080 1352.560 1271.340 1352.820 ;
        RECT 1271.080 1303.940 1271.340 1304.200 ;
        RECT 1271.080 1256.000 1271.340 1256.260 ;
        RECT 1271.080 1159.100 1271.340 1159.360 ;
        RECT 1272.000 1159.100 1272.260 1159.360 ;
        RECT 1271.080 1062.540 1271.340 1062.800 ;
        RECT 1272.000 1062.540 1272.260 1062.800 ;
        RECT 1271.080 982.980 1271.340 983.240 ;
        RECT 1272.000 982.980 1272.260 983.240 ;
        RECT 1271.080 820.800 1271.340 821.060 ;
        RECT 1272.000 820.800 1272.260 821.060 ;
        RECT 1271.080 724.240 1271.340 724.500 ;
        RECT 1272.000 724.240 1272.260 724.500 ;
        RECT 1271.080 627.680 1271.340 627.940 ;
        RECT 1271.080 579.740 1271.340 580.000 ;
        RECT 1271.080 400.220 1271.340 400.480 ;
        RECT 1271.080 399.540 1271.340 399.800 ;
        RECT 1270.620 282.580 1270.880 282.840 ;
        RECT 1270.620 234.640 1270.880 234.900 ;
        RECT 1270.620 186.360 1270.880 186.620 ;
        RECT 1271.080 186.360 1271.340 186.620 ;
        RECT 1269.700 161.880 1269.960 162.140 ;
        RECT 1271.080 161.880 1271.340 162.140 ;
        RECT 1269.700 113.600 1269.960 113.860 ;
        RECT 1270.620 48.320 1270.880 48.580 ;
        RECT 335.900 26.220 336.160 26.480 ;
        RECT 1270.620 26.220 1270.880 26.480 ;
      LAYER met2 ;
        RECT 1275.605 1700.410 1275.885 1704.000 ;
        RECT 1273.900 1700.270 1275.885 1700.410 ;
        RECT 1273.900 1690.210 1274.040 1700.270 ;
        RECT 1275.605 1700.000 1275.885 1700.270 ;
        RECT 1272.060 1690.070 1274.040 1690.210 ;
        RECT 1272.060 1677.290 1272.200 1690.070 ;
        RECT 1271.140 1677.150 1272.200 1677.290 ;
        RECT 1271.140 1642.190 1271.280 1677.150 ;
        RECT 1271.080 1641.870 1271.340 1642.190 ;
        RECT 1271.540 1641.870 1271.800 1642.190 ;
        RECT 1271.600 1611.330 1271.740 1641.870 ;
        RECT 1270.680 1611.190 1271.740 1611.330 ;
        RECT 1270.680 1580.050 1270.820 1611.190 ;
        RECT 1270.680 1579.910 1271.740 1580.050 ;
        RECT 1271.600 1532.370 1271.740 1579.910 ;
        RECT 1270.620 1532.050 1270.880 1532.370 ;
        RECT 1271.540 1532.050 1271.800 1532.370 ;
        RECT 1270.680 1531.885 1270.820 1532.050 ;
        RECT 1269.690 1531.515 1269.970 1531.885 ;
        RECT 1270.610 1531.515 1270.890 1531.885 ;
        RECT 1269.760 1483.750 1269.900 1531.515 ;
        RECT 1269.700 1483.430 1269.960 1483.750 ;
        RECT 1271.080 1483.430 1271.340 1483.750 ;
        RECT 1271.140 1463.350 1271.280 1483.430 ;
        RECT 1271.080 1463.030 1271.340 1463.350 ;
        RECT 1271.080 1462.350 1271.340 1462.670 ;
        RECT 1271.140 1400.790 1271.280 1462.350 ;
        RECT 1271.080 1400.470 1271.340 1400.790 ;
        RECT 1271.080 1352.530 1271.340 1352.850 ;
        RECT 1271.140 1304.230 1271.280 1352.530 ;
        RECT 1271.080 1303.910 1271.340 1304.230 ;
        RECT 1271.080 1255.970 1271.340 1256.290 ;
        RECT 1271.140 1207.525 1271.280 1255.970 ;
        RECT 1271.070 1207.155 1271.350 1207.525 ;
        RECT 1271.990 1207.155 1272.270 1207.525 ;
        RECT 1272.060 1159.390 1272.200 1207.155 ;
        RECT 1271.080 1159.070 1271.340 1159.390 ;
        RECT 1272.000 1159.070 1272.260 1159.390 ;
        RECT 1271.140 1110.965 1271.280 1159.070 ;
        RECT 1271.070 1110.595 1271.350 1110.965 ;
        RECT 1271.990 1110.595 1272.270 1110.965 ;
        RECT 1272.060 1062.830 1272.200 1110.595 ;
        RECT 1271.080 1062.510 1271.340 1062.830 ;
        RECT 1272.000 1062.510 1272.260 1062.830 ;
        RECT 1271.140 983.270 1271.280 1062.510 ;
        RECT 1271.080 982.950 1271.340 983.270 ;
        RECT 1272.000 982.950 1272.260 983.270 ;
        RECT 1272.060 959.325 1272.200 982.950 ;
        RECT 1271.070 958.955 1271.350 959.325 ;
        RECT 1271.990 958.955 1272.270 959.325 ;
        RECT 1271.140 821.090 1271.280 958.955 ;
        RECT 1271.080 820.770 1271.340 821.090 ;
        RECT 1272.000 820.770 1272.260 821.090 ;
        RECT 1272.060 773.005 1272.200 820.770 ;
        RECT 1271.070 772.635 1271.350 773.005 ;
        RECT 1271.990 772.635 1272.270 773.005 ;
        RECT 1271.140 724.530 1271.280 772.635 ;
        RECT 1271.080 724.210 1271.340 724.530 ;
        RECT 1272.000 724.210 1272.260 724.530 ;
        RECT 1272.060 676.445 1272.200 724.210 ;
        RECT 1271.070 676.075 1271.350 676.445 ;
        RECT 1271.990 676.075 1272.270 676.445 ;
        RECT 1271.140 627.970 1271.280 676.075 ;
        RECT 1271.080 627.650 1271.340 627.970 ;
        RECT 1271.080 579.710 1271.340 580.030 ;
        RECT 1271.140 497.490 1271.280 579.710 ;
        RECT 1270.680 497.350 1271.280 497.490 ;
        RECT 1270.680 496.810 1270.820 497.350 ;
        RECT 1270.680 496.670 1271.280 496.810 ;
        RECT 1271.140 400.510 1271.280 496.670 ;
        RECT 1271.080 400.190 1271.340 400.510 ;
        RECT 1271.080 399.510 1271.340 399.830 ;
        RECT 1271.140 283.290 1271.280 399.510 ;
        RECT 1270.680 283.150 1271.280 283.290 ;
        RECT 1270.680 282.870 1270.820 283.150 ;
        RECT 1270.620 282.550 1270.880 282.870 ;
        RECT 1270.620 234.610 1270.880 234.930 ;
        RECT 1270.680 186.650 1270.820 234.610 ;
        RECT 1270.620 186.330 1270.880 186.650 ;
        RECT 1271.080 186.330 1271.340 186.650 ;
        RECT 1271.140 162.170 1271.280 186.330 ;
        RECT 1269.700 161.850 1269.960 162.170 ;
        RECT 1271.080 161.850 1271.340 162.170 ;
        RECT 1269.760 113.890 1269.900 161.850 ;
        RECT 1269.700 113.570 1269.960 113.890 ;
        RECT 1270.620 48.290 1270.880 48.610 ;
        RECT 1270.680 26.510 1270.820 48.290 ;
        RECT 335.900 26.190 336.160 26.510 ;
        RECT 1270.620 26.190 1270.880 26.510 ;
        RECT 335.960 2.400 336.100 26.190 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1269.690 1531.560 1269.970 1531.840 ;
        RECT 1270.610 1531.560 1270.890 1531.840 ;
        RECT 1271.070 1207.200 1271.350 1207.480 ;
        RECT 1271.990 1207.200 1272.270 1207.480 ;
        RECT 1271.070 1110.640 1271.350 1110.920 ;
        RECT 1271.990 1110.640 1272.270 1110.920 ;
        RECT 1271.070 959.000 1271.350 959.280 ;
        RECT 1271.990 959.000 1272.270 959.280 ;
        RECT 1271.070 772.680 1271.350 772.960 ;
        RECT 1271.990 772.680 1272.270 772.960 ;
        RECT 1271.070 676.120 1271.350 676.400 ;
        RECT 1271.990 676.120 1272.270 676.400 ;
      LAYER met3 ;
        RECT 1269.665 1531.850 1269.995 1531.865 ;
        RECT 1270.585 1531.850 1270.915 1531.865 ;
        RECT 1269.665 1531.550 1270.915 1531.850 ;
        RECT 1269.665 1531.535 1269.995 1531.550 ;
        RECT 1270.585 1531.535 1270.915 1531.550 ;
        RECT 1271.045 1207.490 1271.375 1207.505 ;
        RECT 1271.965 1207.490 1272.295 1207.505 ;
        RECT 1271.045 1207.190 1272.295 1207.490 ;
        RECT 1271.045 1207.175 1271.375 1207.190 ;
        RECT 1271.965 1207.175 1272.295 1207.190 ;
        RECT 1271.045 1110.930 1271.375 1110.945 ;
        RECT 1271.965 1110.930 1272.295 1110.945 ;
        RECT 1271.045 1110.630 1272.295 1110.930 ;
        RECT 1271.045 1110.615 1271.375 1110.630 ;
        RECT 1271.965 1110.615 1272.295 1110.630 ;
        RECT 1271.045 959.290 1271.375 959.305 ;
        RECT 1271.965 959.290 1272.295 959.305 ;
        RECT 1271.045 958.990 1272.295 959.290 ;
        RECT 1271.045 958.975 1271.375 958.990 ;
        RECT 1271.965 958.975 1272.295 958.990 ;
        RECT 1271.045 772.970 1271.375 772.985 ;
        RECT 1271.965 772.970 1272.295 772.985 ;
        RECT 1271.045 772.670 1272.295 772.970 ;
        RECT 1271.045 772.655 1271.375 772.670 ;
        RECT 1271.965 772.655 1272.295 772.670 ;
        RECT 1271.045 676.410 1271.375 676.425 ;
        RECT 1271.965 676.410 1272.295 676.425 ;
        RECT 1271.045 676.110 1272.295 676.410 ;
        RECT 1271.045 676.095 1271.375 676.110 ;
        RECT 1271.965 676.095 1272.295 676.110 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1277.030 1678.140 1277.350 1678.200 ;
        RECT 1280.710 1678.140 1281.030 1678.200 ;
        RECT 1277.030 1678.000 1281.030 1678.140 ;
        RECT 1277.030 1677.940 1277.350 1678.000 ;
        RECT 1280.710 1677.940 1281.030 1678.000 ;
        RECT 358.410 65.860 358.730 65.920 ;
        RECT 1277.030 65.860 1277.350 65.920 ;
        RECT 358.410 65.720 1277.350 65.860 ;
        RECT 358.410 65.660 358.730 65.720 ;
        RECT 1277.030 65.660 1277.350 65.720 ;
        RECT 353.350 16.560 353.670 16.620 ;
        RECT 358.410 16.560 358.730 16.620 ;
        RECT 353.350 16.420 358.730 16.560 ;
        RECT 353.350 16.360 353.670 16.420 ;
        RECT 358.410 16.360 358.730 16.420 ;
      LAYER via ;
        RECT 1277.060 1677.940 1277.320 1678.200 ;
        RECT 1280.740 1677.940 1281.000 1678.200 ;
        RECT 358.440 65.660 358.700 65.920 ;
        RECT 1277.060 65.660 1277.320 65.920 ;
        RECT 353.380 16.360 353.640 16.620 ;
        RECT 358.440 16.360 358.700 16.620 ;
      LAYER met2 ;
        RECT 1282.045 1700.410 1282.325 1704.000 ;
        RECT 1280.800 1700.270 1282.325 1700.410 ;
        RECT 1280.800 1678.230 1280.940 1700.270 ;
        RECT 1282.045 1700.000 1282.325 1700.270 ;
        RECT 1277.060 1677.910 1277.320 1678.230 ;
        RECT 1280.740 1677.910 1281.000 1678.230 ;
        RECT 1277.120 65.950 1277.260 1677.910 ;
        RECT 358.440 65.630 358.700 65.950 ;
        RECT 1277.060 65.630 1277.320 65.950 ;
        RECT 358.500 16.650 358.640 65.630 ;
        RECT 353.380 16.330 353.640 16.650 ;
        RECT 358.440 16.330 358.700 16.650 ;
        RECT 353.440 2.400 353.580 16.330 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.930 1670.320 1284.250 1670.380 ;
        RECT 1287.150 1670.320 1287.470 1670.380 ;
        RECT 1283.930 1670.180 1287.470 1670.320 ;
        RECT 1283.930 1670.120 1284.250 1670.180 ;
        RECT 1287.150 1670.120 1287.470 1670.180 ;
        RECT 372.210 72.660 372.530 72.720 ;
        RECT 1283.930 72.660 1284.250 72.720 ;
        RECT 372.210 72.520 1284.250 72.660 ;
        RECT 372.210 72.460 372.530 72.520 ;
        RECT 1283.930 72.460 1284.250 72.520 ;
      LAYER via ;
        RECT 1283.960 1670.120 1284.220 1670.380 ;
        RECT 1287.180 1670.120 1287.440 1670.380 ;
        RECT 372.240 72.460 372.500 72.720 ;
        RECT 1283.960 72.460 1284.220 72.720 ;
      LAYER met2 ;
        RECT 1288.945 1700.410 1289.225 1704.000 ;
        RECT 1287.240 1700.270 1289.225 1700.410 ;
        RECT 1287.240 1670.410 1287.380 1700.270 ;
        RECT 1288.945 1700.000 1289.225 1700.270 ;
        RECT 1283.960 1670.090 1284.220 1670.410 ;
        RECT 1287.180 1670.090 1287.440 1670.410 ;
        RECT 1284.020 72.750 1284.160 1670.090 ;
        RECT 372.240 72.430 372.500 72.750 ;
        RECT 1283.960 72.430 1284.220 72.750 ;
        RECT 372.300 16.900 372.440 72.430 ;
        RECT 371.380 16.760 372.440 16.900 ;
        RECT 371.380 2.400 371.520 16.760 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1290.830 1678.140 1291.150 1678.200 ;
        RECT 1294.510 1678.140 1294.830 1678.200 ;
        RECT 1290.830 1678.000 1294.830 1678.140 ;
        RECT 1290.830 1677.940 1291.150 1678.000 ;
        RECT 1294.510 1677.940 1294.830 1678.000 ;
        RECT 392.910 73.000 393.230 73.060 ;
        RECT 1290.830 73.000 1291.150 73.060 ;
        RECT 392.910 72.860 1291.150 73.000 ;
        RECT 392.910 72.800 393.230 72.860 ;
        RECT 1290.830 72.800 1291.150 72.860 ;
        RECT 389.230 16.220 389.550 16.280 ;
        RECT 392.910 16.220 393.230 16.280 ;
        RECT 389.230 16.080 393.230 16.220 ;
        RECT 389.230 16.020 389.550 16.080 ;
        RECT 392.910 16.020 393.230 16.080 ;
      LAYER via ;
        RECT 1290.860 1677.940 1291.120 1678.200 ;
        RECT 1294.540 1677.940 1294.800 1678.200 ;
        RECT 392.940 72.800 393.200 73.060 ;
        RECT 1290.860 72.800 1291.120 73.060 ;
        RECT 389.260 16.020 389.520 16.280 ;
        RECT 392.940 16.020 393.200 16.280 ;
      LAYER met2 ;
        RECT 1295.845 1700.410 1296.125 1704.000 ;
        RECT 1294.600 1700.270 1296.125 1700.410 ;
        RECT 1294.600 1678.230 1294.740 1700.270 ;
        RECT 1295.845 1700.000 1296.125 1700.270 ;
        RECT 1290.860 1677.910 1291.120 1678.230 ;
        RECT 1294.540 1677.910 1294.800 1678.230 ;
        RECT 1290.920 73.090 1291.060 1677.910 ;
        RECT 392.940 72.770 393.200 73.090 ;
        RECT 1290.860 72.770 1291.120 73.090 ;
        RECT 393.000 16.310 393.140 72.770 ;
        RECT 389.260 15.990 389.520 16.310 ;
        RECT 392.940 15.990 393.200 16.310 ;
        RECT 389.320 2.400 389.460 15.990 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1297.730 1678.140 1298.050 1678.200 ;
        RECT 1300.950 1678.140 1301.270 1678.200 ;
        RECT 1297.730 1678.000 1301.270 1678.140 ;
        RECT 1297.730 1677.940 1298.050 1678.000 ;
        RECT 1300.950 1677.940 1301.270 1678.000 ;
        RECT 413.610 73.340 413.930 73.400 ;
        RECT 1297.730 73.340 1298.050 73.400 ;
        RECT 413.610 73.200 1298.050 73.340 ;
        RECT 413.610 73.140 413.930 73.200 ;
        RECT 1297.730 73.140 1298.050 73.200 ;
        RECT 407.170 16.220 407.490 16.280 ;
        RECT 413.610 16.220 413.930 16.280 ;
        RECT 407.170 16.080 413.930 16.220 ;
        RECT 407.170 16.020 407.490 16.080 ;
        RECT 413.610 16.020 413.930 16.080 ;
      LAYER via ;
        RECT 1297.760 1677.940 1298.020 1678.200 ;
        RECT 1300.980 1677.940 1301.240 1678.200 ;
        RECT 413.640 73.140 413.900 73.400 ;
        RECT 1297.760 73.140 1298.020 73.400 ;
        RECT 407.200 16.020 407.460 16.280 ;
        RECT 413.640 16.020 413.900 16.280 ;
      LAYER met2 ;
        RECT 1302.285 1700.410 1302.565 1704.000 ;
        RECT 1301.040 1700.270 1302.565 1700.410 ;
        RECT 1301.040 1678.230 1301.180 1700.270 ;
        RECT 1302.285 1700.000 1302.565 1700.270 ;
        RECT 1297.760 1677.910 1298.020 1678.230 ;
        RECT 1300.980 1677.910 1301.240 1678.230 ;
        RECT 1297.820 73.430 1297.960 1677.910 ;
        RECT 413.640 73.110 413.900 73.430 ;
        RECT 1297.760 73.110 1298.020 73.430 ;
        RECT 413.700 16.310 413.840 73.110 ;
        RECT 407.200 15.990 407.460 16.310 ;
        RECT 413.640 15.990 413.900 16.310 ;
        RECT 407.260 2.400 407.400 15.990 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1174.065 1587.205 1174.235 1635.315 ;
        RECT 1174.525 1490.645 1174.695 1538.755 ;
        RECT 1174.525 1152.345 1174.695 1200.455 ;
        RECT 1174.065 961.265 1174.235 1007.335 ;
        RECT 1174.525 704.225 1174.695 806.735 ;
        RECT 1174.065 672.945 1174.235 703.715 ;
        RECT 1174.065 460.105 1174.235 503.795 ;
        RECT 1174.525 503.625 1174.695 600.355 ;
        RECT 1174.065 372.725 1174.235 420.835 ;
        RECT 1174.065 276.165 1174.235 324.275 ;
        RECT 1174.065 179.605 1174.235 227.715 ;
        RECT 1174.065 44.625 1174.235 131.155 ;
      LAYER mcon ;
        RECT 1174.065 1635.145 1174.235 1635.315 ;
        RECT 1174.525 1538.585 1174.695 1538.755 ;
        RECT 1174.525 1200.285 1174.695 1200.455 ;
        RECT 1174.065 1007.165 1174.235 1007.335 ;
        RECT 1174.525 806.565 1174.695 806.735 ;
        RECT 1174.065 703.545 1174.235 703.715 ;
        RECT 1174.525 600.185 1174.695 600.355 ;
        RECT 1174.065 503.625 1174.235 503.795 ;
        RECT 1174.065 420.665 1174.235 420.835 ;
        RECT 1174.065 324.105 1174.235 324.275 ;
        RECT 1174.065 227.545 1174.235 227.715 ;
        RECT 1174.065 130.985 1174.235 131.155 ;
      LAYER met1 ;
        RECT 1173.990 1635.300 1174.310 1635.360 ;
        RECT 1173.795 1635.160 1174.310 1635.300 ;
        RECT 1173.990 1635.100 1174.310 1635.160 ;
        RECT 1174.005 1587.360 1174.295 1587.405 ;
        RECT 1174.450 1587.360 1174.770 1587.420 ;
        RECT 1174.005 1587.220 1174.770 1587.360 ;
        RECT 1174.005 1587.175 1174.295 1587.220 ;
        RECT 1174.450 1587.160 1174.770 1587.220 ;
        RECT 1174.450 1538.740 1174.770 1538.800 ;
        RECT 1174.255 1538.600 1174.770 1538.740 ;
        RECT 1174.450 1538.540 1174.770 1538.600 ;
        RECT 1174.450 1490.800 1174.770 1490.860 ;
        RECT 1174.255 1490.660 1174.770 1490.800 ;
        RECT 1174.450 1490.600 1174.770 1490.660 ;
        RECT 1173.070 1297.340 1173.390 1297.400 ;
        RECT 1174.450 1297.340 1174.770 1297.400 ;
        RECT 1173.070 1297.200 1174.770 1297.340 ;
        RECT 1173.070 1297.140 1173.390 1297.200 ;
        RECT 1174.450 1297.140 1174.770 1297.200 ;
        RECT 1174.450 1256.000 1174.770 1256.260 ;
        RECT 1174.540 1255.520 1174.680 1256.000 ;
        RECT 1174.910 1255.520 1175.230 1255.580 ;
        RECT 1174.540 1255.380 1175.230 1255.520 ;
        RECT 1174.910 1255.320 1175.230 1255.380 ;
        RECT 1174.450 1207.580 1174.770 1207.640 ;
        RECT 1174.910 1207.580 1175.230 1207.640 ;
        RECT 1174.450 1207.440 1175.230 1207.580 ;
        RECT 1174.450 1207.380 1174.770 1207.440 ;
        RECT 1174.910 1207.380 1175.230 1207.440 ;
        RECT 1174.450 1200.440 1174.770 1200.500 ;
        RECT 1174.255 1200.300 1174.770 1200.440 ;
        RECT 1174.450 1200.240 1174.770 1200.300 ;
        RECT 1174.450 1152.500 1174.770 1152.560 ;
        RECT 1174.255 1152.360 1174.770 1152.500 ;
        RECT 1174.450 1152.300 1174.770 1152.360 ;
        RECT 1173.990 1014.460 1174.310 1014.520 ;
        RECT 1174.450 1014.460 1174.770 1014.520 ;
        RECT 1173.990 1014.320 1174.770 1014.460 ;
        RECT 1173.990 1014.260 1174.310 1014.320 ;
        RECT 1174.450 1014.260 1174.770 1014.320 ;
        RECT 1173.990 1007.320 1174.310 1007.380 ;
        RECT 1173.795 1007.180 1174.310 1007.320 ;
        RECT 1173.990 1007.120 1174.310 1007.180 ;
        RECT 1173.990 961.420 1174.310 961.480 ;
        RECT 1173.795 961.280 1174.310 961.420 ;
        RECT 1173.990 961.220 1174.310 961.280 ;
        RECT 1173.990 869.620 1174.310 869.680 ;
        RECT 1174.450 869.620 1174.770 869.680 ;
        RECT 1173.990 869.480 1174.770 869.620 ;
        RECT 1173.990 869.420 1174.310 869.480 ;
        RECT 1174.450 869.420 1174.770 869.480 ;
        RECT 1174.450 806.720 1174.770 806.780 ;
        RECT 1174.255 806.580 1174.770 806.720 ;
        RECT 1174.450 806.520 1174.770 806.580 ;
        RECT 1173.990 704.380 1174.310 704.440 ;
        RECT 1174.465 704.380 1174.755 704.425 ;
        RECT 1173.990 704.240 1174.755 704.380 ;
        RECT 1173.990 704.180 1174.310 704.240 ;
        RECT 1174.465 704.195 1174.755 704.240 ;
        RECT 1173.990 703.700 1174.310 703.760 ;
        RECT 1173.795 703.560 1174.310 703.700 ;
        RECT 1173.990 703.500 1174.310 703.560 ;
        RECT 1174.005 673.100 1174.295 673.145 ;
        RECT 1174.910 673.100 1175.230 673.160 ;
        RECT 1174.005 672.960 1175.230 673.100 ;
        RECT 1174.005 672.915 1174.295 672.960 ;
        RECT 1174.910 672.900 1175.230 672.960 ;
        RECT 1174.450 600.340 1174.770 600.400 ;
        RECT 1174.255 600.200 1174.770 600.340 ;
        RECT 1174.450 600.140 1174.770 600.200 ;
        RECT 1174.005 503.780 1174.295 503.825 ;
        RECT 1174.465 503.780 1174.755 503.825 ;
        RECT 1174.005 503.640 1174.755 503.780 ;
        RECT 1174.005 503.595 1174.295 503.640 ;
        RECT 1174.465 503.595 1174.755 503.640 ;
        RECT 1173.990 460.260 1174.310 460.320 ;
        RECT 1173.795 460.120 1174.310 460.260 ;
        RECT 1173.990 460.060 1174.310 460.120 ;
        RECT 1173.990 420.820 1174.310 420.880 ;
        RECT 1173.795 420.680 1174.310 420.820 ;
        RECT 1173.990 420.620 1174.310 420.680 ;
        RECT 1173.990 372.880 1174.310 372.940 ;
        RECT 1173.795 372.740 1174.310 372.880 ;
        RECT 1173.990 372.680 1174.310 372.740 ;
        RECT 1173.990 324.260 1174.310 324.320 ;
        RECT 1173.795 324.120 1174.310 324.260 ;
        RECT 1173.990 324.060 1174.310 324.120 ;
        RECT 1173.990 276.320 1174.310 276.380 ;
        RECT 1173.795 276.180 1174.310 276.320 ;
        RECT 1173.990 276.120 1174.310 276.180 ;
        RECT 1173.990 227.700 1174.310 227.760 ;
        RECT 1173.795 227.560 1174.310 227.700 ;
        RECT 1173.990 227.500 1174.310 227.560 ;
        RECT 1173.990 179.760 1174.310 179.820 ;
        RECT 1173.795 179.620 1174.310 179.760 ;
        RECT 1173.990 179.560 1174.310 179.620 ;
        RECT 1173.990 131.140 1174.310 131.200 ;
        RECT 1173.795 131.000 1174.310 131.140 ;
        RECT 1173.990 130.940 1174.310 131.000 ;
        RECT 68.150 44.780 68.470 44.840 ;
        RECT 1174.005 44.780 1174.295 44.825 ;
        RECT 68.150 44.640 1174.295 44.780 ;
        RECT 68.150 44.580 68.470 44.640 ;
        RECT 1174.005 44.595 1174.295 44.640 ;
      LAYER via ;
        RECT 1174.020 1635.100 1174.280 1635.360 ;
        RECT 1174.480 1587.160 1174.740 1587.420 ;
        RECT 1174.480 1538.540 1174.740 1538.800 ;
        RECT 1174.480 1490.600 1174.740 1490.860 ;
        RECT 1173.100 1297.140 1173.360 1297.400 ;
        RECT 1174.480 1297.140 1174.740 1297.400 ;
        RECT 1174.480 1256.000 1174.740 1256.260 ;
        RECT 1174.940 1255.320 1175.200 1255.580 ;
        RECT 1174.480 1207.380 1174.740 1207.640 ;
        RECT 1174.940 1207.380 1175.200 1207.640 ;
        RECT 1174.480 1200.240 1174.740 1200.500 ;
        RECT 1174.480 1152.300 1174.740 1152.560 ;
        RECT 1174.020 1014.260 1174.280 1014.520 ;
        RECT 1174.480 1014.260 1174.740 1014.520 ;
        RECT 1174.020 1007.120 1174.280 1007.380 ;
        RECT 1174.020 961.220 1174.280 961.480 ;
        RECT 1174.020 869.420 1174.280 869.680 ;
        RECT 1174.480 869.420 1174.740 869.680 ;
        RECT 1174.480 806.520 1174.740 806.780 ;
        RECT 1174.020 704.180 1174.280 704.440 ;
        RECT 1174.020 703.500 1174.280 703.760 ;
        RECT 1174.940 672.900 1175.200 673.160 ;
        RECT 1174.480 600.140 1174.740 600.400 ;
        RECT 1174.020 460.060 1174.280 460.320 ;
        RECT 1174.020 420.620 1174.280 420.880 ;
        RECT 1174.020 372.680 1174.280 372.940 ;
        RECT 1174.020 324.060 1174.280 324.320 ;
        RECT 1174.020 276.120 1174.280 276.380 ;
        RECT 1174.020 227.500 1174.280 227.760 ;
        RECT 1174.020 179.560 1174.280 179.820 ;
        RECT 1174.020 130.940 1174.280 131.200 ;
        RECT 68.180 44.580 68.440 44.840 ;
      LAYER met2 ;
        RECT 1174.405 1700.000 1174.685 1704.000 ;
        RECT 1174.540 1642.610 1174.680 1700.000 ;
        RECT 1174.080 1642.470 1174.680 1642.610 ;
        RECT 1174.080 1635.390 1174.220 1642.470 ;
        RECT 1174.020 1635.070 1174.280 1635.390 ;
        RECT 1174.480 1587.130 1174.740 1587.450 ;
        RECT 1174.540 1538.830 1174.680 1587.130 ;
        RECT 1174.480 1538.510 1174.740 1538.830 ;
        RECT 1174.480 1490.570 1174.740 1490.890 ;
        RECT 1174.540 1393.730 1174.680 1490.570 ;
        RECT 1174.080 1393.590 1174.680 1393.730 ;
        RECT 1174.080 1387.045 1174.220 1393.590 ;
        RECT 1173.090 1386.675 1173.370 1387.045 ;
        RECT 1174.010 1386.675 1174.290 1387.045 ;
        RECT 1173.160 1297.430 1173.300 1386.675 ;
        RECT 1173.100 1297.110 1173.360 1297.430 ;
        RECT 1174.480 1297.110 1174.740 1297.430 ;
        RECT 1174.540 1256.290 1174.680 1297.110 ;
        RECT 1174.480 1255.970 1174.740 1256.290 ;
        RECT 1174.940 1255.290 1175.200 1255.610 ;
        RECT 1175.000 1207.670 1175.140 1255.290 ;
        RECT 1174.480 1207.350 1174.740 1207.670 ;
        RECT 1174.940 1207.350 1175.200 1207.670 ;
        RECT 1174.540 1200.530 1174.680 1207.350 ;
        RECT 1174.480 1200.210 1174.740 1200.530 ;
        RECT 1174.480 1152.270 1174.740 1152.590 ;
        RECT 1174.540 1104.165 1174.680 1152.270 ;
        RECT 1174.470 1103.795 1174.750 1104.165 ;
        RECT 1175.850 1103.795 1176.130 1104.165 ;
        RECT 1175.920 1055.885 1176.060 1103.795 ;
        RECT 1174.470 1055.515 1174.750 1055.885 ;
        RECT 1175.850 1055.515 1176.130 1055.885 ;
        RECT 1174.540 1014.550 1174.680 1055.515 ;
        RECT 1174.020 1014.230 1174.280 1014.550 ;
        RECT 1174.480 1014.230 1174.740 1014.550 ;
        RECT 1174.080 1007.410 1174.220 1014.230 ;
        RECT 1174.020 1007.090 1174.280 1007.410 ;
        RECT 1174.020 961.190 1174.280 961.510 ;
        RECT 1174.080 869.710 1174.220 961.190 ;
        RECT 1174.020 869.390 1174.280 869.710 ;
        RECT 1174.480 869.450 1174.740 869.710 ;
        RECT 1174.480 869.390 1175.140 869.450 ;
        RECT 1174.540 869.310 1175.140 869.390 ;
        RECT 1175.000 815.730 1175.140 869.310 ;
        RECT 1175.000 815.590 1175.600 815.730 ;
        RECT 1175.460 814.485 1175.600 815.590 ;
        RECT 1174.470 814.115 1174.750 814.485 ;
        RECT 1175.390 814.115 1175.670 814.485 ;
        RECT 1174.540 806.810 1174.680 814.115 ;
        RECT 1174.480 806.490 1174.740 806.810 ;
        RECT 1174.020 704.150 1174.280 704.470 ;
        RECT 1174.080 703.790 1174.220 704.150 ;
        RECT 1174.020 703.470 1174.280 703.790 ;
        RECT 1174.940 672.870 1175.200 673.190 ;
        RECT 1175.000 607.650 1175.140 672.870 ;
        RECT 1174.540 607.510 1175.140 607.650 ;
        RECT 1174.540 600.430 1174.680 607.510 ;
        RECT 1174.480 600.110 1174.740 600.430 ;
        RECT 1174.020 460.030 1174.280 460.350 ;
        RECT 1174.080 428.925 1174.220 460.030 ;
        RECT 1174.010 428.555 1174.290 428.925 ;
        RECT 1174.010 427.875 1174.290 428.245 ;
        RECT 1174.080 420.910 1174.220 427.875 ;
        RECT 1174.020 420.590 1174.280 420.910 ;
        RECT 1174.020 372.650 1174.280 372.970 ;
        RECT 1174.080 324.350 1174.220 372.650 ;
        RECT 1174.020 324.030 1174.280 324.350 ;
        RECT 1174.020 276.090 1174.280 276.410 ;
        RECT 1174.080 227.790 1174.220 276.090 ;
        RECT 1174.020 227.470 1174.280 227.790 ;
        RECT 1174.020 179.530 1174.280 179.850 ;
        RECT 1174.080 131.230 1174.220 179.530 ;
        RECT 1174.020 130.910 1174.280 131.230 ;
        RECT 68.180 44.550 68.440 44.870 ;
        RECT 68.240 2.400 68.380 44.550 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 1173.090 1386.720 1173.370 1387.000 ;
        RECT 1174.010 1386.720 1174.290 1387.000 ;
        RECT 1174.470 1103.840 1174.750 1104.120 ;
        RECT 1175.850 1103.840 1176.130 1104.120 ;
        RECT 1174.470 1055.560 1174.750 1055.840 ;
        RECT 1175.850 1055.560 1176.130 1055.840 ;
        RECT 1174.470 814.160 1174.750 814.440 ;
        RECT 1175.390 814.160 1175.670 814.440 ;
        RECT 1174.010 428.600 1174.290 428.880 ;
        RECT 1174.010 427.920 1174.290 428.200 ;
      LAYER met3 ;
        RECT 1173.065 1387.010 1173.395 1387.025 ;
        RECT 1173.985 1387.010 1174.315 1387.025 ;
        RECT 1173.065 1386.710 1174.315 1387.010 ;
        RECT 1173.065 1386.695 1173.395 1386.710 ;
        RECT 1173.985 1386.695 1174.315 1386.710 ;
        RECT 1174.445 1104.130 1174.775 1104.145 ;
        RECT 1175.825 1104.130 1176.155 1104.145 ;
        RECT 1174.445 1103.830 1176.155 1104.130 ;
        RECT 1174.445 1103.815 1174.775 1103.830 ;
        RECT 1175.825 1103.815 1176.155 1103.830 ;
        RECT 1174.445 1055.850 1174.775 1055.865 ;
        RECT 1175.825 1055.850 1176.155 1055.865 ;
        RECT 1174.445 1055.550 1176.155 1055.850 ;
        RECT 1174.445 1055.535 1174.775 1055.550 ;
        RECT 1175.825 1055.535 1176.155 1055.550 ;
        RECT 1174.445 814.450 1174.775 814.465 ;
        RECT 1175.365 814.450 1175.695 814.465 ;
        RECT 1174.445 814.150 1175.695 814.450 ;
        RECT 1174.445 814.135 1174.775 814.150 ;
        RECT 1175.365 814.135 1175.695 814.150 ;
        RECT 1173.985 428.890 1174.315 428.905 ;
        RECT 1173.985 428.575 1174.530 428.890 ;
        RECT 1174.230 428.225 1174.530 428.575 ;
        RECT 1173.985 427.910 1174.530 428.225 ;
        RECT 1173.985 427.895 1174.315 427.910 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1306.545 766.105 1306.715 814.215 ;
        RECT 1306.085 593.045 1306.255 620.755 ;
        RECT 1306.085 241.485 1306.255 265.795 ;
        RECT 1306.085 138.125 1306.255 159.035 ;
      LAYER mcon ;
        RECT 1306.545 814.045 1306.715 814.215 ;
        RECT 1306.085 620.585 1306.255 620.755 ;
        RECT 1306.085 265.625 1306.255 265.795 ;
        RECT 1306.085 158.865 1306.255 159.035 ;
      LAYER met1 ;
        RECT 1306.010 1607.900 1306.330 1608.160 ;
        RECT 1306.100 1607.080 1306.240 1607.900 ;
        RECT 1306.470 1607.080 1306.790 1607.140 ;
        RECT 1306.100 1606.940 1306.790 1607.080 ;
        RECT 1306.470 1606.880 1306.790 1606.940 ;
        RECT 1306.010 1449.320 1306.330 1449.380 ;
        RECT 1306.470 1449.320 1306.790 1449.380 ;
        RECT 1306.010 1449.180 1306.790 1449.320 ;
        RECT 1306.010 1449.120 1306.330 1449.180 ;
        RECT 1306.470 1449.120 1306.790 1449.180 ;
        RECT 1306.010 1365.820 1306.330 1366.080 ;
        RECT 1306.100 1365.400 1306.240 1365.820 ;
        RECT 1306.010 1365.140 1306.330 1365.400 ;
        RECT 1306.010 1269.260 1306.330 1269.520 ;
        RECT 1306.100 1268.840 1306.240 1269.260 ;
        RECT 1306.010 1268.580 1306.330 1268.840 ;
        RECT 1306.010 1172.700 1306.330 1172.960 ;
        RECT 1306.100 1172.280 1306.240 1172.700 ;
        RECT 1306.010 1172.020 1306.330 1172.280 ;
        RECT 1306.010 1080.080 1306.330 1080.140 ;
        RECT 1306.930 1080.080 1307.250 1080.140 ;
        RECT 1306.010 1079.940 1307.250 1080.080 ;
        RECT 1306.010 1079.880 1306.330 1079.940 ;
        RECT 1306.930 1079.880 1307.250 1079.940 ;
        RECT 1306.010 931.980 1306.330 932.240 ;
        RECT 1306.100 931.560 1306.240 931.980 ;
        RECT 1306.010 931.300 1306.330 931.560 ;
        RECT 1306.010 869.620 1306.330 869.680 ;
        RECT 1306.470 869.620 1306.790 869.680 ;
        RECT 1306.010 869.480 1306.790 869.620 ;
        RECT 1306.010 869.420 1306.330 869.480 ;
        RECT 1306.470 869.420 1306.790 869.480 ;
        RECT 1306.485 814.200 1306.775 814.245 ;
        RECT 1306.930 814.200 1307.250 814.260 ;
        RECT 1306.485 814.060 1307.250 814.200 ;
        RECT 1306.485 814.015 1306.775 814.060 ;
        RECT 1306.930 814.000 1307.250 814.060 ;
        RECT 1306.470 766.260 1306.790 766.320 ;
        RECT 1306.275 766.120 1306.790 766.260 ;
        RECT 1306.470 766.060 1306.790 766.120 ;
        RECT 1306.025 620.740 1306.315 620.785 ;
        RECT 1306.470 620.740 1306.790 620.800 ;
        RECT 1306.025 620.600 1306.790 620.740 ;
        RECT 1306.025 620.555 1306.315 620.600 ;
        RECT 1306.470 620.540 1306.790 620.600 ;
        RECT 1306.010 593.200 1306.330 593.260 ;
        RECT 1305.815 593.060 1306.330 593.200 ;
        RECT 1306.010 593.000 1306.330 593.060 ;
        RECT 1305.550 385.940 1305.870 386.200 ;
        RECT 1305.640 385.800 1305.780 385.940 ;
        RECT 1306.470 385.800 1306.790 385.860 ;
        RECT 1305.640 385.660 1306.790 385.800 ;
        RECT 1306.470 385.600 1306.790 385.660 ;
        RECT 1306.470 304.200 1306.790 304.260 ;
        RECT 1306.100 304.060 1306.790 304.200 ;
        RECT 1306.100 303.580 1306.240 304.060 ;
        RECT 1306.470 304.000 1306.790 304.060 ;
        RECT 1306.010 303.320 1306.330 303.580 ;
        RECT 1306.010 265.780 1306.330 265.840 ;
        RECT 1305.815 265.640 1306.330 265.780 ;
        RECT 1306.010 265.580 1306.330 265.640 ;
        RECT 1306.025 241.640 1306.315 241.685 ;
        RECT 1306.470 241.640 1306.790 241.700 ;
        RECT 1306.025 241.500 1306.790 241.640 ;
        RECT 1306.025 241.455 1306.315 241.500 ;
        RECT 1306.470 241.440 1306.790 241.500 ;
        RECT 1306.010 159.020 1306.330 159.080 ;
        RECT 1305.815 158.880 1306.330 159.020 ;
        RECT 1306.010 158.820 1306.330 158.880 ;
        RECT 1306.010 138.280 1306.330 138.340 ;
        RECT 1305.815 138.140 1306.330 138.280 ;
        RECT 1306.010 138.080 1306.330 138.140 ;
        RECT 1305.550 96.800 1305.870 96.860 ;
        RECT 1306.010 96.800 1306.330 96.860 ;
        RECT 1305.550 96.660 1306.330 96.800 ;
        RECT 1305.550 96.600 1305.870 96.660 ;
        RECT 1306.010 96.600 1306.330 96.660 ;
        RECT 427.410 73.680 427.730 73.740 ;
        RECT 1305.550 73.680 1305.870 73.740 ;
        RECT 427.410 73.540 1305.870 73.680 ;
        RECT 427.410 73.480 427.730 73.540 ;
        RECT 1305.550 73.480 1305.870 73.540 ;
        RECT 424.650 16.220 424.970 16.280 ;
        RECT 427.410 16.220 427.730 16.280 ;
        RECT 424.650 16.080 427.730 16.220 ;
        RECT 424.650 16.020 424.970 16.080 ;
        RECT 427.410 16.020 427.730 16.080 ;
      LAYER via ;
        RECT 1306.040 1607.900 1306.300 1608.160 ;
        RECT 1306.500 1606.880 1306.760 1607.140 ;
        RECT 1306.040 1449.120 1306.300 1449.380 ;
        RECT 1306.500 1449.120 1306.760 1449.380 ;
        RECT 1306.040 1365.820 1306.300 1366.080 ;
        RECT 1306.040 1365.140 1306.300 1365.400 ;
        RECT 1306.040 1269.260 1306.300 1269.520 ;
        RECT 1306.040 1268.580 1306.300 1268.840 ;
        RECT 1306.040 1172.700 1306.300 1172.960 ;
        RECT 1306.040 1172.020 1306.300 1172.280 ;
        RECT 1306.040 1079.880 1306.300 1080.140 ;
        RECT 1306.960 1079.880 1307.220 1080.140 ;
        RECT 1306.040 931.980 1306.300 932.240 ;
        RECT 1306.040 931.300 1306.300 931.560 ;
        RECT 1306.040 869.420 1306.300 869.680 ;
        RECT 1306.500 869.420 1306.760 869.680 ;
        RECT 1306.960 814.000 1307.220 814.260 ;
        RECT 1306.500 766.060 1306.760 766.320 ;
        RECT 1306.500 620.540 1306.760 620.800 ;
        RECT 1306.040 593.000 1306.300 593.260 ;
        RECT 1305.580 385.940 1305.840 386.200 ;
        RECT 1306.500 385.600 1306.760 385.860 ;
        RECT 1306.500 304.000 1306.760 304.260 ;
        RECT 1306.040 303.320 1306.300 303.580 ;
        RECT 1306.040 265.580 1306.300 265.840 ;
        RECT 1306.500 241.440 1306.760 241.700 ;
        RECT 1306.040 158.820 1306.300 159.080 ;
        RECT 1306.040 138.080 1306.300 138.340 ;
        RECT 1305.580 96.600 1305.840 96.860 ;
        RECT 1306.040 96.600 1306.300 96.860 ;
        RECT 427.440 73.480 427.700 73.740 ;
        RECT 1305.580 73.480 1305.840 73.740 ;
        RECT 424.680 16.020 424.940 16.280 ;
        RECT 427.440 16.020 427.700 16.280 ;
      LAYER met2 ;
        RECT 1309.185 1700.410 1309.465 1704.000 ;
        RECT 1307.940 1700.270 1309.465 1700.410 ;
        RECT 1307.940 1656.210 1308.080 1700.270 ;
        RECT 1309.185 1700.000 1309.465 1700.270 ;
        RECT 1306.100 1656.070 1308.080 1656.210 ;
        RECT 1306.100 1608.190 1306.240 1656.070 ;
        RECT 1306.040 1607.870 1306.300 1608.190 ;
        RECT 1306.500 1606.850 1306.760 1607.170 ;
        RECT 1306.560 1449.410 1306.700 1606.850 ;
        RECT 1306.040 1449.090 1306.300 1449.410 ;
        RECT 1306.500 1449.090 1306.760 1449.410 ;
        RECT 1306.100 1366.110 1306.240 1449.090 ;
        RECT 1306.040 1365.790 1306.300 1366.110 ;
        RECT 1306.040 1365.110 1306.300 1365.430 ;
        RECT 1306.100 1269.550 1306.240 1365.110 ;
        RECT 1306.040 1269.230 1306.300 1269.550 ;
        RECT 1306.040 1268.550 1306.300 1268.870 ;
        RECT 1306.100 1172.990 1306.240 1268.550 ;
        RECT 1306.040 1172.670 1306.300 1172.990 ;
        RECT 1306.040 1171.990 1306.300 1172.310 ;
        RECT 1306.100 1080.170 1306.240 1171.990 ;
        RECT 1306.040 1079.850 1306.300 1080.170 ;
        RECT 1306.960 1079.850 1307.220 1080.170 ;
        RECT 1307.020 1055.885 1307.160 1079.850 ;
        RECT 1306.030 1055.515 1306.310 1055.885 ;
        RECT 1306.950 1055.515 1307.230 1055.885 ;
        RECT 1306.100 932.270 1306.240 1055.515 ;
        RECT 1306.040 931.950 1306.300 932.270 ;
        RECT 1306.040 931.270 1306.300 931.590 ;
        RECT 1306.100 869.710 1306.240 931.270 ;
        RECT 1306.040 869.390 1306.300 869.710 ;
        RECT 1306.500 869.390 1306.760 869.710 ;
        RECT 1306.560 855.170 1306.700 869.390 ;
        RECT 1306.560 855.030 1307.160 855.170 ;
        RECT 1307.020 814.290 1307.160 855.030 ;
        RECT 1306.960 813.970 1307.220 814.290 ;
        RECT 1306.500 766.030 1306.760 766.350 ;
        RECT 1306.560 669.530 1306.700 766.030 ;
        RECT 1306.560 669.390 1307.160 669.530 ;
        RECT 1307.020 628.845 1307.160 669.390 ;
        RECT 1306.950 628.475 1307.230 628.845 ;
        RECT 1306.490 627.795 1306.770 628.165 ;
        RECT 1306.560 620.830 1306.700 627.795 ;
        RECT 1306.500 620.510 1306.760 620.830 ;
        RECT 1306.040 592.970 1306.300 593.290 ;
        RECT 1306.100 497.490 1306.240 592.970 ;
        RECT 1305.640 497.350 1306.240 497.490 ;
        RECT 1305.640 496.810 1305.780 497.350 ;
        RECT 1305.640 496.670 1306.240 496.810 ;
        RECT 1306.100 411.130 1306.240 496.670 ;
        RECT 1305.640 410.990 1306.240 411.130 ;
        RECT 1305.640 386.230 1305.780 410.990 ;
        RECT 1305.580 385.910 1305.840 386.230 ;
        RECT 1306.500 385.570 1306.760 385.890 ;
        RECT 1306.560 304.290 1306.700 385.570 ;
        RECT 1306.500 303.970 1306.760 304.290 ;
        RECT 1306.040 303.290 1306.300 303.610 ;
        RECT 1306.100 265.870 1306.240 303.290 ;
        RECT 1306.040 265.550 1306.300 265.870 ;
        RECT 1306.500 241.410 1306.760 241.730 ;
        RECT 1306.560 186.730 1306.700 241.410 ;
        RECT 1306.100 186.590 1306.700 186.730 ;
        RECT 1306.100 159.110 1306.240 186.590 ;
        RECT 1306.040 158.790 1306.300 159.110 ;
        RECT 1306.040 138.050 1306.300 138.370 ;
        RECT 1306.100 96.890 1306.240 138.050 ;
        RECT 1305.580 96.570 1305.840 96.890 ;
        RECT 1306.040 96.570 1306.300 96.890 ;
        RECT 1305.640 73.770 1305.780 96.570 ;
        RECT 427.440 73.450 427.700 73.770 ;
        RECT 1305.580 73.450 1305.840 73.770 ;
        RECT 427.500 16.310 427.640 73.450 ;
        RECT 424.680 15.990 424.940 16.310 ;
        RECT 427.440 15.990 427.700 16.310 ;
        RECT 424.740 2.400 424.880 15.990 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 1306.030 1055.560 1306.310 1055.840 ;
        RECT 1306.950 1055.560 1307.230 1055.840 ;
        RECT 1306.950 628.520 1307.230 628.800 ;
        RECT 1306.490 627.840 1306.770 628.120 ;
      LAYER met3 ;
        RECT 1306.005 1055.850 1306.335 1055.865 ;
        RECT 1306.925 1055.850 1307.255 1055.865 ;
        RECT 1306.005 1055.550 1307.255 1055.850 ;
        RECT 1306.005 1055.535 1306.335 1055.550 ;
        RECT 1306.925 1055.535 1307.255 1055.550 ;
        RECT 1306.925 628.810 1307.255 628.825 ;
        RECT 1306.710 628.495 1307.255 628.810 ;
        RECT 1306.710 628.145 1307.010 628.495 ;
        RECT 1306.465 627.830 1307.010 628.145 ;
        RECT 1306.465 627.815 1306.795 627.830 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1313.445 1560.685 1313.615 1593.835 ;
        RECT 1312.985 1449.505 1313.155 1497.275 ;
        RECT 1312.525 1394.085 1312.695 1441.855 ;
        RECT 1312.525 1317.245 1312.695 1393.575 ;
        RECT 1312.985 1256.045 1313.155 1304.155 ;
        RECT 1312.985 917.405 1313.155 959.055 ;
        RECT 1312.525 766.105 1312.695 814.215 ;
        RECT 1313.445 648.805 1313.615 696.915 ;
        RECT 1313.445 510.765 1313.615 600.355 ;
        RECT 1312.525 434.605 1312.695 497.335 ;
        RECT 1313.905 331.245 1314.075 379.355 ;
        RECT 1314.365 186.405 1314.535 234.515 ;
        RECT 1312.985 96.645 1313.155 120.955 ;
      LAYER mcon ;
        RECT 1313.445 1593.665 1313.615 1593.835 ;
        RECT 1312.985 1497.105 1313.155 1497.275 ;
        RECT 1312.525 1441.685 1312.695 1441.855 ;
        RECT 1312.525 1393.405 1312.695 1393.575 ;
        RECT 1312.985 1303.985 1313.155 1304.155 ;
        RECT 1312.985 958.885 1313.155 959.055 ;
        RECT 1312.525 814.045 1312.695 814.215 ;
        RECT 1313.445 696.745 1313.615 696.915 ;
        RECT 1313.445 600.185 1313.615 600.355 ;
        RECT 1312.525 497.165 1312.695 497.335 ;
        RECT 1313.905 379.185 1314.075 379.355 ;
        RECT 1314.365 234.345 1314.535 234.515 ;
        RECT 1312.985 120.785 1313.155 120.955 ;
      LAYER met1 ;
        RECT 1313.370 1642.440 1313.690 1642.500 ;
        RECT 1315.210 1642.440 1315.530 1642.500 ;
        RECT 1313.370 1642.300 1315.530 1642.440 ;
        RECT 1313.370 1642.240 1313.690 1642.300 ;
        RECT 1315.210 1642.240 1315.530 1642.300 ;
        RECT 1313.370 1593.820 1313.690 1593.880 ;
        RECT 1313.175 1593.680 1313.690 1593.820 ;
        RECT 1313.370 1593.620 1313.690 1593.680 ;
        RECT 1313.370 1560.840 1313.690 1560.900 ;
        RECT 1313.175 1560.700 1313.690 1560.840 ;
        RECT 1313.370 1560.640 1313.690 1560.700 ;
        RECT 1312.925 1497.260 1313.215 1497.305 ;
        RECT 1313.370 1497.260 1313.690 1497.320 ;
        RECT 1312.925 1497.120 1313.690 1497.260 ;
        RECT 1312.925 1497.075 1313.215 1497.120 ;
        RECT 1313.370 1497.060 1313.690 1497.120 ;
        RECT 1312.910 1449.660 1313.230 1449.720 ;
        RECT 1312.715 1449.520 1313.230 1449.660 ;
        RECT 1312.910 1449.460 1313.230 1449.520 ;
        RECT 1312.465 1441.840 1312.755 1441.885 ;
        RECT 1312.910 1441.840 1313.230 1441.900 ;
        RECT 1312.465 1441.700 1313.230 1441.840 ;
        RECT 1312.465 1441.655 1312.755 1441.700 ;
        RECT 1312.910 1441.640 1313.230 1441.700 ;
        RECT 1312.450 1394.240 1312.770 1394.300 ;
        RECT 1312.255 1394.100 1312.770 1394.240 ;
        RECT 1312.450 1394.040 1312.770 1394.100 ;
        RECT 1312.450 1393.560 1312.770 1393.620 ;
        RECT 1312.255 1393.420 1312.770 1393.560 ;
        RECT 1312.450 1393.360 1312.770 1393.420 ;
        RECT 1312.465 1317.400 1312.755 1317.445 ;
        RECT 1313.370 1317.400 1313.690 1317.460 ;
        RECT 1312.465 1317.260 1313.690 1317.400 ;
        RECT 1312.465 1317.215 1312.755 1317.260 ;
        RECT 1313.370 1317.200 1313.690 1317.260 ;
        RECT 1312.925 1304.140 1313.215 1304.185 ;
        RECT 1313.370 1304.140 1313.690 1304.200 ;
        RECT 1312.925 1304.000 1313.690 1304.140 ;
        RECT 1312.925 1303.955 1313.215 1304.000 ;
        RECT 1313.370 1303.940 1313.690 1304.000 ;
        RECT 1312.910 1256.200 1313.230 1256.260 ;
        RECT 1312.715 1256.060 1313.230 1256.200 ;
        RECT 1312.910 1256.000 1313.230 1256.060 ;
        RECT 1313.830 1207.580 1314.150 1207.640 ;
        RECT 1314.290 1207.580 1314.610 1207.640 ;
        RECT 1313.830 1207.440 1314.610 1207.580 ;
        RECT 1313.830 1207.380 1314.150 1207.440 ;
        RECT 1314.290 1207.380 1314.610 1207.440 ;
        RECT 1312.910 1159.300 1313.230 1159.360 ;
        RECT 1314.290 1159.300 1314.610 1159.360 ;
        RECT 1312.910 1159.160 1314.610 1159.300 ;
        RECT 1312.910 1159.100 1313.230 1159.160 ;
        RECT 1314.290 1159.100 1314.610 1159.160 ;
        RECT 1312.450 1111.020 1312.770 1111.080 ;
        RECT 1314.290 1111.020 1314.610 1111.080 ;
        RECT 1312.450 1110.880 1314.610 1111.020 ;
        RECT 1312.450 1110.820 1312.770 1110.880 ;
        RECT 1314.290 1110.820 1314.610 1110.880 ;
        RECT 1312.910 1062.740 1313.230 1062.800 ;
        RECT 1314.290 1062.740 1314.610 1062.800 ;
        RECT 1312.910 1062.600 1314.610 1062.740 ;
        RECT 1312.910 1062.540 1313.230 1062.600 ;
        RECT 1314.290 1062.540 1314.610 1062.600 ;
        RECT 1312.910 966.660 1313.230 966.920 ;
        RECT 1313.000 966.240 1313.140 966.660 ;
        RECT 1312.910 965.980 1313.230 966.240 ;
        RECT 1312.910 959.040 1313.230 959.100 ;
        RECT 1312.715 958.900 1313.230 959.040 ;
        RECT 1312.910 958.840 1313.230 958.900 ;
        RECT 1312.910 917.560 1313.230 917.620 ;
        RECT 1312.715 917.420 1313.230 917.560 ;
        RECT 1312.910 917.360 1313.230 917.420 ;
        RECT 1313.370 869.420 1313.690 869.680 ;
        RECT 1313.460 868.940 1313.600 869.420 ;
        RECT 1313.830 868.940 1314.150 869.000 ;
        RECT 1313.460 868.800 1314.150 868.940 ;
        RECT 1313.830 868.740 1314.150 868.800 ;
        RECT 1313.370 821.340 1313.690 821.400 ;
        RECT 1313.830 821.340 1314.150 821.400 ;
        RECT 1313.370 821.200 1314.150 821.340 ;
        RECT 1313.370 821.140 1313.690 821.200 ;
        RECT 1313.830 821.140 1314.150 821.200 ;
        RECT 1312.465 814.200 1312.755 814.245 ;
        RECT 1313.370 814.200 1313.690 814.260 ;
        RECT 1312.465 814.060 1313.690 814.200 ;
        RECT 1312.465 814.015 1312.755 814.060 ;
        RECT 1313.370 814.000 1313.690 814.060 ;
        RECT 1312.450 766.260 1312.770 766.320 ;
        RECT 1312.255 766.120 1312.770 766.260 ;
        RECT 1312.450 766.060 1312.770 766.120 ;
        RECT 1313.370 696.900 1313.690 696.960 ;
        RECT 1313.175 696.760 1313.690 696.900 ;
        RECT 1313.370 696.700 1313.690 696.760 ;
        RECT 1313.385 648.960 1313.675 649.005 ;
        RECT 1314.290 648.960 1314.610 649.020 ;
        RECT 1313.385 648.820 1314.610 648.960 ;
        RECT 1313.385 648.775 1313.675 648.820 ;
        RECT 1314.290 648.760 1314.610 648.820 ;
        RECT 1313.385 600.340 1313.675 600.385 ;
        RECT 1314.290 600.340 1314.610 600.400 ;
        RECT 1313.385 600.200 1314.610 600.340 ;
        RECT 1313.385 600.155 1313.675 600.200 ;
        RECT 1314.290 600.140 1314.610 600.200 ;
        RECT 1313.370 510.920 1313.690 510.980 ;
        RECT 1313.175 510.780 1313.690 510.920 ;
        RECT 1313.370 510.720 1313.690 510.780 ;
        RECT 1312.465 497.320 1312.755 497.365 ;
        RECT 1313.370 497.320 1313.690 497.380 ;
        RECT 1312.465 497.180 1313.690 497.320 ;
        RECT 1312.465 497.135 1312.755 497.180 ;
        RECT 1313.370 497.120 1313.690 497.180 ;
        RECT 1312.450 434.760 1312.770 434.820 ;
        RECT 1312.255 434.620 1312.770 434.760 ;
        RECT 1312.450 434.560 1312.770 434.620 ;
        RECT 1312.450 386.140 1312.770 386.200 ;
        RECT 1314.290 386.140 1314.610 386.200 ;
        RECT 1312.450 386.000 1314.610 386.140 ;
        RECT 1312.450 385.940 1312.770 386.000 ;
        RECT 1314.290 385.940 1314.610 386.000 ;
        RECT 1313.845 379.340 1314.135 379.385 ;
        RECT 1314.290 379.340 1314.610 379.400 ;
        RECT 1313.845 379.200 1314.610 379.340 ;
        RECT 1313.845 379.155 1314.135 379.200 ;
        RECT 1314.290 379.140 1314.610 379.200 ;
        RECT 1313.830 331.400 1314.150 331.460 ;
        RECT 1313.635 331.260 1314.150 331.400 ;
        RECT 1313.830 331.200 1314.150 331.260 ;
        RECT 1313.370 283.120 1313.690 283.180 ;
        RECT 1314.290 283.120 1314.610 283.180 ;
        RECT 1313.370 282.980 1314.610 283.120 ;
        RECT 1313.370 282.920 1313.690 282.980 ;
        RECT 1314.290 282.920 1314.610 282.980 ;
        RECT 1313.370 282.440 1313.690 282.500 ;
        RECT 1314.290 282.440 1314.610 282.500 ;
        RECT 1313.370 282.300 1314.610 282.440 ;
        RECT 1313.370 282.240 1313.690 282.300 ;
        RECT 1314.290 282.240 1314.610 282.300 ;
        RECT 1314.290 234.500 1314.610 234.560 ;
        RECT 1314.290 234.360 1314.805 234.500 ;
        RECT 1314.290 234.300 1314.610 234.360 ;
        RECT 1313.370 186.560 1313.690 186.620 ;
        RECT 1314.305 186.560 1314.595 186.605 ;
        RECT 1313.370 186.420 1314.595 186.560 ;
        RECT 1313.370 186.360 1313.690 186.420 ;
        RECT 1314.305 186.375 1314.595 186.420 ;
        RECT 1312.925 120.940 1313.215 120.985 ;
        RECT 1313.370 120.940 1313.690 121.000 ;
        RECT 1312.925 120.800 1313.690 120.940 ;
        RECT 1312.925 120.755 1313.215 120.800 ;
        RECT 1313.370 120.740 1313.690 120.800 ;
        RECT 1312.910 96.800 1313.230 96.860 ;
        RECT 1312.715 96.660 1313.230 96.800 ;
        RECT 1312.910 96.600 1313.230 96.660 ;
        RECT 448.110 74.020 448.430 74.080 ;
        RECT 1312.910 74.020 1313.230 74.080 ;
        RECT 448.110 73.880 1313.230 74.020 ;
        RECT 448.110 73.820 448.430 73.880 ;
        RECT 1312.910 73.820 1313.230 73.880 ;
        RECT 442.590 16.220 442.910 16.280 ;
        RECT 448.110 16.220 448.430 16.280 ;
        RECT 442.590 16.080 448.430 16.220 ;
        RECT 442.590 16.020 442.910 16.080 ;
        RECT 448.110 16.020 448.430 16.080 ;
      LAYER via ;
        RECT 1313.400 1642.240 1313.660 1642.500 ;
        RECT 1315.240 1642.240 1315.500 1642.500 ;
        RECT 1313.400 1593.620 1313.660 1593.880 ;
        RECT 1313.400 1560.640 1313.660 1560.900 ;
        RECT 1313.400 1497.060 1313.660 1497.320 ;
        RECT 1312.940 1449.460 1313.200 1449.720 ;
        RECT 1312.940 1441.640 1313.200 1441.900 ;
        RECT 1312.480 1394.040 1312.740 1394.300 ;
        RECT 1312.480 1393.360 1312.740 1393.620 ;
        RECT 1313.400 1317.200 1313.660 1317.460 ;
        RECT 1313.400 1303.940 1313.660 1304.200 ;
        RECT 1312.940 1256.000 1313.200 1256.260 ;
        RECT 1313.860 1207.380 1314.120 1207.640 ;
        RECT 1314.320 1207.380 1314.580 1207.640 ;
        RECT 1312.940 1159.100 1313.200 1159.360 ;
        RECT 1314.320 1159.100 1314.580 1159.360 ;
        RECT 1312.480 1110.820 1312.740 1111.080 ;
        RECT 1314.320 1110.820 1314.580 1111.080 ;
        RECT 1312.940 1062.540 1313.200 1062.800 ;
        RECT 1314.320 1062.540 1314.580 1062.800 ;
        RECT 1312.940 966.660 1313.200 966.920 ;
        RECT 1312.940 965.980 1313.200 966.240 ;
        RECT 1312.940 958.840 1313.200 959.100 ;
        RECT 1312.940 917.360 1313.200 917.620 ;
        RECT 1313.400 869.420 1313.660 869.680 ;
        RECT 1313.860 868.740 1314.120 869.000 ;
        RECT 1313.400 821.140 1313.660 821.400 ;
        RECT 1313.860 821.140 1314.120 821.400 ;
        RECT 1313.400 814.000 1313.660 814.260 ;
        RECT 1312.480 766.060 1312.740 766.320 ;
        RECT 1313.400 696.700 1313.660 696.960 ;
        RECT 1314.320 648.760 1314.580 649.020 ;
        RECT 1314.320 600.140 1314.580 600.400 ;
        RECT 1313.400 510.720 1313.660 510.980 ;
        RECT 1313.400 497.120 1313.660 497.380 ;
        RECT 1312.480 434.560 1312.740 434.820 ;
        RECT 1312.480 385.940 1312.740 386.200 ;
        RECT 1314.320 385.940 1314.580 386.200 ;
        RECT 1314.320 379.140 1314.580 379.400 ;
        RECT 1313.860 331.200 1314.120 331.460 ;
        RECT 1313.400 282.920 1313.660 283.180 ;
        RECT 1314.320 282.920 1314.580 283.180 ;
        RECT 1313.400 282.240 1313.660 282.500 ;
        RECT 1314.320 282.240 1314.580 282.500 ;
        RECT 1314.320 234.300 1314.580 234.560 ;
        RECT 1313.400 186.360 1313.660 186.620 ;
        RECT 1313.400 120.740 1313.660 121.000 ;
        RECT 1312.940 96.600 1313.200 96.860 ;
        RECT 448.140 73.820 448.400 74.080 ;
        RECT 1312.940 73.820 1313.200 74.080 ;
        RECT 442.620 16.020 442.880 16.280 ;
        RECT 448.140 16.020 448.400 16.280 ;
      LAYER met2 ;
        RECT 1316.085 1700.410 1316.365 1704.000 ;
        RECT 1315.300 1700.270 1316.365 1700.410 ;
        RECT 1315.300 1642.530 1315.440 1700.270 ;
        RECT 1316.085 1700.000 1316.365 1700.270 ;
        RECT 1313.400 1642.210 1313.660 1642.530 ;
        RECT 1315.240 1642.210 1315.500 1642.530 ;
        RECT 1313.460 1593.910 1313.600 1642.210 ;
        RECT 1313.400 1593.590 1313.660 1593.910 ;
        RECT 1313.400 1560.610 1313.660 1560.930 ;
        RECT 1313.460 1497.350 1313.600 1560.610 ;
        RECT 1313.400 1497.030 1313.660 1497.350 ;
        RECT 1312.940 1449.430 1313.200 1449.750 ;
        RECT 1313.000 1441.930 1313.140 1449.430 ;
        RECT 1312.940 1441.610 1313.200 1441.930 ;
        RECT 1312.480 1394.010 1312.740 1394.330 ;
        RECT 1312.540 1393.650 1312.680 1394.010 ;
        RECT 1312.480 1393.330 1312.740 1393.650 ;
        RECT 1313.400 1317.170 1313.660 1317.490 ;
        RECT 1313.460 1304.230 1313.600 1317.170 ;
        RECT 1313.400 1303.910 1313.660 1304.230 ;
        RECT 1312.940 1255.970 1313.200 1256.290 ;
        RECT 1313.000 1231.890 1313.140 1255.970 ;
        RECT 1313.000 1231.750 1314.060 1231.890 ;
        RECT 1313.920 1207.670 1314.060 1231.750 ;
        RECT 1313.860 1207.350 1314.120 1207.670 ;
        RECT 1314.320 1207.350 1314.580 1207.670 ;
        RECT 1314.380 1159.390 1314.520 1207.350 ;
        RECT 1312.940 1159.070 1313.200 1159.390 ;
        RECT 1314.320 1159.070 1314.580 1159.390 ;
        RECT 1313.000 1135.330 1313.140 1159.070 ;
        RECT 1312.540 1135.190 1313.140 1135.330 ;
        RECT 1312.540 1111.110 1312.680 1135.190 ;
        RECT 1312.480 1110.790 1312.740 1111.110 ;
        RECT 1314.320 1110.790 1314.580 1111.110 ;
        RECT 1314.380 1062.830 1314.520 1110.790 ;
        RECT 1312.940 1062.510 1313.200 1062.830 ;
        RECT 1314.320 1062.510 1314.580 1062.830 ;
        RECT 1313.000 966.950 1313.140 1062.510 ;
        RECT 1312.940 966.630 1313.200 966.950 ;
        RECT 1312.940 965.950 1313.200 966.270 ;
        RECT 1313.000 959.130 1313.140 965.950 ;
        RECT 1312.940 958.810 1313.200 959.130 ;
        RECT 1312.940 917.330 1313.200 917.650 ;
        RECT 1313.000 910.930 1313.140 917.330 ;
        RECT 1313.000 910.790 1313.600 910.930 ;
        RECT 1313.460 869.710 1313.600 910.790 ;
        RECT 1313.400 869.390 1313.660 869.710 ;
        RECT 1313.860 868.710 1314.120 869.030 ;
        RECT 1313.920 821.430 1314.060 868.710 ;
        RECT 1313.400 821.110 1313.660 821.430 ;
        RECT 1313.860 821.110 1314.120 821.430 ;
        RECT 1313.460 814.290 1313.600 821.110 ;
        RECT 1313.400 813.970 1313.660 814.290 ;
        RECT 1312.480 766.030 1312.740 766.350 ;
        RECT 1312.540 724.725 1312.680 766.030 ;
        RECT 1312.470 724.355 1312.750 724.725 ;
        RECT 1313.390 724.355 1313.670 724.725 ;
        RECT 1313.460 696.990 1313.600 724.355 ;
        RECT 1313.400 696.670 1313.660 696.990 ;
        RECT 1314.320 648.730 1314.580 649.050 ;
        RECT 1314.380 600.430 1314.520 648.730 ;
        RECT 1314.320 600.110 1314.580 600.430 ;
        RECT 1313.400 510.690 1313.660 511.010 ;
        RECT 1313.460 497.410 1313.600 510.690 ;
        RECT 1313.400 497.090 1313.660 497.410 ;
        RECT 1312.480 434.530 1312.740 434.850 ;
        RECT 1312.540 386.230 1312.680 434.530 ;
        RECT 1312.480 385.910 1312.740 386.230 ;
        RECT 1314.320 385.910 1314.580 386.230 ;
        RECT 1314.380 379.430 1314.520 385.910 ;
        RECT 1314.320 379.110 1314.580 379.430 ;
        RECT 1313.860 331.170 1314.120 331.490 ;
        RECT 1313.920 330.890 1314.060 331.170 ;
        RECT 1313.920 330.750 1314.520 330.890 ;
        RECT 1314.380 283.210 1314.520 330.750 ;
        RECT 1313.400 282.890 1313.660 283.210 ;
        RECT 1314.320 282.890 1314.580 283.210 ;
        RECT 1313.460 282.530 1313.600 282.890 ;
        RECT 1313.400 282.210 1313.660 282.530 ;
        RECT 1314.320 282.210 1314.580 282.530 ;
        RECT 1314.380 234.590 1314.520 282.210 ;
        RECT 1314.320 234.270 1314.580 234.590 ;
        RECT 1313.400 186.330 1313.660 186.650 ;
        RECT 1313.460 121.030 1313.600 186.330 ;
        RECT 1313.400 120.710 1313.660 121.030 ;
        RECT 1312.940 96.570 1313.200 96.890 ;
        RECT 1313.000 74.110 1313.140 96.570 ;
        RECT 448.140 73.790 448.400 74.110 ;
        RECT 1312.940 73.790 1313.200 74.110 ;
        RECT 448.200 16.310 448.340 73.790 ;
        RECT 442.620 15.990 442.880 16.310 ;
        RECT 448.140 15.990 448.400 16.310 ;
        RECT 442.680 2.400 442.820 15.990 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 1312.470 724.400 1312.750 724.680 ;
        RECT 1313.390 724.400 1313.670 724.680 ;
      LAYER met3 ;
        RECT 1312.445 724.690 1312.775 724.705 ;
        RECT 1313.365 724.690 1313.695 724.705 ;
        RECT 1312.445 724.390 1313.695 724.690 ;
        RECT 1312.445 724.375 1312.775 724.390 ;
        RECT 1313.365 724.375 1313.695 724.390 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1318.430 1678.140 1318.750 1678.200 ;
        RECT 1321.190 1678.140 1321.510 1678.200 ;
        RECT 1318.430 1678.000 1321.510 1678.140 ;
        RECT 1318.430 1677.940 1318.750 1678.000 ;
        RECT 1321.190 1677.940 1321.510 1678.000 ;
        RECT 461.910 74.360 462.230 74.420 ;
        RECT 1318.430 74.360 1318.750 74.420 ;
        RECT 461.910 74.220 1318.750 74.360 ;
        RECT 461.910 74.160 462.230 74.220 ;
        RECT 1318.430 74.160 1318.750 74.220 ;
      LAYER via ;
        RECT 1318.460 1677.940 1318.720 1678.200 ;
        RECT 1321.220 1677.940 1321.480 1678.200 ;
        RECT 461.940 74.160 462.200 74.420 ;
        RECT 1318.460 74.160 1318.720 74.420 ;
      LAYER met2 ;
        RECT 1322.525 1700.410 1322.805 1704.000 ;
        RECT 1321.280 1700.270 1322.805 1700.410 ;
        RECT 1321.280 1678.230 1321.420 1700.270 ;
        RECT 1322.525 1700.000 1322.805 1700.270 ;
        RECT 1318.460 1677.910 1318.720 1678.230 ;
        RECT 1321.220 1677.910 1321.480 1678.230 ;
        RECT 1318.520 74.450 1318.660 1677.910 ;
        RECT 461.940 74.130 462.200 74.450 ;
        RECT 1318.460 74.130 1318.720 74.450 ;
        RECT 462.000 17.410 462.140 74.130 ;
        RECT 460.620 17.270 462.140 17.410 ;
        RECT 460.620 2.400 460.760 17.270 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1325.330 1671.680 1325.650 1671.740 ;
        RECT 1327.630 1671.680 1327.950 1671.740 ;
        RECT 1325.330 1671.540 1327.950 1671.680 ;
        RECT 1325.330 1671.480 1325.650 1671.540 ;
        RECT 1327.630 1671.480 1327.950 1671.540 ;
        RECT 482.610 74.700 482.930 74.760 ;
        RECT 1325.330 74.700 1325.650 74.760 ;
        RECT 482.610 74.560 1325.650 74.700 ;
        RECT 482.610 74.500 482.930 74.560 ;
        RECT 1325.330 74.500 1325.650 74.560 ;
        RECT 478.470 15.540 478.790 15.600 ;
        RECT 482.610 15.540 482.930 15.600 ;
        RECT 478.470 15.400 482.930 15.540 ;
        RECT 478.470 15.340 478.790 15.400 ;
        RECT 482.610 15.340 482.930 15.400 ;
      LAYER via ;
        RECT 1325.360 1671.480 1325.620 1671.740 ;
        RECT 1327.660 1671.480 1327.920 1671.740 ;
        RECT 482.640 74.500 482.900 74.760 ;
        RECT 1325.360 74.500 1325.620 74.760 ;
        RECT 478.500 15.340 478.760 15.600 ;
        RECT 482.640 15.340 482.900 15.600 ;
      LAYER met2 ;
        RECT 1329.425 1700.410 1329.705 1704.000 ;
        RECT 1327.720 1700.270 1329.705 1700.410 ;
        RECT 1327.720 1671.770 1327.860 1700.270 ;
        RECT 1329.425 1700.000 1329.705 1700.270 ;
        RECT 1325.360 1671.450 1325.620 1671.770 ;
        RECT 1327.660 1671.450 1327.920 1671.770 ;
        RECT 1325.420 74.790 1325.560 1671.450 ;
        RECT 482.640 74.470 482.900 74.790 ;
        RECT 1325.360 74.470 1325.620 74.790 ;
        RECT 482.700 15.630 482.840 74.470 ;
        RECT 478.500 15.310 478.760 15.630 ;
        RECT 482.640 15.310 482.900 15.630 ;
        RECT 478.560 2.400 478.700 15.310 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1332.230 1678.140 1332.550 1678.200 ;
        RECT 1334.990 1678.140 1335.310 1678.200 ;
        RECT 1332.230 1678.000 1335.310 1678.140 ;
        RECT 1332.230 1677.940 1332.550 1678.000 ;
        RECT 1334.990 1677.940 1335.310 1678.000 ;
        RECT 496.410 75.040 496.730 75.100 ;
        RECT 1332.230 75.040 1332.550 75.100 ;
        RECT 496.410 74.900 1332.550 75.040 ;
        RECT 496.410 74.840 496.730 74.900 ;
        RECT 1332.230 74.840 1332.550 74.900 ;
      LAYER via ;
        RECT 1332.260 1677.940 1332.520 1678.200 ;
        RECT 1335.020 1677.940 1335.280 1678.200 ;
        RECT 496.440 74.840 496.700 75.100 ;
        RECT 1332.260 74.840 1332.520 75.100 ;
      LAYER met2 ;
        RECT 1336.325 1700.410 1336.605 1704.000 ;
        RECT 1335.080 1700.270 1336.605 1700.410 ;
        RECT 1335.080 1678.230 1335.220 1700.270 ;
        RECT 1336.325 1700.000 1336.605 1700.270 ;
        RECT 1332.260 1677.910 1332.520 1678.230 ;
        RECT 1335.020 1677.910 1335.280 1678.230 ;
        RECT 1332.320 75.130 1332.460 1677.910 ;
        RECT 496.440 74.810 496.700 75.130 ;
        RECT 1332.260 74.810 1332.520 75.130 ;
        RECT 496.500 2.400 496.640 74.810 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1339.130 1678.140 1339.450 1678.200 ;
        RECT 1341.430 1678.140 1341.750 1678.200 ;
        RECT 1339.130 1678.000 1341.750 1678.140 ;
        RECT 1339.130 1677.940 1339.450 1678.000 ;
        RECT 1341.430 1677.940 1341.750 1678.000 ;
        RECT 517.110 75.380 517.430 75.440 ;
        RECT 1339.130 75.380 1339.450 75.440 ;
        RECT 517.110 75.240 1339.450 75.380 ;
        RECT 517.110 75.180 517.430 75.240 ;
        RECT 1339.130 75.180 1339.450 75.240 ;
        RECT 513.890 15.540 514.210 15.600 ;
        RECT 517.110 15.540 517.430 15.600 ;
        RECT 513.890 15.400 517.430 15.540 ;
        RECT 513.890 15.340 514.210 15.400 ;
        RECT 517.110 15.340 517.430 15.400 ;
      LAYER via ;
        RECT 1339.160 1677.940 1339.420 1678.200 ;
        RECT 1341.460 1677.940 1341.720 1678.200 ;
        RECT 517.140 75.180 517.400 75.440 ;
        RECT 1339.160 75.180 1339.420 75.440 ;
        RECT 513.920 15.340 514.180 15.600 ;
        RECT 517.140 15.340 517.400 15.600 ;
      LAYER met2 ;
        RECT 1342.765 1700.410 1343.045 1704.000 ;
        RECT 1341.520 1700.270 1343.045 1700.410 ;
        RECT 1341.520 1678.230 1341.660 1700.270 ;
        RECT 1342.765 1700.000 1343.045 1700.270 ;
        RECT 1339.160 1677.910 1339.420 1678.230 ;
        RECT 1341.460 1677.910 1341.720 1678.230 ;
        RECT 1339.220 75.470 1339.360 1677.910 ;
        RECT 517.140 75.150 517.400 75.470 ;
        RECT 1339.160 75.150 1339.420 75.470 ;
        RECT 517.200 15.630 517.340 75.150 ;
        RECT 513.920 15.310 514.180 15.630 ;
        RECT 517.140 15.310 517.400 15.630 ;
        RECT 513.980 2.400 514.120 15.310 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.030 1678.140 1346.350 1678.200 ;
        RECT 1347.870 1678.140 1348.190 1678.200 ;
        RECT 1346.030 1678.000 1348.190 1678.140 ;
        RECT 1346.030 1677.940 1346.350 1678.000 ;
        RECT 1347.870 1677.940 1348.190 1678.000 ;
        RECT 537.350 75.720 537.670 75.780 ;
        RECT 1346.030 75.720 1346.350 75.780 ;
        RECT 537.350 75.580 1346.350 75.720 ;
        RECT 537.350 75.520 537.670 75.580 ;
        RECT 1346.030 75.520 1346.350 75.580 ;
        RECT 531.830 15.540 532.150 15.600 ;
        RECT 537.350 15.540 537.670 15.600 ;
        RECT 531.830 15.400 537.670 15.540 ;
        RECT 531.830 15.340 532.150 15.400 ;
        RECT 537.350 15.340 537.670 15.400 ;
      LAYER via ;
        RECT 1346.060 1677.940 1346.320 1678.200 ;
        RECT 1347.900 1677.940 1348.160 1678.200 ;
        RECT 537.380 75.520 537.640 75.780 ;
        RECT 1346.060 75.520 1346.320 75.780 ;
        RECT 531.860 15.340 532.120 15.600 ;
        RECT 537.380 15.340 537.640 15.600 ;
      LAYER met2 ;
        RECT 1349.665 1700.410 1349.945 1704.000 ;
        RECT 1347.960 1700.270 1349.945 1700.410 ;
        RECT 1347.960 1678.230 1348.100 1700.270 ;
        RECT 1349.665 1700.000 1349.945 1700.270 ;
        RECT 1346.060 1677.910 1346.320 1678.230 ;
        RECT 1347.900 1677.910 1348.160 1678.230 ;
        RECT 1346.120 75.810 1346.260 1677.910 ;
        RECT 537.380 75.490 537.640 75.810 ;
        RECT 1346.060 75.490 1346.320 75.810 ;
        RECT 537.440 15.630 537.580 75.490 ;
        RECT 531.860 15.310 532.120 15.630 ;
        RECT 537.380 15.310 537.640 15.630 ;
        RECT 531.920 2.400 532.060 15.310 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.930 1692.080 1353.250 1692.140 ;
        RECT 1356.150 1692.080 1356.470 1692.140 ;
        RECT 1352.930 1691.940 1356.470 1692.080 ;
        RECT 1352.930 1691.880 1353.250 1691.940 ;
        RECT 1356.150 1691.880 1356.470 1691.940 ;
        RECT 551.610 71.980 551.930 72.040 ;
        RECT 1352.930 71.980 1353.250 72.040 ;
        RECT 551.610 71.840 1353.250 71.980 ;
        RECT 551.610 71.780 551.930 71.840 ;
        RECT 1352.930 71.780 1353.250 71.840 ;
      LAYER via ;
        RECT 1352.960 1691.880 1353.220 1692.140 ;
        RECT 1356.180 1691.880 1356.440 1692.140 ;
        RECT 551.640 71.780 551.900 72.040 ;
        RECT 1352.960 71.780 1353.220 72.040 ;
      LAYER met2 ;
        RECT 1356.105 1700.000 1356.385 1704.000 ;
        RECT 1356.240 1692.170 1356.380 1700.000 ;
        RECT 1352.960 1691.850 1353.220 1692.170 ;
        RECT 1356.180 1691.850 1356.440 1692.170 ;
        RECT 1353.020 72.070 1353.160 1691.850 ;
        RECT 551.640 71.750 551.900 72.070 ;
        RECT 1352.960 71.750 1353.220 72.070 ;
        RECT 551.700 16.730 551.840 71.750 ;
        RECT 549.860 16.590 551.840 16.730 ;
        RECT 549.860 2.400 550.000 16.590 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1359.830 1678.140 1360.150 1678.200 ;
        RECT 1361.670 1678.140 1361.990 1678.200 ;
        RECT 1359.830 1678.000 1361.990 1678.140 ;
        RECT 1359.830 1677.940 1360.150 1678.000 ;
        RECT 1361.670 1677.940 1361.990 1678.000 ;
        RECT 572.310 71.640 572.630 71.700 ;
        RECT 1359.830 71.640 1360.150 71.700 ;
        RECT 572.310 71.500 1360.150 71.640 ;
        RECT 572.310 71.440 572.630 71.500 ;
        RECT 1359.830 71.440 1360.150 71.500 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 1359.860 1677.940 1360.120 1678.200 ;
        RECT 1361.700 1677.940 1361.960 1678.200 ;
        RECT 572.340 71.440 572.600 71.700 ;
        RECT 1359.860 71.440 1360.120 71.700 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1363.005 1700.410 1363.285 1704.000 ;
        RECT 1361.760 1700.270 1363.285 1700.410 ;
        RECT 1361.760 1678.230 1361.900 1700.270 ;
        RECT 1363.005 1700.000 1363.285 1700.270 ;
        RECT 1359.860 1677.910 1360.120 1678.230 ;
        RECT 1361.700 1677.910 1361.960 1678.230 ;
        RECT 1359.920 71.730 1360.060 1677.910 ;
        RECT 572.340 71.410 572.600 71.730 ;
        RECT 1359.860 71.410 1360.120 71.730 ;
        RECT 572.400 14.950 572.540 71.410 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.400 567.940 14.630 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.730 1666.580 1367.050 1666.640 ;
        RECT 1368.110 1666.580 1368.430 1666.640 ;
        RECT 1366.730 1666.440 1368.430 1666.580 ;
        RECT 1366.730 1666.380 1367.050 1666.440 ;
        RECT 1368.110 1666.380 1368.430 1666.440 ;
        RECT 1366.730 1076.340 1367.050 1076.400 ;
        RECT 1367.650 1076.340 1367.970 1076.400 ;
        RECT 1366.730 1076.200 1367.970 1076.340 ;
        RECT 1366.730 1076.140 1367.050 1076.200 ;
        RECT 1367.650 1076.140 1367.970 1076.200 ;
        RECT 1366.730 980.120 1367.050 980.180 ;
        RECT 1367.650 980.120 1367.970 980.180 ;
        RECT 1366.730 979.980 1367.970 980.120 ;
        RECT 1366.730 979.920 1367.050 979.980 ;
        RECT 1367.650 979.920 1367.970 979.980 ;
        RECT 1366.730 303.320 1367.050 303.580 ;
        RECT 1366.820 303.180 1366.960 303.320 ;
        RECT 1367.650 303.180 1367.970 303.240 ;
        RECT 1366.820 303.040 1367.970 303.180 ;
        RECT 1367.650 302.980 1367.970 303.040 ;
        RECT 1366.270 193.360 1366.590 193.420 ;
        RECT 1367.650 193.360 1367.970 193.420 ;
        RECT 1366.270 193.220 1367.970 193.360 ;
        RECT 1366.270 193.160 1366.590 193.220 ;
        RECT 1367.650 193.160 1367.970 193.220 ;
        RECT 586.110 71.300 586.430 71.360 ;
        RECT 1366.730 71.300 1367.050 71.360 ;
        RECT 586.110 71.160 1367.050 71.300 ;
        RECT 586.110 71.100 586.430 71.160 ;
        RECT 1366.730 71.100 1367.050 71.160 ;
      LAYER via ;
        RECT 1366.760 1666.380 1367.020 1666.640 ;
        RECT 1368.140 1666.380 1368.400 1666.640 ;
        RECT 1366.760 1076.140 1367.020 1076.400 ;
        RECT 1367.680 1076.140 1367.940 1076.400 ;
        RECT 1366.760 979.920 1367.020 980.180 ;
        RECT 1367.680 979.920 1367.940 980.180 ;
        RECT 1366.760 303.320 1367.020 303.580 ;
        RECT 1367.680 302.980 1367.940 303.240 ;
        RECT 1366.300 193.160 1366.560 193.420 ;
        RECT 1367.680 193.160 1367.940 193.420 ;
        RECT 586.140 71.100 586.400 71.360 ;
        RECT 1366.760 71.100 1367.020 71.360 ;
      LAYER met2 ;
        RECT 1369.905 1700.410 1370.185 1704.000 ;
        RECT 1368.200 1700.270 1370.185 1700.410 ;
        RECT 1368.200 1666.670 1368.340 1700.270 ;
        RECT 1369.905 1700.000 1370.185 1700.270 ;
        RECT 1366.760 1666.350 1367.020 1666.670 ;
        RECT 1368.140 1666.350 1368.400 1666.670 ;
        RECT 1366.820 1076.430 1366.960 1666.350 ;
        RECT 1366.760 1076.110 1367.020 1076.430 ;
        RECT 1367.680 1076.110 1367.940 1076.430 ;
        RECT 1367.740 980.210 1367.880 1076.110 ;
        RECT 1366.760 979.890 1367.020 980.210 ;
        RECT 1367.680 979.890 1367.940 980.210 ;
        RECT 1366.820 303.610 1366.960 979.890 ;
        RECT 1366.760 303.290 1367.020 303.610 ;
        RECT 1367.680 302.950 1367.940 303.270 ;
        RECT 1367.740 193.450 1367.880 302.950 ;
        RECT 1366.300 193.130 1366.560 193.450 ;
        RECT 1367.680 193.130 1367.940 193.450 ;
        RECT 1366.360 158.170 1366.500 193.130 ;
        RECT 1366.360 158.030 1366.960 158.170 ;
        RECT 1366.820 71.390 1366.960 158.030 ;
        RECT 586.140 71.070 586.400 71.390 ;
        RECT 1366.760 71.070 1367.020 71.390 ;
        RECT 586.200 17.410 586.340 71.070 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1180.430 1678.140 1180.750 1678.200 ;
        RECT 1182.270 1678.140 1182.590 1678.200 ;
        RECT 1180.430 1678.000 1182.590 1678.140 ;
        RECT 1180.430 1677.940 1180.750 1678.000 ;
        RECT 1182.270 1677.940 1182.590 1678.000 ;
        RECT 91.610 58.720 91.930 58.780 ;
        RECT 1180.430 58.720 1180.750 58.780 ;
        RECT 91.610 58.580 1180.750 58.720 ;
        RECT 91.610 58.520 91.930 58.580 ;
        RECT 1180.430 58.520 1180.750 58.580 ;
      LAYER via ;
        RECT 1180.460 1677.940 1180.720 1678.200 ;
        RECT 1182.300 1677.940 1182.560 1678.200 ;
        RECT 91.640 58.520 91.900 58.780 ;
        RECT 1180.460 58.520 1180.720 58.780 ;
      LAYER met2 ;
        RECT 1183.605 1700.410 1183.885 1704.000 ;
        RECT 1182.360 1700.270 1183.885 1700.410 ;
        RECT 1182.360 1678.230 1182.500 1700.270 ;
        RECT 1183.605 1700.000 1183.885 1700.270 ;
        RECT 1180.460 1677.910 1180.720 1678.230 ;
        RECT 1182.300 1677.910 1182.560 1678.230 ;
        RECT 1180.520 58.810 1180.660 1677.910 ;
        RECT 91.640 58.490 91.900 58.810 ;
        RECT 1180.460 58.490 1180.720 58.810 ;
        RECT 91.700 2.400 91.840 58.490 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1373.630 1678.140 1373.950 1678.200 ;
        RECT 1374.550 1678.140 1374.870 1678.200 ;
        RECT 1373.630 1678.000 1374.870 1678.140 ;
        RECT 1373.630 1677.940 1373.950 1678.000 ;
        RECT 1374.550 1677.940 1374.870 1678.000 ;
        RECT 606.810 70.960 607.130 71.020 ;
        RECT 1373.630 70.960 1373.950 71.020 ;
        RECT 606.810 70.820 1373.950 70.960 ;
        RECT 606.810 70.760 607.130 70.820 ;
        RECT 1373.630 70.760 1373.950 70.820 ;
        RECT 603.130 14.860 603.450 14.920 ;
        RECT 606.810 14.860 607.130 14.920 ;
        RECT 603.130 14.720 607.130 14.860 ;
        RECT 603.130 14.660 603.450 14.720 ;
        RECT 606.810 14.660 607.130 14.720 ;
      LAYER via ;
        RECT 1373.660 1677.940 1373.920 1678.200 ;
        RECT 1374.580 1677.940 1374.840 1678.200 ;
        RECT 606.840 70.760 607.100 71.020 ;
        RECT 1373.660 70.760 1373.920 71.020 ;
        RECT 603.160 14.660 603.420 14.920 ;
        RECT 606.840 14.660 607.100 14.920 ;
      LAYER met2 ;
        RECT 1376.345 1700.410 1376.625 1704.000 ;
        RECT 1374.640 1700.270 1376.625 1700.410 ;
        RECT 1374.640 1678.230 1374.780 1700.270 ;
        RECT 1376.345 1700.000 1376.625 1700.270 ;
        RECT 1373.660 1677.910 1373.920 1678.230 ;
        RECT 1374.580 1677.910 1374.840 1678.230 ;
        RECT 1373.720 71.050 1373.860 1677.910 ;
        RECT 606.840 70.730 607.100 71.050 ;
        RECT 1373.660 70.730 1373.920 71.050 ;
        RECT 606.900 14.950 607.040 70.730 ;
        RECT 603.160 14.630 603.420 14.950 ;
        RECT 606.840 14.630 607.100 14.950 ;
        RECT 603.220 2.400 603.360 14.630 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1381.450 932.180 1381.770 932.240 ;
        RECT 1380.620 932.040 1381.770 932.180 ;
        RECT 1380.620 931.900 1380.760 932.040 ;
        RECT 1381.450 931.980 1381.770 932.040 ;
        RECT 1380.530 931.640 1380.850 931.900 ;
        RECT 1380.530 883.020 1380.850 883.280 ;
        RECT 1380.620 882.880 1380.760 883.020 ;
        RECT 1381.450 882.880 1381.770 882.940 ;
        RECT 1380.620 882.740 1381.770 882.880 ;
        RECT 1381.450 882.680 1381.770 882.740 ;
        RECT 1381.450 352.480 1381.770 352.540 ;
        RECT 1380.620 352.340 1381.770 352.480 ;
        RECT 1380.620 352.200 1380.760 352.340 ;
        RECT 1381.450 352.280 1381.770 352.340 ;
        RECT 1380.530 351.940 1380.850 352.200 ;
        RECT 627.050 70.620 627.370 70.680 ;
        RECT 1380.530 70.620 1380.850 70.680 ;
        RECT 627.050 70.480 1380.850 70.620 ;
        RECT 627.050 70.420 627.370 70.480 ;
        RECT 1380.530 70.420 1380.850 70.480 ;
        RECT 621.070 20.980 621.390 21.040 ;
        RECT 627.050 20.980 627.370 21.040 ;
        RECT 621.070 20.840 627.370 20.980 ;
        RECT 621.070 20.780 621.390 20.840 ;
        RECT 627.050 20.780 627.370 20.840 ;
      LAYER via ;
        RECT 1381.480 931.980 1381.740 932.240 ;
        RECT 1380.560 931.640 1380.820 931.900 ;
        RECT 1380.560 883.020 1380.820 883.280 ;
        RECT 1381.480 882.680 1381.740 882.940 ;
        RECT 1381.480 352.280 1381.740 352.540 ;
        RECT 1380.560 351.940 1380.820 352.200 ;
        RECT 627.080 70.420 627.340 70.680 ;
        RECT 1380.560 70.420 1380.820 70.680 ;
        RECT 621.100 20.780 621.360 21.040 ;
        RECT 627.080 20.780 627.340 21.040 ;
      LAYER met2 ;
        RECT 1383.245 1700.410 1383.525 1704.000 ;
        RECT 1381.540 1700.270 1383.525 1700.410 ;
        RECT 1381.540 932.270 1381.680 1700.270 ;
        RECT 1383.245 1700.000 1383.525 1700.270 ;
        RECT 1381.480 931.950 1381.740 932.270 ;
        RECT 1380.560 931.610 1380.820 931.930 ;
        RECT 1380.620 883.310 1380.760 931.610 ;
        RECT 1380.560 882.990 1380.820 883.310 ;
        RECT 1381.480 882.650 1381.740 882.970 ;
        RECT 1381.540 352.570 1381.680 882.650 ;
        RECT 1381.480 352.250 1381.740 352.570 ;
        RECT 1380.560 351.910 1380.820 352.230 ;
        RECT 1380.620 70.710 1380.760 351.910 ;
        RECT 627.080 70.390 627.340 70.710 ;
        RECT 1380.560 70.390 1380.820 70.710 ;
        RECT 627.140 21.070 627.280 70.390 ;
        RECT 621.100 20.750 621.360 21.070 ;
        RECT 627.080 20.750 627.340 21.070 ;
        RECT 621.160 2.400 621.300 20.750 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1187.330 1678.140 1187.650 1678.200 ;
        RECT 1190.550 1678.140 1190.870 1678.200 ;
        RECT 1187.330 1678.000 1190.870 1678.140 ;
        RECT 1187.330 1677.940 1187.650 1678.000 ;
        RECT 1190.550 1677.940 1190.870 1678.000 ;
        RECT 116.910 65.520 117.230 65.580 ;
        RECT 1187.330 65.520 1187.650 65.580 ;
        RECT 116.910 65.380 1187.650 65.520 ;
        RECT 116.910 65.320 117.230 65.380 ;
        RECT 1187.330 65.320 1187.650 65.380 ;
        RECT 115.530 2.960 115.850 3.020 ;
        RECT 116.910 2.960 117.230 3.020 ;
        RECT 115.530 2.820 117.230 2.960 ;
        RECT 115.530 2.760 115.850 2.820 ;
        RECT 116.910 2.760 117.230 2.820 ;
      LAYER via ;
        RECT 1187.360 1677.940 1187.620 1678.200 ;
        RECT 1190.580 1677.940 1190.840 1678.200 ;
        RECT 116.940 65.320 117.200 65.580 ;
        RECT 1187.360 65.320 1187.620 65.580 ;
        RECT 115.560 2.760 115.820 3.020 ;
        RECT 116.940 2.760 117.200 3.020 ;
      LAYER met2 ;
        RECT 1192.345 1700.410 1192.625 1704.000 ;
        RECT 1190.640 1700.270 1192.625 1700.410 ;
        RECT 1190.640 1678.230 1190.780 1700.270 ;
        RECT 1192.345 1700.000 1192.625 1700.270 ;
        RECT 1187.360 1677.910 1187.620 1678.230 ;
        RECT 1190.580 1677.910 1190.840 1678.230 ;
        RECT 1187.420 65.610 1187.560 1677.910 ;
        RECT 116.940 65.290 117.200 65.610 ;
        RECT 1187.360 65.290 1187.620 65.610 ;
        RECT 117.000 3.050 117.140 65.290 ;
        RECT 115.560 2.730 115.820 3.050 ;
        RECT 116.940 2.730 117.200 3.050 ;
        RECT 115.620 2.400 115.760 2.730 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1170.770 1686.980 1171.090 1687.040 ;
        RECT 1201.590 1686.980 1201.910 1687.040 ;
        RECT 1170.770 1686.840 1201.910 1686.980 ;
        RECT 1170.770 1686.780 1171.090 1686.840 ;
        RECT 1201.590 1686.780 1201.910 1686.840 ;
        RECT 139.450 45.120 139.770 45.180 ;
        RECT 1169.390 45.120 1169.710 45.180 ;
        RECT 139.450 44.980 1169.710 45.120 ;
        RECT 139.450 44.920 139.770 44.980 ;
        RECT 1169.390 44.920 1169.710 44.980 ;
      LAYER via ;
        RECT 1170.800 1686.780 1171.060 1687.040 ;
        RECT 1201.620 1686.780 1201.880 1687.040 ;
        RECT 139.480 44.920 139.740 45.180 ;
        RECT 1169.420 44.920 1169.680 45.180 ;
      LAYER met2 ;
        RECT 1201.545 1700.000 1201.825 1704.000 ;
        RECT 1201.680 1687.070 1201.820 1700.000 ;
        RECT 1170.800 1686.750 1171.060 1687.070 ;
        RECT 1201.620 1686.750 1201.880 1687.070 ;
        RECT 1170.860 1671.850 1171.000 1686.750 ;
        RECT 1169.480 1671.710 1171.000 1671.850 ;
        RECT 1169.480 45.210 1169.620 1671.710 ;
        RECT 139.480 44.890 139.740 45.210 ;
        RECT 1169.420 44.890 1169.680 45.210 ;
        RECT 139.540 2.400 139.680 44.890 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 72.320 158.630 72.380 ;
        RECT 1208.490 72.320 1208.810 72.380 ;
        RECT 158.310 72.180 1208.810 72.320 ;
        RECT 158.310 72.120 158.630 72.180 ;
        RECT 1208.490 72.120 1208.810 72.180 ;
      LAYER via ;
        RECT 158.340 72.120 158.600 72.380 ;
        RECT 1208.520 72.120 1208.780 72.380 ;
      LAYER met2 ;
        RECT 1207.985 1700.410 1208.265 1704.000 ;
        RECT 1207.985 1700.270 1208.720 1700.410 ;
        RECT 1207.985 1700.000 1208.265 1700.270 ;
        RECT 1208.580 72.410 1208.720 1700.270 ;
        RECT 158.340 72.090 158.600 72.410 ;
        RECT 1208.520 72.090 1208.780 72.410 ;
        RECT 158.400 3.130 158.540 72.090 ;
        RECT 157.480 2.990 158.540 3.130 ;
        RECT 157.480 2.400 157.620 2.990 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 286.190 1689.020 286.510 1689.080 ;
        RECT 1214.930 1689.020 1215.250 1689.080 ;
        RECT 286.190 1688.880 1215.250 1689.020 ;
        RECT 286.190 1688.820 286.510 1688.880 ;
        RECT 1214.930 1688.820 1215.250 1688.880 ;
        RECT 174.870 16.900 175.190 16.960 ;
        RECT 286.190 16.900 286.510 16.960 ;
        RECT 174.870 16.760 286.510 16.900 ;
        RECT 174.870 16.700 175.190 16.760 ;
        RECT 286.190 16.700 286.510 16.760 ;
      LAYER via ;
        RECT 286.220 1688.820 286.480 1689.080 ;
        RECT 1214.960 1688.820 1215.220 1689.080 ;
        RECT 174.900 16.700 175.160 16.960 ;
        RECT 286.220 16.700 286.480 16.960 ;
      LAYER met2 ;
        RECT 1214.885 1700.000 1215.165 1704.000 ;
        RECT 1215.020 1689.110 1215.160 1700.000 ;
        RECT 286.220 1688.790 286.480 1689.110 ;
        RECT 1214.960 1688.790 1215.220 1689.110 ;
        RECT 286.280 16.990 286.420 1688.790 ;
        RECT 174.900 16.670 175.160 16.990 ;
        RECT 286.220 16.670 286.480 16.990 ;
        RECT 174.960 2.400 175.100 16.670 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.830 1656.180 1222.150 1656.440 ;
        RECT 1221.920 1655.760 1222.060 1656.180 ;
        RECT 1221.830 1655.500 1222.150 1655.760 ;
        RECT 192.810 18.940 193.130 19.000 ;
        RECT 1222.290 18.940 1222.610 19.000 ;
        RECT 192.810 18.800 1222.610 18.940 ;
        RECT 192.810 18.740 193.130 18.800 ;
        RECT 1222.290 18.740 1222.610 18.800 ;
      LAYER via ;
        RECT 1221.860 1656.180 1222.120 1656.440 ;
        RECT 1221.860 1655.500 1222.120 1655.760 ;
        RECT 192.840 18.740 193.100 19.000 ;
        RECT 1222.320 18.740 1222.580 19.000 ;
      LAYER met2 ;
        RECT 1221.785 1700.000 1222.065 1704.000 ;
        RECT 1221.920 1656.470 1222.060 1700.000 ;
        RECT 1221.860 1656.150 1222.120 1656.470 ;
        RECT 1221.860 1655.470 1222.120 1655.790 ;
        RECT 1221.920 26.250 1222.060 1655.470 ;
        RECT 1221.920 26.110 1222.520 26.250 ;
        RECT 1222.380 19.030 1222.520 26.110 ;
        RECT 192.840 18.710 193.100 19.030 ;
        RECT 1222.320 18.710 1222.580 19.030 ;
        RECT 192.900 2.400 193.040 18.710 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 334.490 1689.700 334.810 1689.760 ;
        RECT 1228.270 1689.700 1228.590 1689.760 ;
        RECT 334.490 1689.560 1228.590 1689.700 ;
        RECT 334.490 1689.500 334.810 1689.560 ;
        RECT 1228.270 1689.500 1228.590 1689.560 ;
        RECT 210.750 16.560 211.070 16.620 ;
        RECT 334.490 16.560 334.810 16.620 ;
        RECT 210.750 16.420 334.810 16.560 ;
        RECT 210.750 16.360 211.070 16.420 ;
        RECT 334.490 16.360 334.810 16.420 ;
      LAYER via ;
        RECT 334.520 1689.500 334.780 1689.760 ;
        RECT 1228.300 1689.500 1228.560 1689.760 ;
        RECT 210.780 16.360 211.040 16.620 ;
        RECT 334.520 16.360 334.780 16.620 ;
      LAYER met2 ;
        RECT 1228.225 1700.000 1228.505 1704.000 ;
        RECT 1228.360 1689.790 1228.500 1700.000 ;
        RECT 334.520 1689.470 334.780 1689.790 ;
        RECT 1228.300 1689.470 1228.560 1689.790 ;
        RECT 334.580 16.650 334.720 1689.470 ;
        RECT 210.780 16.330 211.040 16.650 ;
        RECT 334.520 16.330 334.780 16.650 ;
        RECT 210.840 2.400 210.980 16.330 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1231.490 1686.300 1231.810 1686.360 ;
        RECT 1235.170 1686.300 1235.490 1686.360 ;
        RECT 1231.490 1686.160 1235.490 1686.300 ;
        RECT 1231.490 1686.100 1231.810 1686.160 ;
        RECT 1235.170 1686.100 1235.490 1686.160 ;
        RECT 228.690 19.620 229.010 19.680 ;
        RECT 1231.490 19.620 1231.810 19.680 ;
        RECT 228.690 19.480 1231.810 19.620 ;
        RECT 228.690 19.420 229.010 19.480 ;
        RECT 1231.490 19.420 1231.810 19.480 ;
      LAYER via ;
        RECT 1231.520 1686.100 1231.780 1686.360 ;
        RECT 1235.200 1686.100 1235.460 1686.360 ;
        RECT 228.720 19.420 228.980 19.680 ;
        RECT 1231.520 19.420 1231.780 19.680 ;
      LAYER met2 ;
        RECT 1235.125 1700.000 1235.405 1704.000 ;
        RECT 1235.260 1686.390 1235.400 1700.000 ;
        RECT 1231.520 1686.070 1231.780 1686.390 ;
        RECT 1235.200 1686.070 1235.460 1686.390 ;
        RECT 1231.580 19.710 1231.720 1686.070 ;
        RECT 228.720 19.390 228.980 19.710 ;
        RECT 1231.520 19.390 1231.780 19.710 ;
        RECT 228.780 2.400 228.920 19.390 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 65.390 1686.980 65.710 1687.040 ;
        RECT 1168.010 1686.980 1168.330 1687.040 ;
        RECT 65.390 1686.840 1168.330 1686.980 ;
        RECT 65.390 1686.780 65.710 1686.840 ;
        RECT 1168.010 1686.780 1168.330 1686.840 ;
        RECT 50.210 16.560 50.530 16.620 ;
        RECT 65.390 16.560 65.710 16.620 ;
        RECT 50.210 16.420 65.710 16.560 ;
        RECT 50.210 16.360 50.530 16.420 ;
        RECT 65.390 16.360 65.710 16.420 ;
      LAYER via ;
        RECT 65.420 1686.780 65.680 1687.040 ;
        RECT 1168.040 1686.780 1168.300 1687.040 ;
        RECT 50.240 16.360 50.500 16.620 ;
        RECT 65.420 16.360 65.680 16.620 ;
      LAYER met2 ;
        RECT 1167.965 1700.000 1168.245 1704.000 ;
        RECT 1168.100 1687.070 1168.240 1700.000 ;
        RECT 65.420 1686.750 65.680 1687.070 ;
        RECT 1168.040 1686.750 1168.300 1687.070 ;
        RECT 65.480 16.650 65.620 1686.750 ;
        RECT 50.240 16.330 50.500 16.650 ;
        RECT 65.420 16.330 65.680 16.650 ;
        RECT 50.300 2.400 50.440 16.330 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1238.850 1686.300 1239.170 1686.360 ;
        RECT 1243.910 1686.300 1244.230 1686.360 ;
        RECT 1238.850 1686.160 1244.230 1686.300 ;
        RECT 1238.850 1686.100 1239.170 1686.160 ;
        RECT 1243.910 1686.100 1244.230 1686.160 ;
        RECT 252.610 20.300 252.930 20.360 ;
        RECT 1238.390 20.300 1238.710 20.360 ;
        RECT 252.610 20.160 1238.710 20.300 ;
        RECT 252.610 20.100 252.930 20.160 ;
        RECT 1238.390 20.100 1238.710 20.160 ;
      LAYER via ;
        RECT 1238.880 1686.100 1239.140 1686.360 ;
        RECT 1243.940 1686.100 1244.200 1686.360 ;
        RECT 252.640 20.100 252.900 20.360 ;
        RECT 1238.420 20.100 1238.680 20.360 ;
      LAYER met2 ;
        RECT 1243.865 1700.000 1244.145 1704.000 ;
        RECT 1244.000 1686.390 1244.140 1700.000 ;
        RECT 1238.880 1686.070 1239.140 1686.390 ;
        RECT 1243.940 1686.070 1244.200 1686.390 ;
        RECT 1238.940 1677.290 1239.080 1686.070 ;
        RECT 1238.480 1677.150 1239.080 1677.290 ;
        RECT 1238.480 20.390 1238.620 1677.150 ;
        RECT 252.640 20.070 252.900 20.390 ;
        RECT 1238.420 20.070 1238.680 20.390 ;
        RECT 252.700 2.400 252.840 20.070 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 355.190 1690.040 355.510 1690.100 ;
        RECT 1250.810 1690.040 1251.130 1690.100 ;
        RECT 355.190 1689.900 1251.130 1690.040 ;
        RECT 355.190 1689.840 355.510 1689.900 ;
        RECT 1250.810 1689.840 1251.130 1689.900 ;
        RECT 270.090 15.880 270.410 15.940 ;
        RECT 355.190 15.880 355.510 15.940 ;
        RECT 270.090 15.740 355.510 15.880 ;
        RECT 270.090 15.680 270.410 15.740 ;
        RECT 355.190 15.680 355.510 15.740 ;
      LAYER via ;
        RECT 355.220 1689.840 355.480 1690.100 ;
        RECT 1250.840 1689.840 1251.100 1690.100 ;
        RECT 270.120 15.680 270.380 15.940 ;
        RECT 355.220 15.680 355.480 15.940 ;
      LAYER met2 ;
        RECT 1250.765 1700.000 1251.045 1704.000 ;
        RECT 1250.900 1690.130 1251.040 1700.000 ;
        RECT 355.220 1689.810 355.480 1690.130 ;
        RECT 1250.840 1689.810 1251.100 1690.130 ;
        RECT 355.280 15.970 355.420 1689.810 ;
        RECT 270.120 15.650 270.380 15.970 ;
        RECT 355.220 15.650 355.480 15.970 ;
        RECT 270.180 2.400 270.320 15.650 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.290 1686.300 1245.610 1686.360 ;
        RECT 1257.710 1686.300 1258.030 1686.360 ;
        RECT 1245.290 1686.160 1258.030 1686.300 ;
        RECT 1245.290 1686.100 1245.610 1686.160 ;
        RECT 1257.710 1686.100 1258.030 1686.160 ;
        RECT 288.030 20.640 288.350 20.700 ;
        RECT 1245.290 20.640 1245.610 20.700 ;
        RECT 288.030 20.500 1245.610 20.640 ;
        RECT 288.030 20.440 288.350 20.500 ;
        RECT 1245.290 20.440 1245.610 20.500 ;
      LAYER via ;
        RECT 1245.320 1686.100 1245.580 1686.360 ;
        RECT 1257.740 1686.100 1258.000 1686.360 ;
        RECT 288.060 20.440 288.320 20.700 ;
        RECT 1245.320 20.440 1245.580 20.700 ;
      LAYER met2 ;
        RECT 1257.665 1700.000 1257.945 1704.000 ;
        RECT 1257.800 1686.390 1257.940 1700.000 ;
        RECT 1245.320 1686.070 1245.580 1686.390 ;
        RECT 1257.740 1686.070 1258.000 1686.390 ;
        RECT 1245.380 20.730 1245.520 1686.070 ;
        RECT 288.060 20.410 288.320 20.730 ;
        RECT 1245.320 20.410 1245.580 20.730 ;
        RECT 288.120 2.400 288.260 20.410 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1264.150 1686.980 1264.470 1687.040 ;
        RECT 1230.660 1686.840 1264.470 1686.980 ;
        RECT 389.690 1686.300 390.010 1686.360 ;
        RECT 1230.660 1686.300 1230.800 1686.840 ;
        RECT 1264.150 1686.780 1264.470 1686.840 ;
        RECT 389.690 1686.160 1230.800 1686.300 ;
        RECT 389.690 1686.100 390.010 1686.160 ;
        RECT 305.970 15.540 306.290 15.600 ;
        RECT 389.690 15.540 390.010 15.600 ;
        RECT 305.970 15.400 390.010 15.540 ;
        RECT 305.970 15.340 306.290 15.400 ;
        RECT 389.690 15.340 390.010 15.400 ;
      LAYER via ;
        RECT 389.720 1686.100 389.980 1686.360 ;
        RECT 1264.180 1686.780 1264.440 1687.040 ;
        RECT 306.000 15.340 306.260 15.600 ;
        RECT 389.720 15.340 389.980 15.600 ;
      LAYER met2 ;
        RECT 1264.105 1700.000 1264.385 1704.000 ;
        RECT 1264.240 1687.070 1264.380 1700.000 ;
        RECT 1264.180 1686.750 1264.440 1687.070 ;
        RECT 389.720 1686.070 389.980 1686.390 ;
        RECT 389.780 15.630 389.920 1686.070 ;
        RECT 306.000 15.310 306.260 15.630 ;
        RECT 389.720 15.310 389.980 15.630 ;
        RECT 306.060 2.400 306.200 15.310 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1252.190 1689.360 1252.510 1689.420 ;
        RECT 1271.050 1689.360 1271.370 1689.420 ;
        RECT 1252.190 1689.220 1271.370 1689.360 ;
        RECT 1252.190 1689.160 1252.510 1689.220 ;
        RECT 1271.050 1689.160 1271.370 1689.220 ;
        RECT 323.450 16.900 323.770 16.960 ;
        RECT 1252.190 16.900 1252.510 16.960 ;
        RECT 323.450 16.760 1252.510 16.900 ;
        RECT 323.450 16.700 323.770 16.760 ;
        RECT 1252.190 16.700 1252.510 16.760 ;
      LAYER via ;
        RECT 1252.220 1689.160 1252.480 1689.420 ;
        RECT 1271.080 1689.160 1271.340 1689.420 ;
        RECT 323.480 16.700 323.740 16.960 ;
        RECT 1252.220 16.700 1252.480 16.960 ;
      LAYER met2 ;
        RECT 1271.005 1700.000 1271.285 1704.000 ;
        RECT 1271.140 1689.450 1271.280 1700.000 ;
        RECT 1252.220 1689.130 1252.480 1689.450 ;
        RECT 1271.080 1689.130 1271.340 1689.450 ;
        RECT 1252.280 16.990 1252.420 1689.130 ;
        RECT 323.480 16.670 323.740 16.990 ;
        RECT 1252.220 16.670 1252.480 16.990 ;
        RECT 323.540 8.570 323.680 16.670 ;
        RECT 323.540 8.430 324.140 8.570 ;
        RECT 324.000 2.400 324.140 8.430 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 513.890 1684.260 514.210 1684.320 ;
        RECT 1277.950 1684.260 1278.270 1684.320 ;
        RECT 513.890 1684.120 1278.270 1684.260 ;
        RECT 513.890 1684.060 514.210 1684.120 ;
        RECT 1277.950 1684.060 1278.270 1684.120 ;
        RECT 341.390 15.200 341.710 15.260 ;
        RECT 512.970 15.200 513.290 15.260 ;
        RECT 341.390 15.060 513.290 15.200 ;
        RECT 341.390 15.000 341.710 15.060 ;
        RECT 512.970 15.000 513.290 15.060 ;
      LAYER via ;
        RECT 513.920 1684.060 514.180 1684.320 ;
        RECT 1277.980 1684.060 1278.240 1684.320 ;
        RECT 341.420 15.000 341.680 15.260 ;
        RECT 513.000 15.000 513.260 15.260 ;
      LAYER met2 ;
        RECT 1277.905 1700.000 1278.185 1704.000 ;
        RECT 1278.040 1684.350 1278.180 1700.000 ;
        RECT 513.920 1684.030 514.180 1684.350 ;
        RECT 1277.980 1684.030 1278.240 1684.350 ;
        RECT 513.980 16.050 514.120 1684.030 ;
        RECT 513.060 15.910 514.120 16.050 ;
        RECT 513.060 15.290 513.200 15.910 ;
        RECT 341.420 14.970 341.680 15.290 ;
        RECT 513.000 14.970 513.260 15.290 ;
        RECT 341.480 2.400 341.620 14.970 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1259.090 1689.700 1259.410 1689.760 ;
        RECT 1284.390 1689.700 1284.710 1689.760 ;
        RECT 1259.090 1689.560 1284.710 1689.700 ;
        RECT 1259.090 1689.500 1259.410 1689.560 ;
        RECT 1284.390 1689.500 1284.710 1689.560 ;
        RECT 359.330 16.560 359.650 16.620 ;
        RECT 1259.090 16.560 1259.410 16.620 ;
        RECT 359.330 16.420 1259.410 16.560 ;
        RECT 359.330 16.360 359.650 16.420 ;
        RECT 1259.090 16.360 1259.410 16.420 ;
      LAYER via ;
        RECT 1259.120 1689.500 1259.380 1689.760 ;
        RECT 1284.420 1689.500 1284.680 1689.760 ;
        RECT 359.360 16.360 359.620 16.620 ;
        RECT 1259.120 16.360 1259.380 16.620 ;
      LAYER met2 ;
        RECT 1284.345 1700.000 1284.625 1704.000 ;
        RECT 1284.480 1689.790 1284.620 1700.000 ;
        RECT 1259.120 1689.470 1259.380 1689.790 ;
        RECT 1284.420 1689.470 1284.680 1689.790 ;
        RECT 1259.180 16.650 1259.320 1689.470 ;
        RECT 359.360 16.330 359.620 16.650 ;
        RECT 1259.120 16.330 1259.380 16.650 ;
        RECT 359.420 2.400 359.560 16.330 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 396.590 1690.380 396.910 1690.440 ;
        RECT 1291.290 1690.380 1291.610 1690.440 ;
        RECT 396.590 1690.240 1291.610 1690.380 ;
        RECT 396.590 1690.180 396.910 1690.240 ;
        RECT 1291.290 1690.180 1291.610 1690.240 ;
        RECT 377.270 15.880 377.590 15.940 ;
        RECT 396.590 15.880 396.910 15.940 ;
        RECT 377.270 15.740 396.910 15.880 ;
        RECT 377.270 15.680 377.590 15.740 ;
        RECT 396.590 15.680 396.910 15.740 ;
      LAYER via ;
        RECT 396.620 1690.180 396.880 1690.440 ;
        RECT 1291.320 1690.180 1291.580 1690.440 ;
        RECT 377.300 15.680 377.560 15.940 ;
        RECT 396.620 15.680 396.880 15.940 ;
      LAYER met2 ;
        RECT 1291.245 1700.000 1291.525 1704.000 ;
        RECT 1291.380 1690.470 1291.520 1700.000 ;
        RECT 396.620 1690.150 396.880 1690.470 ;
        RECT 1291.320 1690.150 1291.580 1690.470 ;
        RECT 396.680 15.970 396.820 1690.150 ;
        RECT 377.300 15.650 377.560 15.970 ;
        RECT 396.620 15.650 396.880 15.970 ;
        RECT 377.360 2.400 377.500 15.650 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 414.605 14.705 414.775 15.895 ;
      LAYER mcon ;
        RECT 414.605 15.725 414.775 15.895 ;
      LAYER met1 ;
        RECT 1265.990 1686.300 1266.310 1686.360 ;
        RECT 1298.190 1686.300 1298.510 1686.360 ;
        RECT 1265.990 1686.160 1298.510 1686.300 ;
        RECT 1265.990 1686.100 1266.310 1686.160 ;
        RECT 1298.190 1686.100 1298.510 1686.160 ;
        RECT 1265.990 16.220 1266.310 16.280 ;
        RECT 448.660 16.080 1266.310 16.220 ;
        RECT 414.545 15.880 414.835 15.925 ;
        RECT 448.660 15.880 448.800 16.080 ;
        RECT 1265.990 16.020 1266.310 16.080 ;
        RECT 414.545 15.740 448.800 15.880 ;
        RECT 414.545 15.695 414.835 15.740 ;
        RECT 395.210 14.860 395.530 14.920 ;
        RECT 414.545 14.860 414.835 14.905 ;
        RECT 395.210 14.720 414.835 14.860 ;
        RECT 395.210 14.660 395.530 14.720 ;
        RECT 414.545 14.675 414.835 14.720 ;
      LAYER via ;
        RECT 1266.020 1686.100 1266.280 1686.360 ;
        RECT 1298.220 1686.100 1298.480 1686.360 ;
        RECT 1266.020 16.020 1266.280 16.280 ;
        RECT 395.240 14.660 395.500 14.920 ;
      LAYER met2 ;
        RECT 1298.145 1700.000 1298.425 1704.000 ;
        RECT 1298.280 1686.390 1298.420 1700.000 ;
        RECT 1266.020 1686.070 1266.280 1686.390 ;
        RECT 1298.220 1686.070 1298.480 1686.390 ;
        RECT 1266.080 16.310 1266.220 1686.070 ;
        RECT 1266.020 15.990 1266.280 16.310 ;
        RECT 395.240 14.630 395.500 14.950 ;
        RECT 395.300 2.400 395.440 14.630 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1269.285 1687.165 1269.455 1689.035 ;
        RECT 1296.885 1688.525 1297.055 1689.375 ;
        RECT 448.185 1685.465 448.355 1686.655 ;
        RECT 496.945 1684.445 497.115 1686.655 ;
        RECT 544.785 1684.445 544.955 1686.655 ;
        RECT 593.545 1683.765 593.715 1686.655 ;
        RECT 641.385 1683.425 641.555 1686.655 ;
      LAYER mcon ;
        RECT 1296.885 1689.205 1297.055 1689.375 ;
        RECT 1269.285 1688.865 1269.455 1689.035 ;
        RECT 448.185 1686.485 448.355 1686.655 ;
        RECT 496.945 1686.485 497.115 1686.655 ;
        RECT 544.785 1686.485 544.955 1686.655 ;
        RECT 593.545 1686.485 593.715 1686.655 ;
        RECT 641.385 1686.485 641.555 1686.655 ;
      LAYER met1 ;
        RECT 1296.825 1689.360 1297.115 1689.405 ;
        RECT 1271.600 1689.220 1297.115 1689.360 ;
        RECT 1269.225 1689.020 1269.515 1689.065 ;
        RECT 1271.600 1689.020 1271.740 1689.220 ;
        RECT 1296.825 1689.175 1297.115 1689.220 ;
        RECT 1304.630 1689.020 1304.950 1689.080 ;
        RECT 1269.225 1688.880 1271.740 1689.020 ;
        RECT 1297.820 1688.880 1304.950 1689.020 ;
        RECT 1269.225 1688.835 1269.515 1688.880 ;
        RECT 1296.825 1688.680 1297.115 1688.725 ;
        RECT 1297.820 1688.680 1297.960 1688.880 ;
        RECT 1304.630 1688.820 1304.950 1688.880 ;
        RECT 1296.825 1688.540 1297.960 1688.680 ;
        RECT 1296.825 1688.495 1297.115 1688.540 ;
        RECT 1269.225 1687.320 1269.515 1687.365 ;
        RECT 1202.140 1687.180 1269.515 1687.320 ;
        RECT 448.125 1686.640 448.415 1686.685 ;
        RECT 496.885 1686.640 497.175 1686.685 ;
        RECT 448.125 1686.500 497.175 1686.640 ;
        RECT 448.125 1686.455 448.415 1686.500 ;
        RECT 496.885 1686.455 497.175 1686.500 ;
        RECT 544.725 1686.640 545.015 1686.685 ;
        RECT 593.485 1686.640 593.775 1686.685 ;
        RECT 544.725 1686.500 593.775 1686.640 ;
        RECT 544.725 1686.455 545.015 1686.500 ;
        RECT 593.485 1686.455 593.775 1686.500 ;
        RECT 641.325 1686.640 641.615 1686.685 ;
        RECT 690.070 1686.640 690.390 1686.700 ;
        RECT 641.325 1686.500 690.390 1686.640 ;
        RECT 641.325 1686.455 641.615 1686.500 ;
        RECT 690.070 1686.440 690.390 1686.500 ;
        RECT 737.910 1686.640 738.230 1686.700 ;
        RECT 786.670 1686.640 786.990 1686.700 ;
        RECT 737.910 1686.500 786.990 1686.640 ;
        RECT 737.910 1686.440 738.230 1686.500 ;
        RECT 786.670 1686.440 786.990 1686.500 ;
        RECT 834.510 1686.640 834.830 1686.700 ;
        RECT 883.270 1686.640 883.590 1686.700 ;
        RECT 834.510 1686.500 883.590 1686.640 ;
        RECT 834.510 1686.440 834.830 1686.500 ;
        RECT 883.270 1686.440 883.590 1686.500 ;
        RECT 931.110 1686.640 931.430 1686.700 ;
        RECT 979.870 1686.640 980.190 1686.700 ;
        RECT 931.110 1686.500 980.190 1686.640 ;
        RECT 931.110 1686.440 931.430 1686.500 ;
        RECT 979.870 1686.440 980.190 1686.500 ;
        RECT 1027.710 1686.640 1028.030 1686.700 ;
        RECT 1076.470 1686.640 1076.790 1686.700 ;
        RECT 1027.710 1686.500 1076.790 1686.640 ;
        RECT 1027.710 1686.440 1028.030 1686.500 ;
        RECT 1076.470 1686.440 1076.790 1686.500 ;
        RECT 1124.310 1686.640 1124.630 1686.700 ;
        RECT 1202.140 1686.640 1202.280 1687.180 ;
        RECT 1269.225 1687.135 1269.515 1687.180 ;
        RECT 1124.310 1686.500 1202.280 1686.640 ;
        RECT 1124.310 1686.440 1124.630 1686.500 ;
        RECT 424.190 1685.620 424.510 1685.680 ;
        RECT 448.125 1685.620 448.415 1685.665 ;
        RECT 424.190 1685.480 448.415 1685.620 ;
        RECT 424.190 1685.420 424.510 1685.480 ;
        RECT 448.125 1685.435 448.415 1685.480 ;
        RECT 496.885 1684.600 497.175 1684.645 ;
        RECT 544.725 1684.600 545.015 1684.645 ;
        RECT 496.885 1684.460 545.015 1684.600 ;
        RECT 496.885 1684.415 497.175 1684.460 ;
        RECT 544.725 1684.415 545.015 1684.460 ;
        RECT 593.485 1683.920 593.775 1683.965 ;
        RECT 593.485 1683.780 627.280 1683.920 ;
        RECT 593.485 1683.735 593.775 1683.780 ;
        RECT 627.140 1683.580 627.280 1683.780 ;
        RECT 641.325 1683.580 641.615 1683.625 ;
        RECT 627.140 1683.440 641.615 1683.580 ;
        RECT 641.325 1683.395 641.615 1683.440 ;
        RECT 424.190 16.220 424.510 16.280 ;
        RECT 414.160 16.080 424.510 16.220 ;
        RECT 413.150 15.880 413.470 15.940 ;
        RECT 414.160 15.880 414.300 16.080 ;
        RECT 424.190 16.020 424.510 16.080 ;
        RECT 413.150 15.740 414.300 15.880 ;
        RECT 413.150 15.680 413.470 15.740 ;
      LAYER via ;
        RECT 1304.660 1688.820 1304.920 1689.080 ;
        RECT 690.100 1686.440 690.360 1686.700 ;
        RECT 737.940 1686.440 738.200 1686.700 ;
        RECT 786.700 1686.440 786.960 1686.700 ;
        RECT 834.540 1686.440 834.800 1686.700 ;
        RECT 883.300 1686.440 883.560 1686.700 ;
        RECT 931.140 1686.440 931.400 1686.700 ;
        RECT 979.900 1686.440 980.160 1686.700 ;
        RECT 1027.740 1686.440 1028.000 1686.700 ;
        RECT 1076.500 1686.440 1076.760 1686.700 ;
        RECT 1124.340 1686.440 1124.600 1686.700 ;
        RECT 424.220 1685.420 424.480 1685.680 ;
        RECT 413.180 15.680 413.440 15.940 ;
        RECT 424.220 16.020 424.480 16.280 ;
      LAYER met2 ;
        RECT 1304.585 1700.000 1304.865 1704.000 ;
        RECT 1304.720 1689.110 1304.860 1700.000 ;
        RECT 1304.660 1688.790 1304.920 1689.110 ;
        RECT 690.100 1686.410 690.360 1686.730 ;
        RECT 737.940 1686.410 738.200 1686.730 ;
        RECT 786.700 1686.410 786.960 1686.730 ;
        RECT 834.540 1686.410 834.800 1686.730 ;
        RECT 883.300 1686.410 883.560 1686.730 ;
        RECT 931.140 1686.410 931.400 1686.730 ;
        RECT 979.900 1686.410 980.160 1686.730 ;
        RECT 1027.740 1686.410 1028.000 1686.730 ;
        RECT 1076.500 1686.410 1076.760 1686.730 ;
        RECT 1124.340 1686.410 1124.600 1686.730 ;
        RECT 690.160 1686.245 690.300 1686.410 ;
        RECT 738.000 1686.245 738.140 1686.410 ;
        RECT 786.760 1686.245 786.900 1686.410 ;
        RECT 834.600 1686.245 834.740 1686.410 ;
        RECT 883.360 1686.245 883.500 1686.410 ;
        RECT 931.200 1686.245 931.340 1686.410 ;
        RECT 979.960 1686.245 980.100 1686.410 ;
        RECT 1027.800 1686.245 1027.940 1686.410 ;
        RECT 1076.560 1686.245 1076.700 1686.410 ;
        RECT 1124.400 1686.245 1124.540 1686.410 ;
        RECT 690.090 1685.875 690.370 1686.245 ;
        RECT 737.930 1685.875 738.210 1686.245 ;
        RECT 786.690 1685.875 786.970 1686.245 ;
        RECT 834.530 1685.875 834.810 1686.245 ;
        RECT 883.290 1685.875 883.570 1686.245 ;
        RECT 931.130 1685.875 931.410 1686.245 ;
        RECT 979.890 1685.875 980.170 1686.245 ;
        RECT 1027.730 1685.875 1028.010 1686.245 ;
        RECT 1076.490 1685.875 1076.770 1686.245 ;
        RECT 1124.330 1685.875 1124.610 1686.245 ;
        RECT 424.220 1685.390 424.480 1685.710 ;
        RECT 424.280 16.310 424.420 1685.390 ;
        RECT 424.220 15.990 424.480 16.310 ;
        RECT 413.180 15.650 413.440 15.970 ;
        RECT 413.240 2.400 413.380 15.650 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 690.090 1685.920 690.370 1686.200 ;
        RECT 737.930 1685.920 738.210 1686.200 ;
        RECT 786.690 1685.920 786.970 1686.200 ;
        RECT 834.530 1685.920 834.810 1686.200 ;
        RECT 883.290 1685.920 883.570 1686.200 ;
        RECT 931.130 1685.920 931.410 1686.200 ;
        RECT 979.890 1685.920 980.170 1686.200 ;
        RECT 1027.730 1685.920 1028.010 1686.200 ;
        RECT 1076.490 1685.920 1076.770 1686.200 ;
        RECT 1124.330 1685.920 1124.610 1686.200 ;
      LAYER met3 ;
        RECT 690.065 1686.210 690.395 1686.225 ;
        RECT 737.905 1686.210 738.235 1686.225 ;
        RECT 690.065 1685.910 738.235 1686.210 ;
        RECT 690.065 1685.895 690.395 1685.910 ;
        RECT 737.905 1685.895 738.235 1685.910 ;
        RECT 786.665 1686.210 786.995 1686.225 ;
        RECT 834.505 1686.210 834.835 1686.225 ;
        RECT 786.665 1685.910 834.835 1686.210 ;
        RECT 786.665 1685.895 786.995 1685.910 ;
        RECT 834.505 1685.895 834.835 1685.910 ;
        RECT 883.265 1686.210 883.595 1686.225 ;
        RECT 931.105 1686.210 931.435 1686.225 ;
        RECT 883.265 1685.910 931.435 1686.210 ;
        RECT 883.265 1685.895 883.595 1685.910 ;
        RECT 931.105 1685.895 931.435 1685.910 ;
        RECT 979.865 1686.210 980.195 1686.225 ;
        RECT 1027.705 1686.210 1028.035 1686.225 ;
        RECT 979.865 1685.910 1028.035 1686.210 ;
        RECT 979.865 1685.895 980.195 1685.910 ;
        RECT 1027.705 1685.895 1028.035 1685.910 ;
        RECT 1076.465 1686.210 1076.795 1686.225 ;
        RECT 1124.305 1686.210 1124.635 1686.225 ;
        RECT 1076.465 1685.910 1124.635 1686.210 ;
        RECT 1076.465 1685.895 1076.795 1685.910 ;
        RECT 1124.305 1685.895 1124.635 1685.910 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1173.605 55.845 1173.775 62.475 ;
      LAYER mcon ;
        RECT 1173.605 62.305 1173.775 62.475 ;
      LAYER met1 ;
        RECT 1173.530 1678.140 1173.850 1678.200 ;
        RECT 1174.910 1678.140 1175.230 1678.200 ;
        RECT 1173.530 1678.000 1175.230 1678.140 ;
        RECT 1173.530 1677.940 1173.850 1678.000 ;
        RECT 1174.910 1677.940 1175.230 1678.000 ;
        RECT 1173.530 62.460 1173.850 62.520 ;
        RECT 1173.335 62.320 1173.850 62.460 ;
        RECT 1173.530 62.260 1173.850 62.320 ;
        RECT 1173.530 56.000 1173.850 56.060 ;
        RECT 1173.335 55.860 1173.850 56.000 ;
        RECT 1173.530 55.800 1173.850 55.860 ;
        RECT 74.130 17.240 74.450 17.300 ;
        RECT 1173.530 17.240 1173.850 17.300 ;
        RECT 74.130 17.100 1173.850 17.240 ;
        RECT 74.130 17.040 74.450 17.100 ;
        RECT 1173.530 17.040 1173.850 17.100 ;
      LAYER via ;
        RECT 1173.560 1677.940 1173.820 1678.200 ;
        RECT 1174.940 1677.940 1175.200 1678.200 ;
        RECT 1173.560 62.260 1173.820 62.520 ;
        RECT 1173.560 55.800 1173.820 56.060 ;
        RECT 74.160 17.040 74.420 17.300 ;
        RECT 1173.560 17.040 1173.820 17.300 ;
      LAYER met2 ;
        RECT 1176.705 1700.410 1176.985 1704.000 ;
        RECT 1175.000 1700.270 1176.985 1700.410 ;
        RECT 1175.000 1678.230 1175.140 1700.270 ;
        RECT 1176.705 1700.000 1176.985 1700.270 ;
        RECT 1173.560 1677.910 1173.820 1678.230 ;
        RECT 1174.940 1677.910 1175.200 1678.230 ;
        RECT 1173.620 62.550 1173.760 1677.910 ;
        RECT 1173.560 62.230 1173.820 62.550 ;
        RECT 1173.560 55.770 1173.820 56.090 ;
        RECT 1173.620 17.330 1173.760 55.770 ;
        RECT 74.160 17.010 74.420 17.330 ;
        RECT 1173.560 17.010 1173.820 17.330 ;
        RECT 74.220 2.400 74.360 17.010 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 527.690 1684.940 528.010 1685.000 ;
        RECT 1311.530 1684.940 1311.850 1685.000 ;
        RECT 527.690 1684.800 1311.850 1684.940 ;
        RECT 527.690 1684.740 528.010 1684.800 ;
        RECT 1311.530 1684.740 1311.850 1684.800 ;
        RECT 430.630 14.860 430.950 14.920 ;
        RECT 430.630 14.720 487.440 14.860 ;
        RECT 430.630 14.660 430.950 14.720 ;
        RECT 487.300 14.180 487.440 14.720 ;
        RECT 527.690 14.180 528.010 14.240 ;
        RECT 487.300 14.040 528.010 14.180 ;
        RECT 527.690 13.980 528.010 14.040 ;
      LAYER via ;
        RECT 527.720 1684.740 527.980 1685.000 ;
        RECT 1311.560 1684.740 1311.820 1685.000 ;
        RECT 430.660 14.660 430.920 14.920 ;
        RECT 527.720 13.980 527.980 14.240 ;
      LAYER met2 ;
        RECT 1311.485 1700.000 1311.765 1704.000 ;
        RECT 1311.620 1685.030 1311.760 1700.000 ;
        RECT 527.720 1684.710 527.980 1685.030 ;
        RECT 1311.560 1684.710 1311.820 1685.030 ;
        RECT 430.660 14.630 430.920 14.950 ;
        RECT 430.720 2.400 430.860 14.630 ;
        RECT 527.780 14.270 527.920 1684.710 ;
        RECT 527.720 13.950 527.980 14.270 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1297.345 1688.865 1297.515 1690.055 ;
      LAYER mcon ;
        RECT 1297.345 1689.885 1297.515 1690.055 ;
      LAYER met1 ;
        RECT 1297.285 1690.040 1297.575 1690.085 ;
        RECT 1317.970 1690.040 1318.290 1690.100 ;
        RECT 1297.285 1689.900 1318.290 1690.040 ;
        RECT 1297.285 1689.855 1297.575 1689.900 ;
        RECT 1317.970 1689.840 1318.290 1689.900 ;
        RECT 1272.890 1689.020 1273.210 1689.080 ;
        RECT 1297.285 1689.020 1297.575 1689.065 ;
        RECT 1272.890 1688.880 1297.575 1689.020 ;
        RECT 1272.890 1688.820 1273.210 1688.880 ;
        RECT 1297.285 1688.835 1297.575 1688.880 ;
        RECT 1272.890 15.880 1273.210 15.940 ;
        RECT 469.360 15.740 1273.210 15.880 ;
        RECT 448.570 15.540 448.890 15.600 ;
        RECT 469.360 15.540 469.500 15.740 ;
        RECT 1272.890 15.680 1273.210 15.740 ;
        RECT 448.570 15.400 469.500 15.540 ;
        RECT 448.570 15.340 448.890 15.400 ;
      LAYER via ;
        RECT 1318.000 1689.840 1318.260 1690.100 ;
        RECT 1272.920 1688.820 1273.180 1689.080 ;
        RECT 448.600 15.340 448.860 15.600 ;
        RECT 1272.920 15.680 1273.180 15.940 ;
      LAYER met2 ;
        RECT 1317.925 1700.000 1318.205 1704.000 ;
        RECT 1318.060 1690.130 1318.200 1700.000 ;
        RECT 1318.000 1689.810 1318.260 1690.130 ;
        RECT 1272.920 1688.790 1273.180 1689.110 ;
        RECT 1272.980 15.970 1273.120 1688.790 ;
        RECT 1272.920 15.650 1273.180 15.970 ;
        RECT 448.600 15.310 448.860 15.630 ;
        RECT 448.660 2.400 448.800 15.310 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 486.290 1685.960 486.610 1686.020 ;
        RECT 1324.870 1685.960 1325.190 1686.020 ;
        RECT 486.290 1685.820 1325.190 1685.960 ;
        RECT 486.290 1685.760 486.610 1685.820 ;
        RECT 1324.870 1685.760 1325.190 1685.820 ;
        RECT 466.510 14.520 466.830 14.580 ;
        RECT 486.290 14.520 486.610 14.580 ;
        RECT 466.510 14.380 486.610 14.520 ;
        RECT 466.510 14.320 466.830 14.380 ;
        RECT 486.290 14.320 486.610 14.380 ;
      LAYER via ;
        RECT 486.320 1685.760 486.580 1686.020 ;
        RECT 1324.900 1685.760 1325.160 1686.020 ;
        RECT 466.540 14.320 466.800 14.580 ;
        RECT 486.320 14.320 486.580 14.580 ;
      LAYER met2 ;
        RECT 1324.825 1700.000 1325.105 1704.000 ;
        RECT 1324.960 1686.050 1325.100 1700.000 ;
        RECT 486.320 1685.730 486.580 1686.050 ;
        RECT 1324.900 1685.730 1325.160 1686.050 ;
        RECT 486.380 14.610 486.520 1685.730 ;
        RECT 466.540 14.290 466.800 14.610 ;
        RECT 486.320 14.290 486.580 14.610 ;
        RECT 466.600 2.400 466.740 14.290 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 513.965 13.685 514.135 14.875 ;
      LAYER mcon ;
        RECT 513.965 14.705 514.135 14.875 ;
      LAYER met1 ;
        RECT 1297.730 1689.700 1298.050 1689.760 ;
        RECT 1331.770 1689.700 1332.090 1689.760 ;
        RECT 1297.730 1689.560 1332.090 1689.700 ;
        RECT 1297.730 1689.500 1298.050 1689.560 ;
        RECT 1331.770 1689.500 1332.090 1689.560 ;
        RECT 1274.270 1688.340 1274.590 1688.400 ;
        RECT 1297.270 1688.340 1297.590 1688.400 ;
        RECT 1274.270 1688.200 1297.590 1688.340 ;
        RECT 1274.270 1688.140 1274.590 1688.200 ;
        RECT 1297.270 1688.140 1297.590 1688.200 ;
        RECT 1273.350 15.540 1273.670 15.600 ;
        RECT 541.580 15.400 1273.670 15.540 ;
        RECT 513.905 14.860 514.195 14.905 ;
        RECT 541.580 14.860 541.720 15.400 ;
        RECT 1273.350 15.340 1273.670 15.400 ;
        RECT 513.905 14.720 541.720 14.860 ;
        RECT 513.905 14.675 514.195 14.720 ;
        RECT 484.450 14.180 484.770 14.240 ;
        RECT 484.450 14.040 486.980 14.180 ;
        RECT 484.450 13.980 484.770 14.040 ;
        RECT 486.840 13.840 486.980 14.040 ;
        RECT 513.905 13.840 514.195 13.885 ;
        RECT 486.840 13.700 514.195 13.840 ;
        RECT 513.905 13.655 514.195 13.700 ;
      LAYER via ;
        RECT 1297.760 1689.500 1298.020 1689.760 ;
        RECT 1331.800 1689.500 1332.060 1689.760 ;
        RECT 1274.300 1688.140 1274.560 1688.400 ;
        RECT 1297.300 1688.140 1297.560 1688.400 ;
        RECT 1273.380 15.340 1273.640 15.600 ;
        RECT 484.480 13.980 484.740 14.240 ;
      LAYER met2 ;
        RECT 1331.725 1700.000 1332.005 1704.000 ;
        RECT 1331.860 1689.790 1332.000 1700.000 ;
        RECT 1297.760 1689.470 1298.020 1689.790 ;
        RECT 1331.800 1689.470 1332.060 1689.790 ;
        RECT 1274.300 1688.110 1274.560 1688.430 ;
        RECT 1297.300 1688.340 1297.560 1688.430 ;
        RECT 1297.820 1688.340 1297.960 1689.470 ;
        RECT 1297.300 1688.200 1297.960 1688.340 ;
        RECT 1297.300 1688.110 1297.560 1688.200 ;
        RECT 1274.360 1672.530 1274.500 1688.110 ;
        RECT 1273.440 1672.390 1274.500 1672.530 ;
        RECT 1273.440 15.630 1273.580 1672.390 ;
        RECT 1273.380 15.310 1273.640 15.630 ;
        RECT 484.480 13.950 484.740 14.270 ;
        RECT 484.540 2.400 484.680 13.950 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 1685.620 503.630 1685.680 ;
        RECT 1338.210 1685.620 1338.530 1685.680 ;
        RECT 503.310 1685.480 1338.530 1685.620 ;
        RECT 503.310 1685.420 503.630 1685.480 ;
        RECT 1338.210 1685.420 1338.530 1685.480 ;
      LAYER via ;
        RECT 503.340 1685.420 503.600 1685.680 ;
        RECT 1338.240 1685.420 1338.500 1685.680 ;
      LAYER met2 ;
        RECT 1338.165 1700.000 1338.445 1704.000 ;
        RECT 1338.300 1685.710 1338.440 1700.000 ;
        RECT 503.340 1685.390 503.600 1685.710 ;
        RECT 1338.240 1685.390 1338.500 1685.710 ;
        RECT 503.400 16.730 503.540 1685.390 ;
        RECT 502.480 16.590 503.540 16.730 ;
        RECT 502.480 2.400 502.620 16.590 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1343.270 1686.980 1343.590 1687.040 ;
        RECT 1305.180 1686.840 1343.590 1686.980 ;
        RECT 1279.790 1686.640 1280.110 1686.700 ;
        RECT 1305.180 1686.640 1305.320 1686.840 ;
        RECT 1343.270 1686.780 1343.590 1686.840 ;
        RECT 1279.790 1686.500 1305.320 1686.640 ;
        RECT 1279.790 1686.440 1280.110 1686.500 ;
        RECT 1279.790 15.200 1280.110 15.260 ;
        RECT 542.040 15.060 1280.110 15.200 ;
        RECT 519.870 14.520 520.190 14.580 ;
        RECT 542.040 14.520 542.180 15.060 ;
        RECT 1279.790 15.000 1280.110 15.060 ;
        RECT 519.870 14.380 542.180 14.520 ;
        RECT 519.870 14.320 520.190 14.380 ;
      LAYER via ;
        RECT 1279.820 1686.440 1280.080 1686.700 ;
        RECT 1343.300 1686.780 1343.560 1687.040 ;
        RECT 519.900 14.320 520.160 14.580 ;
        RECT 1279.820 15.000 1280.080 15.260 ;
      LAYER met2 ;
        RECT 1345.065 1700.410 1345.345 1704.000 ;
        RECT 1343.360 1700.270 1345.345 1700.410 ;
        RECT 1343.360 1687.070 1343.500 1700.270 ;
        RECT 1345.065 1700.000 1345.345 1700.270 ;
        RECT 1343.300 1686.750 1343.560 1687.070 ;
        RECT 1279.820 1686.410 1280.080 1686.730 ;
        RECT 1279.880 15.290 1280.020 1686.410 ;
        RECT 1279.820 14.970 1280.080 15.290 ;
        RECT 519.900 14.290 520.160 14.610 ;
        RECT 519.960 2.400 520.100 14.290 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 1685.280 538.130 1685.340 ;
        RECT 1352.010 1685.280 1352.330 1685.340 ;
        RECT 537.810 1685.140 1352.330 1685.280 ;
        RECT 537.810 1685.080 538.130 1685.140 ;
        RECT 1352.010 1685.080 1352.330 1685.140 ;
      LAYER via ;
        RECT 537.840 1685.080 538.100 1685.340 ;
        RECT 1352.040 1685.080 1352.300 1685.340 ;
      LAYER met2 ;
        RECT 1351.965 1700.000 1352.245 1704.000 ;
        RECT 1352.100 1685.370 1352.240 1700.000 ;
        RECT 537.840 1685.050 538.100 1685.370 ;
        RECT 1352.040 1685.050 1352.300 1685.370 ;
        RECT 537.900 2.400 538.040 1685.050 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1286.690 1687.320 1287.010 1687.380 ;
        RECT 1358.450 1687.320 1358.770 1687.380 ;
        RECT 1286.690 1687.180 1358.770 1687.320 ;
        RECT 1286.690 1687.120 1287.010 1687.180 ;
        RECT 1358.450 1687.120 1358.770 1687.180 ;
        RECT 1286.690 14.860 1287.010 14.920 ;
        RECT 607.360 14.720 1287.010 14.860 ;
        RECT 555.750 14.520 556.070 14.580 ;
        RECT 607.360 14.520 607.500 14.720 ;
        RECT 1286.690 14.660 1287.010 14.720 ;
        RECT 555.750 14.380 607.500 14.520 ;
        RECT 555.750 14.320 556.070 14.380 ;
      LAYER via ;
        RECT 1286.720 1687.120 1286.980 1687.380 ;
        RECT 1358.480 1687.120 1358.740 1687.380 ;
        RECT 555.780 14.320 556.040 14.580 ;
        RECT 1286.720 14.660 1286.980 14.920 ;
      LAYER met2 ;
        RECT 1358.405 1700.000 1358.685 1704.000 ;
        RECT 1358.540 1687.410 1358.680 1700.000 ;
        RECT 1286.720 1687.090 1286.980 1687.410 ;
        RECT 1358.480 1687.090 1358.740 1687.410 ;
        RECT 1286.780 14.950 1286.920 1687.090 ;
        RECT 1286.720 14.630 1286.980 14.950 ;
        RECT 555.780 14.290 556.040 14.610 ;
        RECT 555.840 2.400 555.980 14.290 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1293.590 1687.660 1293.910 1687.720 ;
        RECT 1365.350 1687.660 1365.670 1687.720 ;
        RECT 1293.590 1687.520 1365.670 1687.660 ;
        RECT 1293.590 1687.460 1293.910 1687.520 ;
        RECT 1365.350 1687.460 1365.670 1687.520 ;
        RECT 1293.590 14.520 1293.910 14.580 ;
        RECT 607.820 14.380 1293.910 14.520 ;
        RECT 573.690 14.180 574.010 14.240 ;
        RECT 607.820 14.180 607.960 14.380 ;
        RECT 1293.590 14.320 1293.910 14.380 ;
        RECT 573.690 14.040 607.960 14.180 ;
        RECT 573.690 13.980 574.010 14.040 ;
      LAYER via ;
        RECT 1293.620 1687.460 1293.880 1687.720 ;
        RECT 1365.380 1687.460 1365.640 1687.720 ;
        RECT 573.720 13.980 573.980 14.240 ;
        RECT 1293.620 14.320 1293.880 14.580 ;
      LAYER met2 ;
        RECT 1365.305 1700.000 1365.585 1704.000 ;
        RECT 1365.440 1687.750 1365.580 1700.000 ;
        RECT 1293.620 1687.430 1293.880 1687.750 ;
        RECT 1365.380 1687.430 1365.640 1687.750 ;
        RECT 1293.680 14.610 1293.820 1687.430 ;
        RECT 1293.620 14.290 1293.880 14.610 ;
        RECT 573.720 13.950 573.980 14.270 ;
        RECT 573.780 2.400 573.920 13.950 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 1684.600 593.330 1684.660 ;
        RECT 1372.250 1684.600 1372.570 1684.660 ;
        RECT 593.010 1684.460 1372.570 1684.600 ;
        RECT 593.010 1684.400 593.330 1684.460 ;
        RECT 1372.250 1684.400 1372.570 1684.460 ;
      LAYER via ;
        RECT 593.040 1684.400 593.300 1684.660 ;
        RECT 1372.280 1684.400 1372.540 1684.660 ;
      LAYER met2 ;
        RECT 1372.205 1700.000 1372.485 1704.000 ;
        RECT 1372.340 1684.690 1372.480 1700.000 ;
        RECT 593.040 1684.370 593.300 1684.690 ;
        RECT 1372.280 1684.370 1372.540 1684.690 ;
        RECT 593.100 16.730 593.240 1684.370 ;
        RECT 591.260 16.590 593.240 16.730 ;
        RECT 591.260 2.400 591.400 16.590 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 141.290 1687.660 141.610 1687.720 ;
        RECT 141.290 1687.520 1148.920 1687.660 ;
        RECT 141.290 1687.460 141.610 1687.520 ;
        RECT 1148.780 1687.320 1148.920 1687.520 ;
        RECT 1185.950 1687.320 1186.270 1687.380 ;
        RECT 1148.780 1687.180 1186.270 1687.320 ;
        RECT 1185.950 1687.120 1186.270 1687.180 ;
        RECT 97.590 16.900 97.910 16.960 ;
        RECT 141.290 16.900 141.610 16.960 ;
        RECT 97.590 16.760 141.610 16.900 ;
        RECT 97.590 16.700 97.910 16.760 ;
        RECT 141.290 16.700 141.610 16.760 ;
      LAYER via ;
        RECT 141.320 1687.460 141.580 1687.720 ;
        RECT 1185.980 1687.120 1186.240 1687.380 ;
        RECT 97.620 16.700 97.880 16.960 ;
        RECT 141.320 16.700 141.580 16.960 ;
      LAYER met2 ;
        RECT 1185.905 1700.000 1186.185 1704.000 ;
        RECT 141.320 1687.430 141.580 1687.750 ;
        RECT 141.380 16.990 141.520 1687.430 ;
        RECT 1186.040 1687.410 1186.180 1700.000 ;
        RECT 1185.980 1687.090 1186.240 1687.410 ;
        RECT 97.620 16.670 97.880 16.990 ;
        RECT 141.320 16.670 141.580 16.990 ;
        RECT 97.680 2.400 97.820 16.670 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1297.805 1687.845 1298.895 1688.015 ;
      LAYER mcon ;
        RECT 1298.725 1687.845 1298.895 1688.015 ;
      LAYER met1 ;
        RECT 1294.050 1688.000 1294.370 1688.060 ;
        RECT 1297.745 1688.000 1298.035 1688.045 ;
        RECT 1294.050 1687.860 1298.035 1688.000 ;
        RECT 1294.050 1687.800 1294.370 1687.860 ;
        RECT 1297.745 1687.815 1298.035 1687.860 ;
        RECT 1298.665 1688.000 1298.955 1688.045 ;
        RECT 1378.690 1688.000 1379.010 1688.060 ;
        RECT 1298.665 1687.860 1379.010 1688.000 ;
        RECT 1298.665 1687.815 1298.955 1687.860 ;
        RECT 1378.690 1687.800 1379.010 1687.860 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 1294.050 14.180 1294.370 14.240 ;
        RECT 609.110 14.040 1294.370 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 1294.050 13.980 1294.370 14.040 ;
      LAYER via ;
        RECT 1294.080 1687.800 1294.340 1688.060 ;
        RECT 1378.720 1687.800 1378.980 1688.060 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 1294.080 13.980 1294.340 14.240 ;
      LAYER met2 ;
        RECT 1378.645 1700.000 1378.925 1704.000 ;
        RECT 1378.780 1688.090 1378.920 1700.000 ;
        RECT 1294.080 1687.770 1294.340 1688.090 ;
        RECT 1378.720 1687.770 1378.980 1688.090 ;
        RECT 1294.140 14.270 1294.280 1687.770 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 1294.080 13.950 1294.340 14.270 ;
        RECT 609.200 2.400 609.340 13.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 1683.920 627.830 1683.980 ;
        RECT 1385.590 1683.920 1385.910 1683.980 ;
        RECT 627.510 1683.780 1385.910 1683.920 ;
        RECT 627.510 1683.720 627.830 1683.780 ;
        RECT 1385.590 1683.720 1385.910 1683.780 ;
      LAYER via ;
        RECT 627.540 1683.720 627.800 1683.980 ;
        RECT 1385.620 1683.720 1385.880 1683.980 ;
      LAYER met2 ;
        RECT 1385.545 1700.000 1385.825 1704.000 ;
        RECT 1385.680 1684.010 1385.820 1700.000 ;
        RECT 627.540 1683.690 627.800 1684.010 ;
        RECT 1385.620 1683.690 1385.880 1684.010 ;
        RECT 627.600 17.410 627.740 1683.690 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1194.305 990.165 1194.475 992.375 ;
        RECT 1194.305 796.705 1194.475 798.575 ;
      LAYER mcon ;
        RECT 1194.305 992.205 1194.475 992.375 ;
        RECT 1194.305 798.405 1194.475 798.575 ;
      LAYER met1 ;
        RECT 1194.230 1548.740 1194.550 1549.000 ;
        RECT 1194.320 1548.320 1194.460 1548.740 ;
        RECT 1194.230 1548.060 1194.550 1548.320 ;
        RECT 1194.230 992.360 1194.550 992.420 ;
        RECT 1194.035 992.220 1194.550 992.360 ;
        RECT 1194.230 992.160 1194.550 992.220 ;
        RECT 1194.230 990.320 1194.550 990.380 ;
        RECT 1194.035 990.180 1194.550 990.320 ;
        RECT 1194.230 990.120 1194.550 990.180 ;
        RECT 1194.230 798.560 1194.550 798.620 ;
        RECT 1194.035 798.420 1194.550 798.560 ;
        RECT 1194.230 798.360 1194.550 798.420 ;
        RECT 1194.230 796.860 1194.550 796.920 ;
        RECT 1194.035 796.720 1194.550 796.860 ;
        RECT 1194.230 796.660 1194.550 796.720 ;
        RECT 1194.230 738.520 1194.550 738.780 ;
        RECT 1194.320 738.100 1194.460 738.520 ;
        RECT 1194.230 737.840 1194.550 738.100 ;
        RECT 121.510 17.920 121.830 17.980 ;
        RECT 1194.230 17.920 1194.550 17.980 ;
        RECT 121.510 17.780 1194.550 17.920 ;
        RECT 121.510 17.720 121.830 17.780 ;
        RECT 1194.230 17.720 1194.550 17.780 ;
      LAYER via ;
        RECT 1194.260 1548.740 1194.520 1549.000 ;
        RECT 1194.260 1548.060 1194.520 1548.320 ;
        RECT 1194.260 992.160 1194.520 992.420 ;
        RECT 1194.260 990.120 1194.520 990.380 ;
        RECT 1194.260 798.360 1194.520 798.620 ;
        RECT 1194.260 796.660 1194.520 796.920 ;
        RECT 1194.260 738.520 1194.520 738.780 ;
        RECT 1194.260 737.840 1194.520 738.100 ;
        RECT 121.540 17.720 121.800 17.980 ;
        RECT 1194.260 17.720 1194.520 17.980 ;
      LAYER met2 ;
        RECT 1194.645 1700.000 1194.925 1704.000 ;
        RECT 1194.780 1656.210 1194.920 1700.000 ;
        RECT 1193.860 1656.070 1194.920 1656.210 ;
        RECT 1193.860 1654.850 1194.000 1656.070 ;
        RECT 1193.860 1654.710 1194.460 1654.850 ;
        RECT 1194.320 1549.030 1194.460 1654.710 ;
        RECT 1194.260 1548.710 1194.520 1549.030 ;
        RECT 1194.260 1548.030 1194.520 1548.350 ;
        RECT 1194.320 992.450 1194.460 1548.030 ;
        RECT 1194.260 992.130 1194.520 992.450 ;
        RECT 1194.260 990.090 1194.520 990.410 ;
        RECT 1194.320 798.650 1194.460 990.090 ;
        RECT 1194.260 798.330 1194.520 798.650 ;
        RECT 1194.260 796.630 1194.520 796.950 ;
        RECT 1194.320 738.810 1194.460 796.630 ;
        RECT 1194.260 738.490 1194.520 738.810 ;
        RECT 1194.260 737.810 1194.520 738.130 ;
        RECT 1194.320 18.010 1194.460 737.810 ;
        RECT 121.540 17.690 121.800 18.010 ;
        RECT 1194.260 17.690 1194.520 18.010 ;
        RECT 121.600 2.400 121.740 17.690 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 1688.000 176.110 1688.060 ;
        RECT 1203.890 1688.000 1204.210 1688.060 ;
        RECT 175.790 1687.860 1204.210 1688.000 ;
        RECT 175.790 1687.800 176.110 1687.860 ;
        RECT 1203.890 1687.800 1204.210 1687.860 ;
        RECT 145.430 16.560 145.750 16.620 ;
        RECT 175.790 16.560 176.110 16.620 ;
        RECT 145.430 16.420 176.110 16.560 ;
        RECT 145.430 16.360 145.750 16.420 ;
        RECT 175.790 16.360 176.110 16.420 ;
      LAYER via ;
        RECT 175.820 1687.800 176.080 1688.060 ;
        RECT 1203.920 1687.800 1204.180 1688.060 ;
        RECT 145.460 16.360 145.720 16.620 ;
        RECT 175.820 16.360 176.080 16.620 ;
      LAYER met2 ;
        RECT 1203.845 1700.000 1204.125 1704.000 ;
        RECT 1203.980 1688.090 1204.120 1700.000 ;
        RECT 175.820 1687.770 176.080 1688.090 ;
        RECT 1203.920 1687.770 1204.180 1688.090 ;
        RECT 175.880 16.650 176.020 1687.770 ;
        RECT 145.460 16.330 145.720 16.650 ;
        RECT 175.820 16.330 176.080 16.650 ;
        RECT 145.520 2.400 145.660 16.330 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1207.570 1678.140 1207.890 1678.200 ;
        RECT 1208.950 1678.140 1209.270 1678.200 ;
        RECT 1207.570 1678.000 1209.270 1678.140 ;
        RECT 1207.570 1677.940 1207.890 1678.000 ;
        RECT 1208.950 1677.940 1209.270 1678.000 ;
        RECT 163.370 18.600 163.690 18.660 ;
        RECT 1207.570 18.600 1207.890 18.660 ;
        RECT 163.370 18.460 1207.890 18.600 ;
        RECT 163.370 18.400 163.690 18.460 ;
        RECT 1207.570 18.400 1207.890 18.460 ;
      LAYER via ;
        RECT 1207.600 1677.940 1207.860 1678.200 ;
        RECT 1208.980 1677.940 1209.240 1678.200 ;
        RECT 163.400 18.400 163.660 18.660 ;
        RECT 1207.600 18.400 1207.860 18.660 ;
      LAYER met2 ;
        RECT 1210.285 1700.410 1210.565 1704.000 ;
        RECT 1209.040 1700.270 1210.565 1700.410 ;
        RECT 1209.040 1678.230 1209.180 1700.270 ;
        RECT 1210.285 1700.000 1210.565 1700.270 ;
        RECT 1207.600 1677.910 1207.860 1678.230 ;
        RECT 1208.980 1677.910 1209.240 1678.230 ;
        RECT 1207.660 18.690 1207.800 1677.910 ;
        RECT 163.400 18.370 163.660 18.690 ;
        RECT 1207.600 18.370 1207.860 18.690 ;
        RECT 163.460 2.400 163.600 18.370 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 196.490 1688.340 196.810 1688.400 ;
        RECT 1217.230 1688.340 1217.550 1688.400 ;
        RECT 196.490 1688.200 1217.550 1688.340 ;
        RECT 196.490 1688.140 196.810 1688.200 ;
        RECT 1217.230 1688.140 1217.550 1688.200 ;
        RECT 180.850 20.640 181.170 20.700 ;
        RECT 196.490 20.640 196.810 20.700 ;
        RECT 180.850 20.500 196.810 20.640 ;
        RECT 180.850 20.440 181.170 20.500 ;
        RECT 196.490 20.440 196.810 20.500 ;
      LAYER via ;
        RECT 196.520 1688.140 196.780 1688.400 ;
        RECT 1217.260 1688.140 1217.520 1688.400 ;
        RECT 180.880 20.440 181.140 20.700 ;
        RECT 196.520 20.440 196.780 20.700 ;
      LAYER met2 ;
        RECT 1217.185 1700.000 1217.465 1704.000 ;
        RECT 1217.320 1688.430 1217.460 1700.000 ;
        RECT 196.520 1688.110 196.780 1688.430 ;
        RECT 1217.260 1688.110 1217.520 1688.430 ;
        RECT 196.580 20.730 196.720 1688.110 ;
        RECT 180.880 20.410 181.140 20.730 ;
        RECT 196.520 20.410 196.780 20.730 ;
        RECT 180.940 2.400 181.080 20.410 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1221.445 1304.325 1221.615 1352.435 ;
        RECT 1221.445 1207.425 1221.615 1255.875 ;
        RECT 1221.445 289.765 1221.615 337.875 ;
      LAYER mcon ;
        RECT 1221.445 1352.265 1221.615 1352.435 ;
        RECT 1221.445 1255.705 1221.615 1255.875 ;
        RECT 1221.445 337.705 1221.615 337.875 ;
      LAYER met1 ;
        RECT 1222.290 1656.720 1222.610 1656.780 ;
        RECT 1221.460 1656.580 1222.610 1656.720 ;
        RECT 1221.460 1656.100 1221.600 1656.580 ;
        RECT 1222.290 1656.520 1222.610 1656.580 ;
        RECT 1221.370 1655.840 1221.690 1656.100 ;
        RECT 1220.910 1497.940 1221.230 1498.000 ;
        RECT 1220.910 1497.800 1221.600 1497.940 ;
        RECT 1220.910 1497.740 1221.230 1497.800 ;
        RECT 1221.460 1497.660 1221.600 1497.800 ;
        RECT 1221.370 1497.400 1221.690 1497.660 ;
        RECT 1221.370 1352.420 1221.690 1352.480 ;
        RECT 1221.175 1352.280 1221.690 1352.420 ;
        RECT 1221.370 1352.220 1221.690 1352.280 ;
        RECT 1221.370 1304.480 1221.690 1304.540 ;
        RECT 1221.175 1304.340 1221.690 1304.480 ;
        RECT 1221.370 1304.280 1221.690 1304.340 ;
        RECT 1221.370 1255.860 1221.690 1255.920 ;
        RECT 1221.175 1255.720 1221.690 1255.860 ;
        RECT 1221.370 1255.660 1221.690 1255.720 ;
        RECT 1221.370 1207.580 1221.690 1207.640 ;
        RECT 1221.175 1207.440 1221.690 1207.580 ;
        RECT 1221.370 1207.380 1221.690 1207.440 ;
        RECT 1220.910 1111.020 1221.230 1111.080 ;
        RECT 1221.370 1111.020 1221.690 1111.080 ;
        RECT 1220.910 1110.880 1221.690 1111.020 ;
        RECT 1220.910 1110.820 1221.230 1110.880 ;
        RECT 1221.370 1110.820 1221.690 1110.880 ;
        RECT 1220.450 966.180 1220.770 966.240 ;
        RECT 1221.370 966.180 1221.690 966.240 ;
        RECT 1220.450 966.040 1221.690 966.180 ;
        RECT 1220.450 965.980 1220.770 966.040 ;
        RECT 1221.370 965.980 1221.690 966.040 ;
        RECT 1221.370 947.140 1221.690 947.200 ;
        RECT 1222.290 947.140 1222.610 947.200 ;
        RECT 1221.370 947.000 1222.610 947.140 ;
        RECT 1221.370 946.940 1221.690 947.000 ;
        RECT 1222.290 946.940 1222.610 947.000 ;
        RECT 1221.370 869.620 1221.690 869.680 ;
        RECT 1222.290 869.620 1222.610 869.680 ;
        RECT 1221.370 869.480 1222.610 869.620 ;
        RECT 1221.370 869.420 1221.690 869.480 ;
        RECT 1222.290 869.420 1222.610 869.480 ;
        RECT 1220.450 724.440 1220.770 724.500 ;
        RECT 1221.370 724.440 1221.690 724.500 ;
        RECT 1220.450 724.300 1221.690 724.440 ;
        RECT 1220.450 724.240 1220.770 724.300 ;
        RECT 1221.370 724.240 1221.690 724.300 ;
        RECT 1221.370 337.860 1221.690 337.920 ;
        RECT 1221.175 337.720 1221.690 337.860 ;
        RECT 1221.370 337.660 1221.690 337.720 ;
        RECT 1221.370 289.920 1221.690 289.980 ;
        RECT 1221.175 289.780 1221.690 289.920 ;
        RECT 1221.370 289.720 1221.690 289.780 ;
        RECT 198.790 19.280 199.110 19.340 ;
        RECT 1221.370 19.280 1221.690 19.340 ;
        RECT 198.790 19.140 1221.690 19.280 ;
        RECT 198.790 19.080 199.110 19.140 ;
        RECT 1221.370 19.080 1221.690 19.140 ;
      LAYER via ;
        RECT 1222.320 1656.520 1222.580 1656.780 ;
        RECT 1221.400 1655.840 1221.660 1656.100 ;
        RECT 1220.940 1497.740 1221.200 1498.000 ;
        RECT 1221.400 1497.400 1221.660 1497.660 ;
        RECT 1221.400 1352.220 1221.660 1352.480 ;
        RECT 1221.400 1304.280 1221.660 1304.540 ;
        RECT 1221.400 1255.660 1221.660 1255.920 ;
        RECT 1221.400 1207.380 1221.660 1207.640 ;
        RECT 1220.940 1110.820 1221.200 1111.080 ;
        RECT 1221.400 1110.820 1221.660 1111.080 ;
        RECT 1220.480 965.980 1220.740 966.240 ;
        RECT 1221.400 965.980 1221.660 966.240 ;
        RECT 1221.400 946.940 1221.660 947.200 ;
        RECT 1222.320 946.940 1222.580 947.200 ;
        RECT 1221.400 869.420 1221.660 869.680 ;
        RECT 1222.320 869.420 1222.580 869.680 ;
        RECT 1220.480 724.240 1220.740 724.500 ;
        RECT 1221.400 724.240 1221.660 724.500 ;
        RECT 1221.400 337.660 1221.660 337.920 ;
        RECT 1221.400 289.720 1221.660 289.980 ;
        RECT 198.820 19.080 199.080 19.340 ;
        RECT 1221.400 19.080 1221.660 19.340 ;
      LAYER met2 ;
        RECT 1224.085 1700.410 1224.365 1704.000 ;
        RECT 1222.380 1700.270 1224.365 1700.410 ;
        RECT 1222.380 1656.810 1222.520 1700.270 ;
        RECT 1224.085 1700.000 1224.365 1700.270 ;
        RECT 1222.320 1656.490 1222.580 1656.810 ;
        RECT 1221.400 1655.810 1221.660 1656.130 ;
        RECT 1221.460 1545.370 1221.600 1655.810 ;
        RECT 1221.000 1545.230 1221.600 1545.370 ;
        RECT 1221.000 1498.030 1221.140 1545.230 ;
        RECT 1220.940 1497.710 1221.200 1498.030 ;
        RECT 1221.400 1497.370 1221.660 1497.690 ;
        RECT 1221.460 1352.510 1221.600 1497.370 ;
        RECT 1221.400 1352.190 1221.660 1352.510 ;
        RECT 1221.400 1304.250 1221.660 1304.570 ;
        RECT 1221.460 1255.950 1221.600 1304.250 ;
        RECT 1221.400 1255.630 1221.660 1255.950 ;
        RECT 1221.400 1207.350 1221.660 1207.670 ;
        RECT 1221.460 1159.130 1221.600 1207.350 ;
        RECT 1221.000 1158.990 1221.600 1159.130 ;
        RECT 1221.000 1111.110 1221.140 1158.990 ;
        RECT 1220.940 1110.790 1221.200 1111.110 ;
        RECT 1221.400 1110.790 1221.660 1111.110 ;
        RECT 1221.460 1014.405 1221.600 1110.790 ;
        RECT 1220.470 1014.035 1220.750 1014.405 ;
        RECT 1221.390 1014.035 1221.670 1014.405 ;
        RECT 1220.540 966.270 1220.680 1014.035 ;
        RECT 1220.480 965.950 1220.740 966.270 ;
        RECT 1221.400 965.950 1221.660 966.270 ;
        RECT 1221.460 947.230 1221.600 965.950 ;
        RECT 1221.400 946.910 1221.660 947.230 ;
        RECT 1222.320 946.910 1222.580 947.230 ;
        RECT 1222.380 869.710 1222.520 946.910 ;
        RECT 1221.400 869.390 1221.660 869.710 ;
        RECT 1222.320 869.390 1222.580 869.710 ;
        RECT 1221.460 724.530 1221.600 869.390 ;
        RECT 1220.480 724.210 1220.740 724.530 ;
        RECT 1221.400 724.210 1221.660 724.530 ;
        RECT 1220.540 676.445 1220.680 724.210 ;
        RECT 1220.470 676.075 1220.750 676.445 ;
        RECT 1221.390 676.075 1221.670 676.445 ;
        RECT 1221.460 337.950 1221.600 676.075 ;
        RECT 1221.400 337.630 1221.660 337.950 ;
        RECT 1221.400 289.690 1221.660 290.010 ;
        RECT 1221.460 19.370 1221.600 289.690 ;
        RECT 198.820 19.050 199.080 19.370 ;
        RECT 1221.400 19.050 1221.660 19.370 ;
        RECT 198.880 2.400 199.020 19.050 ;
        RECT 198.670 -4.800 199.230 2.400 ;
      LAYER via2 ;
        RECT 1220.470 1014.080 1220.750 1014.360 ;
        RECT 1221.390 1014.080 1221.670 1014.360 ;
        RECT 1220.470 676.120 1220.750 676.400 ;
        RECT 1221.390 676.120 1221.670 676.400 ;
      LAYER met3 ;
        RECT 1220.445 1014.370 1220.775 1014.385 ;
        RECT 1221.365 1014.370 1221.695 1014.385 ;
        RECT 1220.445 1014.070 1221.695 1014.370 ;
        RECT 1220.445 1014.055 1220.775 1014.070 ;
        RECT 1221.365 1014.055 1221.695 1014.070 ;
        RECT 1220.445 676.410 1220.775 676.425 ;
        RECT 1221.365 676.410 1221.695 676.425 ;
        RECT 1220.445 676.110 1221.695 676.410 ;
        RECT 1220.445 676.095 1220.775 676.110 ;
        RECT 1221.365 676.095 1221.695 676.110 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 306.890 1689.360 307.210 1689.420 ;
        RECT 1230.570 1689.360 1230.890 1689.420 ;
        RECT 306.890 1689.220 1230.890 1689.360 ;
        RECT 306.890 1689.160 307.210 1689.220 ;
        RECT 1230.570 1689.160 1230.890 1689.220 ;
        RECT 216.730 16.220 217.050 16.280 ;
        RECT 306.890 16.220 307.210 16.280 ;
        RECT 216.730 16.080 307.210 16.220 ;
        RECT 216.730 16.020 217.050 16.080 ;
        RECT 306.890 16.020 307.210 16.080 ;
      LAYER via ;
        RECT 306.920 1689.160 307.180 1689.420 ;
        RECT 1230.600 1689.160 1230.860 1689.420 ;
        RECT 216.760 16.020 217.020 16.280 ;
        RECT 306.920 16.020 307.180 16.280 ;
      LAYER met2 ;
        RECT 1230.525 1700.000 1230.805 1704.000 ;
        RECT 1230.660 1689.450 1230.800 1700.000 ;
        RECT 306.920 1689.130 307.180 1689.450 ;
        RECT 1230.600 1689.130 1230.860 1689.450 ;
        RECT 306.980 16.310 307.120 1689.130 ;
        RECT 216.760 15.990 217.020 16.310 ;
        RECT 306.920 15.990 307.180 16.310 ;
        RECT 216.820 2.400 216.960 15.990 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 234.670 19.960 234.990 20.020 ;
        RECT 1236.090 19.960 1236.410 20.020 ;
        RECT 234.670 19.820 1236.410 19.960 ;
        RECT 234.670 19.760 234.990 19.820 ;
        RECT 1236.090 19.760 1236.410 19.820 ;
      LAYER via ;
        RECT 234.700 19.760 234.960 20.020 ;
        RECT 1236.120 19.760 1236.380 20.020 ;
      LAYER met2 ;
        RECT 1237.425 1700.410 1237.705 1704.000 ;
        RECT 1236.180 1700.270 1237.705 1700.410 ;
        RECT 1236.180 20.050 1236.320 1700.270 ;
        RECT 1237.425 1700.000 1237.705 1700.270 ;
        RECT 234.700 19.730 234.960 20.050 ;
        RECT 1236.120 19.730 1236.380 20.050 ;
        RECT 234.760 2.400 234.900 19.730 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1149.685 1687.335 1149.855 1688.695 ;
        RECT 1148.305 1687.165 1149.855 1687.335 ;
      LAYER mcon ;
        RECT 1149.685 1688.525 1149.855 1688.695 ;
      LAYER met1 ;
        RECT 1149.625 1688.680 1149.915 1688.725 ;
        RECT 1169.850 1688.680 1170.170 1688.740 ;
        RECT 1149.625 1688.540 1170.170 1688.680 ;
        RECT 1149.625 1688.495 1149.915 1688.540 ;
        RECT 1169.850 1688.480 1170.170 1688.540 ;
        RECT 99.890 1687.320 100.210 1687.380 ;
        RECT 1148.245 1687.320 1148.535 1687.365 ;
        RECT 99.890 1687.180 1148.535 1687.320 ;
        RECT 99.890 1687.120 100.210 1687.180 ;
        RECT 1148.245 1687.135 1148.535 1687.180 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 99.890 17.920 100.210 17.980 ;
        RECT 56.190 17.780 100.210 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 99.890 17.720 100.210 17.780 ;
      LAYER via ;
        RECT 1169.880 1688.480 1170.140 1688.740 ;
        RECT 99.920 1687.120 100.180 1687.380 ;
        RECT 56.220 17.720 56.480 17.980 ;
        RECT 99.920 17.720 100.180 17.980 ;
      LAYER met2 ;
        RECT 1169.805 1700.000 1170.085 1704.000 ;
        RECT 1169.940 1688.770 1170.080 1700.000 ;
        RECT 1169.880 1688.450 1170.140 1688.770 ;
        RECT 99.920 1687.090 100.180 1687.410 ;
        RECT 99.980 18.010 100.120 1687.090 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 99.920 17.690 100.180 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1175.445 1635.485 1175.615 1659.795 ;
        RECT 1175.445 1497.445 1175.615 1545.555 ;
        RECT 1175.445 1400.885 1175.615 1490.475 ;
        RECT 1175.445 1304.325 1175.615 1393.575 ;
        RECT 1175.445 1207.425 1175.615 1297.015 ;
        RECT 1175.445 1055.785 1175.615 1103.895 ;
        RECT 1174.985 758.965 1175.155 807.075 ;
        RECT 1175.445 614.125 1175.615 641.835 ;
        RECT 1174.525 83.045 1174.695 131.155 ;
      LAYER mcon ;
        RECT 1175.445 1659.625 1175.615 1659.795 ;
        RECT 1175.445 1545.385 1175.615 1545.555 ;
        RECT 1175.445 1490.305 1175.615 1490.475 ;
        RECT 1175.445 1393.405 1175.615 1393.575 ;
        RECT 1175.445 1296.845 1175.615 1297.015 ;
        RECT 1175.445 1103.725 1175.615 1103.895 ;
        RECT 1174.985 806.905 1175.155 807.075 ;
        RECT 1175.445 641.665 1175.615 641.835 ;
        RECT 1174.525 130.985 1174.695 131.155 ;
      LAYER met1 ;
        RECT 1175.385 1659.780 1175.675 1659.825 ;
        RECT 1177.210 1659.780 1177.530 1659.840 ;
        RECT 1175.385 1659.640 1177.530 1659.780 ;
        RECT 1175.385 1659.595 1175.675 1659.640 ;
        RECT 1177.210 1659.580 1177.530 1659.640 ;
        RECT 1175.370 1635.640 1175.690 1635.700 ;
        RECT 1175.175 1635.500 1175.690 1635.640 ;
        RECT 1175.370 1635.440 1175.690 1635.500 ;
        RECT 1175.370 1545.540 1175.690 1545.600 ;
        RECT 1175.175 1545.400 1175.690 1545.540 ;
        RECT 1175.370 1545.340 1175.690 1545.400 ;
        RECT 1175.370 1497.600 1175.690 1497.660 ;
        RECT 1175.175 1497.460 1175.690 1497.600 ;
        RECT 1175.370 1497.400 1175.690 1497.460 ;
        RECT 1175.370 1490.460 1175.690 1490.520 ;
        RECT 1175.175 1490.320 1175.690 1490.460 ;
        RECT 1175.370 1490.260 1175.690 1490.320 ;
        RECT 1175.370 1401.040 1175.690 1401.100 ;
        RECT 1175.175 1400.900 1175.690 1401.040 ;
        RECT 1175.370 1400.840 1175.690 1400.900 ;
        RECT 1175.370 1393.560 1175.690 1393.620 ;
        RECT 1175.175 1393.420 1175.690 1393.560 ;
        RECT 1175.370 1393.360 1175.690 1393.420 ;
        RECT 1175.370 1304.480 1175.690 1304.540 ;
        RECT 1175.175 1304.340 1175.690 1304.480 ;
        RECT 1175.370 1304.280 1175.690 1304.340 ;
        RECT 1175.370 1297.000 1175.690 1297.060 ;
        RECT 1175.175 1296.860 1175.690 1297.000 ;
        RECT 1175.370 1296.800 1175.690 1296.860 ;
        RECT 1175.370 1207.580 1175.690 1207.640 ;
        RECT 1175.370 1207.440 1175.885 1207.580 ;
        RECT 1175.370 1207.380 1175.690 1207.440 ;
        RECT 1175.370 1152.500 1175.690 1152.560 ;
        RECT 1176.290 1152.500 1176.610 1152.560 ;
        RECT 1175.370 1152.360 1176.610 1152.500 ;
        RECT 1175.370 1152.300 1175.690 1152.360 ;
        RECT 1176.290 1152.300 1176.610 1152.360 ;
        RECT 1175.370 1111.500 1175.690 1111.760 ;
        RECT 1175.460 1111.080 1175.600 1111.500 ;
        RECT 1175.370 1110.820 1175.690 1111.080 ;
        RECT 1175.370 1103.880 1175.690 1103.940 ;
        RECT 1175.175 1103.740 1175.690 1103.880 ;
        RECT 1175.370 1103.680 1175.690 1103.740 ;
        RECT 1175.370 1055.940 1175.690 1056.000 ;
        RECT 1175.175 1055.800 1175.690 1055.940 ;
        RECT 1175.370 1055.740 1175.690 1055.800 ;
        RECT 1175.370 965.980 1175.690 966.240 ;
        RECT 1175.460 965.840 1175.600 965.980 ;
        RECT 1176.290 965.840 1176.610 965.900 ;
        RECT 1175.460 965.700 1176.610 965.840 ;
        RECT 1176.290 965.640 1176.610 965.700 ;
        RECT 1174.910 917.900 1175.230 917.960 ;
        RECT 1176.290 917.900 1176.610 917.960 ;
        RECT 1174.910 917.760 1176.610 917.900 ;
        RECT 1174.910 917.700 1175.230 917.760 ;
        RECT 1176.290 917.700 1176.610 917.760 ;
        RECT 1174.910 896.820 1175.230 896.880 ;
        RECT 1175.830 896.820 1176.150 896.880 ;
        RECT 1174.910 896.680 1176.150 896.820 ;
        RECT 1174.910 896.620 1175.230 896.680 ;
        RECT 1175.830 896.620 1176.150 896.680 ;
        RECT 1174.910 814.880 1175.230 814.940 ;
        RECT 1175.830 814.880 1176.150 814.940 ;
        RECT 1174.910 814.740 1176.150 814.880 ;
        RECT 1174.910 814.680 1175.230 814.740 ;
        RECT 1175.830 814.680 1176.150 814.740 ;
        RECT 1174.910 807.060 1175.230 807.120 ;
        RECT 1174.715 806.920 1175.230 807.060 ;
        RECT 1174.910 806.860 1175.230 806.920 ;
        RECT 1174.925 759.120 1175.215 759.165 ;
        RECT 1175.370 759.120 1175.690 759.180 ;
        RECT 1174.925 758.980 1175.690 759.120 ;
        RECT 1174.925 758.935 1175.215 758.980 ;
        RECT 1175.370 758.920 1175.690 758.980 ;
        RECT 1175.370 641.820 1175.690 641.880 ;
        RECT 1175.175 641.680 1175.690 641.820 ;
        RECT 1175.370 641.620 1175.690 641.680 ;
        RECT 1175.370 614.280 1175.690 614.340 ;
        RECT 1175.175 614.140 1175.690 614.280 ;
        RECT 1175.370 614.080 1175.690 614.140 ;
        RECT 1174.910 572.460 1175.230 572.520 ;
        RECT 1175.370 572.460 1175.690 572.520 ;
        RECT 1174.910 572.320 1175.690 572.460 ;
        RECT 1174.910 572.260 1175.230 572.320 ;
        RECT 1175.370 572.260 1175.690 572.320 ;
        RECT 1174.910 524.180 1175.230 524.240 ;
        RECT 1175.370 524.180 1175.690 524.240 ;
        RECT 1174.910 524.040 1175.690 524.180 ;
        RECT 1174.910 523.980 1175.230 524.040 ;
        RECT 1175.370 523.980 1175.690 524.040 ;
        RECT 1174.910 386.480 1175.230 386.540 ;
        RECT 1175.370 386.480 1175.690 386.540 ;
        RECT 1174.910 386.340 1175.690 386.480 ;
        RECT 1174.910 386.280 1175.230 386.340 ;
        RECT 1175.370 386.280 1175.690 386.340 ;
        RECT 1174.910 227.700 1175.230 227.760 ;
        RECT 1175.830 227.700 1176.150 227.760 ;
        RECT 1174.910 227.560 1176.150 227.700 ;
        RECT 1174.910 227.500 1175.230 227.560 ;
        RECT 1175.830 227.500 1176.150 227.560 ;
        RECT 1174.465 131.140 1174.755 131.185 ;
        RECT 1175.370 131.140 1175.690 131.200 ;
        RECT 1174.465 131.000 1175.690 131.140 ;
        RECT 1174.465 130.955 1174.755 131.000 ;
        RECT 1175.370 130.940 1175.690 131.000 ;
        RECT 1174.450 83.200 1174.770 83.260 ;
        RECT 1174.255 83.060 1174.770 83.200 ;
        RECT 1174.450 83.000 1174.770 83.060 ;
        RECT 1174.450 41.720 1174.770 41.780 ;
        RECT 1175.370 41.720 1175.690 41.780 ;
        RECT 1174.450 41.580 1175.690 41.720 ;
        RECT 1174.450 41.520 1174.770 41.580 ;
        RECT 1175.370 41.520 1175.690 41.580 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 1175.370 17.580 1175.690 17.640 ;
        RECT 80.110 17.440 1175.690 17.580 ;
        RECT 80.110 17.380 80.430 17.440 ;
        RECT 1175.370 17.380 1175.690 17.440 ;
      LAYER via ;
        RECT 1177.240 1659.580 1177.500 1659.840 ;
        RECT 1175.400 1635.440 1175.660 1635.700 ;
        RECT 1175.400 1545.340 1175.660 1545.600 ;
        RECT 1175.400 1497.400 1175.660 1497.660 ;
        RECT 1175.400 1490.260 1175.660 1490.520 ;
        RECT 1175.400 1400.840 1175.660 1401.100 ;
        RECT 1175.400 1393.360 1175.660 1393.620 ;
        RECT 1175.400 1304.280 1175.660 1304.540 ;
        RECT 1175.400 1296.800 1175.660 1297.060 ;
        RECT 1175.400 1207.380 1175.660 1207.640 ;
        RECT 1175.400 1152.300 1175.660 1152.560 ;
        RECT 1176.320 1152.300 1176.580 1152.560 ;
        RECT 1175.400 1111.500 1175.660 1111.760 ;
        RECT 1175.400 1110.820 1175.660 1111.080 ;
        RECT 1175.400 1103.680 1175.660 1103.940 ;
        RECT 1175.400 1055.740 1175.660 1056.000 ;
        RECT 1175.400 965.980 1175.660 966.240 ;
        RECT 1176.320 965.640 1176.580 965.900 ;
        RECT 1174.940 917.700 1175.200 917.960 ;
        RECT 1176.320 917.700 1176.580 917.960 ;
        RECT 1174.940 896.620 1175.200 896.880 ;
        RECT 1175.860 896.620 1176.120 896.880 ;
        RECT 1174.940 814.680 1175.200 814.940 ;
        RECT 1175.860 814.680 1176.120 814.940 ;
        RECT 1174.940 806.860 1175.200 807.120 ;
        RECT 1175.400 758.920 1175.660 759.180 ;
        RECT 1175.400 641.620 1175.660 641.880 ;
        RECT 1175.400 614.080 1175.660 614.340 ;
        RECT 1174.940 572.260 1175.200 572.520 ;
        RECT 1175.400 572.260 1175.660 572.520 ;
        RECT 1174.940 523.980 1175.200 524.240 ;
        RECT 1175.400 523.980 1175.660 524.240 ;
        RECT 1174.940 386.280 1175.200 386.540 ;
        RECT 1175.400 386.280 1175.660 386.540 ;
        RECT 1174.940 227.500 1175.200 227.760 ;
        RECT 1175.860 227.500 1176.120 227.760 ;
        RECT 1175.400 130.940 1175.660 131.200 ;
        RECT 1174.480 83.000 1174.740 83.260 ;
        RECT 1174.480 41.520 1174.740 41.780 ;
        RECT 1175.400 41.520 1175.660 41.780 ;
        RECT 80.140 17.380 80.400 17.640 ;
        RECT 1175.400 17.380 1175.660 17.640 ;
      LAYER met2 ;
        RECT 1179.005 1700.410 1179.285 1704.000 ;
        RECT 1177.300 1700.270 1179.285 1700.410 ;
        RECT 1177.300 1659.870 1177.440 1700.270 ;
        RECT 1179.005 1700.000 1179.285 1700.270 ;
        RECT 1177.240 1659.550 1177.500 1659.870 ;
        RECT 1175.400 1635.410 1175.660 1635.730 ;
        RECT 1175.460 1545.630 1175.600 1635.410 ;
        RECT 1175.400 1545.310 1175.660 1545.630 ;
        RECT 1175.400 1497.370 1175.660 1497.690 ;
        RECT 1175.460 1490.550 1175.600 1497.370 ;
        RECT 1175.400 1490.230 1175.660 1490.550 ;
        RECT 1175.400 1400.810 1175.660 1401.130 ;
        RECT 1175.460 1393.650 1175.600 1400.810 ;
        RECT 1175.400 1393.330 1175.660 1393.650 ;
        RECT 1175.400 1304.250 1175.660 1304.570 ;
        RECT 1175.460 1297.090 1175.600 1304.250 ;
        RECT 1175.400 1296.770 1175.660 1297.090 ;
        RECT 1175.400 1207.350 1175.660 1207.670 ;
        RECT 1175.460 1200.725 1175.600 1207.350 ;
        RECT 1175.390 1200.355 1175.670 1200.725 ;
        RECT 1176.310 1200.355 1176.590 1200.725 ;
        RECT 1176.380 1152.590 1176.520 1200.355 ;
        RECT 1175.400 1152.270 1175.660 1152.590 ;
        RECT 1176.320 1152.270 1176.580 1152.590 ;
        RECT 1175.460 1111.790 1175.600 1152.270 ;
        RECT 1175.400 1111.470 1175.660 1111.790 ;
        RECT 1175.400 1110.790 1175.660 1111.110 ;
        RECT 1175.460 1103.970 1175.600 1110.790 ;
        RECT 1175.400 1103.650 1175.660 1103.970 ;
        RECT 1175.400 1055.710 1175.660 1056.030 ;
        RECT 1175.460 1029.250 1175.600 1055.710 ;
        RECT 1175.000 1029.110 1175.600 1029.250 ;
        RECT 1175.000 1027.890 1175.140 1029.110 ;
        RECT 1175.000 1027.750 1175.600 1027.890 ;
        RECT 1175.460 966.270 1175.600 1027.750 ;
        RECT 1175.400 965.950 1175.660 966.270 ;
        RECT 1176.320 965.610 1176.580 965.930 ;
        RECT 1176.380 917.990 1176.520 965.610 ;
        RECT 1174.940 917.670 1175.200 917.990 ;
        RECT 1176.320 917.670 1176.580 917.990 ;
        RECT 1175.000 896.910 1175.140 917.670 ;
        RECT 1174.940 896.590 1175.200 896.910 ;
        RECT 1175.860 896.590 1176.120 896.910 ;
        RECT 1175.920 814.970 1176.060 896.590 ;
        RECT 1174.940 814.650 1175.200 814.970 ;
        RECT 1175.860 814.650 1176.120 814.970 ;
        RECT 1175.000 807.150 1175.140 814.650 ;
        RECT 1174.940 806.830 1175.200 807.150 ;
        RECT 1175.400 758.890 1175.660 759.210 ;
        RECT 1175.460 718.605 1175.600 758.890 ;
        RECT 1175.390 718.235 1175.670 718.605 ;
        RECT 1175.850 717.555 1176.130 717.925 ;
        RECT 1175.920 662.730 1176.060 717.555 ;
        RECT 1175.460 662.590 1176.060 662.730 ;
        RECT 1175.460 641.910 1175.600 662.590 ;
        RECT 1175.400 641.590 1175.660 641.910 ;
        RECT 1175.400 614.050 1175.660 614.370 ;
        RECT 1175.460 572.550 1175.600 614.050 ;
        RECT 1174.940 572.230 1175.200 572.550 ;
        RECT 1175.400 572.230 1175.660 572.550 ;
        RECT 1175.000 524.270 1175.140 572.230 ;
        RECT 1174.940 523.950 1175.200 524.270 ;
        RECT 1175.400 523.950 1175.660 524.270 ;
        RECT 1175.460 386.570 1175.600 523.950 ;
        RECT 1174.940 386.250 1175.200 386.570 ;
        RECT 1175.400 386.250 1175.660 386.570 ;
        RECT 1175.000 265.610 1175.140 386.250 ;
        RECT 1175.000 265.470 1176.060 265.610 ;
        RECT 1175.920 227.790 1176.060 265.470 ;
        RECT 1174.940 227.470 1175.200 227.790 ;
        RECT 1175.860 227.470 1176.120 227.790 ;
        RECT 1175.000 179.930 1175.140 227.470 ;
        RECT 1175.000 179.790 1175.600 179.930 ;
        RECT 1175.460 131.230 1175.600 179.790 ;
        RECT 1175.400 130.910 1175.660 131.230 ;
        RECT 1174.480 82.970 1174.740 83.290 ;
        RECT 1174.540 41.810 1174.680 82.970 ;
        RECT 1174.480 41.490 1174.740 41.810 ;
        RECT 1175.400 41.490 1175.660 41.810 ;
        RECT 1175.460 17.670 1175.600 41.490 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 1175.400 17.350 1175.660 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 1175.390 1200.400 1175.670 1200.680 ;
        RECT 1176.310 1200.400 1176.590 1200.680 ;
        RECT 1175.390 718.280 1175.670 718.560 ;
        RECT 1175.850 717.600 1176.130 717.880 ;
      LAYER met3 ;
        RECT 1175.365 1200.690 1175.695 1200.705 ;
        RECT 1176.285 1200.690 1176.615 1200.705 ;
        RECT 1175.365 1200.390 1176.615 1200.690 ;
        RECT 1175.365 1200.375 1175.695 1200.390 ;
        RECT 1176.285 1200.375 1176.615 1200.390 ;
        RECT 1175.365 718.570 1175.695 718.585 ;
        RECT 1175.150 718.255 1175.695 718.570 ;
        RECT 1175.150 717.890 1175.450 718.255 ;
        RECT 1175.825 717.890 1176.155 717.905 ;
        RECT 1175.150 717.590 1176.155 717.890 ;
        RECT 1175.825 717.575 1176.155 717.590 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1149.225 1687.505 1149.395 1688.695 ;
      LAYER mcon ;
        RECT 1149.225 1688.525 1149.395 1688.695 ;
      LAYER met1 ;
        RECT 210.290 1688.680 210.610 1688.740 ;
        RECT 1149.165 1688.680 1149.455 1688.725 ;
        RECT 210.290 1688.540 1149.455 1688.680 ;
        RECT 210.290 1688.480 210.610 1688.540 ;
        RECT 1149.165 1688.495 1149.455 1688.540 ;
        RECT 1149.165 1687.660 1149.455 1687.705 ;
        RECT 1187.790 1687.660 1188.110 1687.720 ;
        RECT 1149.165 1687.520 1188.110 1687.660 ;
        RECT 1149.165 1687.475 1149.455 1687.520 ;
        RECT 1187.790 1687.460 1188.110 1687.520 ;
        RECT 103.570 19.620 103.890 19.680 ;
        RECT 210.290 19.620 210.610 19.680 ;
        RECT 103.570 19.480 210.610 19.620 ;
        RECT 103.570 19.420 103.890 19.480 ;
        RECT 210.290 19.420 210.610 19.480 ;
      LAYER via ;
        RECT 210.320 1688.480 210.580 1688.740 ;
        RECT 1187.820 1687.460 1188.080 1687.720 ;
        RECT 103.600 19.420 103.860 19.680 ;
        RECT 210.320 19.420 210.580 19.680 ;
      LAYER met2 ;
        RECT 1187.745 1700.000 1188.025 1704.000 ;
        RECT 210.320 1688.450 210.580 1688.770 ;
        RECT 210.380 19.710 210.520 1688.450 ;
        RECT 1187.880 1687.750 1188.020 1700.000 ;
        RECT 1187.820 1687.430 1188.080 1687.750 ;
        RECT 103.600 19.390 103.860 19.710 ;
        RECT 210.320 19.390 210.580 19.710 ;
        RECT 103.660 2.400 103.800 19.390 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1193.310 1666.580 1193.630 1666.640 ;
        RECT 1195.150 1666.580 1195.470 1666.640 ;
        RECT 1193.310 1666.440 1195.470 1666.580 ;
        RECT 1193.310 1666.380 1193.630 1666.440 ;
        RECT 1195.150 1666.380 1195.470 1666.440 ;
        RECT 1193.770 1607.760 1194.090 1607.820 ;
        RECT 1194.690 1607.760 1195.010 1607.820 ;
        RECT 1193.770 1607.620 1195.010 1607.760 ;
        RECT 1193.770 1607.560 1194.090 1607.620 ;
        RECT 1194.690 1607.560 1195.010 1607.620 ;
        RECT 1193.770 1022.960 1194.090 1023.020 ;
        RECT 1194.690 1022.960 1195.010 1023.020 ;
        RECT 1193.770 1022.820 1195.010 1022.960 ;
        RECT 1193.770 1022.760 1194.090 1022.820 ;
        RECT 1194.690 1022.760 1195.010 1022.820 ;
        RECT 1193.770 931.840 1194.090 931.900 ;
        RECT 1194.690 931.840 1195.010 931.900 ;
        RECT 1193.770 931.700 1195.010 931.840 ;
        RECT 1193.770 931.640 1194.090 931.700 ;
        RECT 1194.690 931.640 1195.010 931.700 ;
        RECT 1193.770 883.220 1194.090 883.280 ;
        RECT 1194.690 883.220 1195.010 883.280 ;
        RECT 1193.770 883.080 1195.010 883.220 ;
        RECT 1193.770 883.020 1194.090 883.080 ;
        RECT 1194.690 883.020 1195.010 883.080 ;
        RECT 1193.770 835.280 1194.090 835.340 ;
        RECT 1194.690 835.280 1195.010 835.340 ;
        RECT 1193.770 835.140 1195.010 835.280 ;
        RECT 1193.770 835.080 1194.090 835.140 ;
        RECT 1194.690 835.080 1195.010 835.140 ;
        RECT 1194.690 738.860 1195.010 739.120 ;
        RECT 1194.780 738.100 1194.920 738.860 ;
        RECT 1194.690 737.840 1195.010 738.100 ;
        RECT 1193.770 717.640 1194.090 717.700 ;
        RECT 1194.690 717.640 1195.010 717.700 ;
        RECT 1193.770 717.500 1195.010 717.640 ;
        RECT 1193.770 717.440 1194.090 717.500 ;
        RECT 1194.690 717.440 1195.010 717.500 ;
        RECT 1193.770 641.480 1194.090 641.540 ;
        RECT 1194.690 641.480 1195.010 641.540 ;
        RECT 1193.770 641.340 1195.010 641.480 ;
        RECT 1193.770 641.280 1194.090 641.340 ;
        RECT 1194.690 641.280 1195.010 641.340 ;
        RECT 1193.770 545.260 1194.090 545.320 ;
        RECT 1194.690 545.260 1195.010 545.320 ;
        RECT 1193.770 545.120 1195.010 545.260 ;
        RECT 1193.770 545.060 1194.090 545.120 ;
        RECT 1194.690 545.060 1195.010 545.120 ;
        RECT 127.490 18.260 127.810 18.320 ;
        RECT 1193.770 18.260 1194.090 18.320 ;
        RECT 127.490 18.120 1194.090 18.260 ;
        RECT 127.490 18.060 127.810 18.120 ;
        RECT 1193.770 18.060 1194.090 18.120 ;
      LAYER via ;
        RECT 1193.340 1666.380 1193.600 1666.640 ;
        RECT 1195.180 1666.380 1195.440 1666.640 ;
        RECT 1193.800 1607.560 1194.060 1607.820 ;
        RECT 1194.720 1607.560 1194.980 1607.820 ;
        RECT 1193.800 1022.760 1194.060 1023.020 ;
        RECT 1194.720 1022.760 1194.980 1023.020 ;
        RECT 1193.800 931.640 1194.060 931.900 ;
        RECT 1194.720 931.640 1194.980 931.900 ;
        RECT 1193.800 883.020 1194.060 883.280 ;
        RECT 1194.720 883.020 1194.980 883.280 ;
        RECT 1193.800 835.080 1194.060 835.340 ;
        RECT 1194.720 835.080 1194.980 835.340 ;
        RECT 1194.720 738.860 1194.980 739.120 ;
        RECT 1194.720 737.840 1194.980 738.100 ;
        RECT 1193.800 717.440 1194.060 717.700 ;
        RECT 1194.720 717.440 1194.980 717.700 ;
        RECT 1193.800 641.280 1194.060 641.540 ;
        RECT 1194.720 641.280 1194.980 641.540 ;
        RECT 1193.800 545.060 1194.060 545.320 ;
        RECT 1194.720 545.060 1194.980 545.320 ;
        RECT 127.520 18.060 127.780 18.320 ;
        RECT 1193.800 18.060 1194.060 18.320 ;
      LAYER met2 ;
        RECT 1196.945 1700.410 1197.225 1704.000 ;
        RECT 1195.240 1700.270 1197.225 1700.410 ;
        RECT 1195.240 1666.670 1195.380 1700.270 ;
        RECT 1196.945 1700.000 1197.225 1700.270 ;
        RECT 1193.340 1666.350 1193.600 1666.670 ;
        RECT 1195.180 1666.350 1195.440 1666.670 ;
        RECT 1193.400 1654.170 1193.540 1666.350 ;
        RECT 1193.400 1654.030 1194.000 1654.170 ;
        RECT 1193.860 1607.850 1194.000 1654.030 ;
        RECT 1193.800 1607.530 1194.060 1607.850 ;
        RECT 1194.720 1607.530 1194.980 1607.850 ;
        RECT 1194.780 1023.050 1194.920 1607.530 ;
        RECT 1193.800 1022.730 1194.060 1023.050 ;
        RECT 1194.720 1022.730 1194.980 1023.050 ;
        RECT 1193.860 991.850 1194.000 1022.730 ;
        RECT 1193.860 991.710 1194.920 991.850 ;
        RECT 1194.780 931.930 1194.920 991.710 ;
        RECT 1193.800 931.610 1194.060 931.930 ;
        RECT 1194.720 931.610 1194.980 931.930 ;
        RECT 1193.860 883.310 1194.000 931.610 ;
        RECT 1193.800 882.990 1194.060 883.310 ;
        RECT 1194.720 882.990 1194.980 883.310 ;
        RECT 1194.780 835.370 1194.920 882.990 ;
        RECT 1193.800 835.050 1194.060 835.370 ;
        RECT 1194.720 835.050 1194.980 835.370 ;
        RECT 1193.860 798.050 1194.000 835.050 ;
        RECT 1193.860 797.910 1194.920 798.050 ;
        RECT 1194.780 739.150 1194.920 797.910 ;
        RECT 1194.720 738.830 1194.980 739.150 ;
        RECT 1194.720 737.810 1194.980 738.130 ;
        RECT 1194.780 717.730 1194.920 737.810 ;
        RECT 1193.800 717.410 1194.060 717.730 ;
        RECT 1194.720 717.410 1194.980 717.730 ;
        RECT 1193.860 641.570 1194.000 717.410 ;
        RECT 1193.800 641.250 1194.060 641.570 ;
        RECT 1194.720 641.250 1194.980 641.570 ;
        RECT 1194.780 545.350 1194.920 641.250 ;
        RECT 1193.800 545.030 1194.060 545.350 ;
        RECT 1194.720 545.030 1194.980 545.350 ;
        RECT 1193.860 18.350 1194.000 545.030 ;
        RECT 127.520 18.030 127.780 18.350 ;
        RECT 1193.800 18.030 1194.060 18.350 ;
        RECT 127.580 2.400 127.720 18.030 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 20.640 26.610 20.700 ;
        RECT 51.590 20.640 51.910 20.700 ;
        RECT 26.290 20.500 51.910 20.640 ;
        RECT 26.290 20.440 26.610 20.500 ;
        RECT 51.590 20.440 51.910 20.500 ;
      LAYER via ;
        RECT 26.320 20.440 26.580 20.700 ;
        RECT 51.620 20.440 51.880 20.700 ;
      LAYER met2 ;
        RECT 1158.765 1700.000 1159.045 1704.000 ;
        RECT 1158.900 1686.925 1159.040 1700.000 ;
        RECT 51.610 1686.555 51.890 1686.925 ;
        RECT 1158.830 1686.555 1159.110 1686.925 ;
        RECT 51.680 20.730 51.820 1686.555 ;
        RECT 26.320 20.410 26.580 20.730 ;
        RECT 51.620 20.410 51.880 20.730 ;
        RECT 26.380 2.400 26.520 20.410 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 51.610 1686.600 51.890 1686.880 ;
        RECT 1158.830 1686.600 1159.110 1686.880 ;
      LAYER met3 ;
        RECT 51.585 1686.890 51.915 1686.905 ;
        RECT 1158.805 1686.890 1159.135 1686.905 ;
        RECT 51.585 1686.590 1159.135 1686.890 ;
        RECT 51.585 1686.575 51.915 1686.590 ;
        RECT 1158.805 1686.575 1159.135 1686.590 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.065 1700.410 1161.345 1704.000 ;
        RECT 1160.740 1700.270 1161.345 1700.410 ;
        RECT 1160.740 16.845 1160.880 1700.270 ;
        RECT 1161.065 1700.000 1161.345 1700.270 ;
        RECT 32.290 16.475 32.570 16.845 ;
        RECT 1160.670 16.475 1160.950 16.845 ;
        RECT 32.360 2.400 32.500 16.475 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 32.290 16.520 32.570 16.800 ;
        RECT 1160.670 16.520 1160.950 16.800 ;
      LAYER met3 ;
        RECT 32.265 16.810 32.595 16.825 ;
        RECT 1160.645 16.810 1160.975 16.825 ;
        RECT 32.265 16.510 1160.975 16.810 ;
        RECT 32.265 16.495 32.595 16.510 ;
        RECT 1160.645 16.495 1160.975 16.510 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1154.535 1710.795 2243.355 2788.085 ;
      LAYER met1 ;
        RECT 1154.145 1707.860 2247.885 2796.120 ;
      LAYER met2 ;
        RECT 1150.025 2795.720 1153.425 2796.150 ;
        RECT 1154.265 2795.720 1162.625 2796.150 ;
        RECT 1163.465 2795.720 1172.285 2796.150 ;
        RECT 1173.125 2795.720 1181.945 2796.150 ;
        RECT 1182.785 2795.720 1191.605 2796.150 ;
        RECT 1192.445 2795.720 1201.265 2796.150 ;
        RECT 1202.105 2795.720 1210.925 2796.150 ;
        RECT 1211.765 2795.720 1220.585 2796.150 ;
        RECT 1221.425 2795.720 1230.245 2796.150 ;
        RECT 1231.085 2795.720 1239.905 2796.150 ;
        RECT 1240.745 2795.720 1249.565 2796.150 ;
        RECT 1250.405 2795.720 1259.225 2796.150 ;
        RECT 1260.065 2795.720 1268.885 2796.150 ;
        RECT 1269.725 2795.720 1278.545 2796.150 ;
        RECT 1279.385 2795.720 1288.205 2796.150 ;
        RECT 1289.045 2795.720 1297.865 2796.150 ;
        RECT 1298.705 2795.720 1307.525 2796.150 ;
        RECT 1308.365 2795.720 1317.185 2796.150 ;
        RECT 1318.025 2795.720 1326.845 2796.150 ;
        RECT 1327.685 2795.720 1336.505 2796.150 ;
        RECT 1337.345 2795.720 1346.165 2796.150 ;
        RECT 1347.005 2795.720 1355.825 2796.150 ;
        RECT 1356.665 2795.720 1365.485 2796.150 ;
        RECT 1366.325 2795.720 1375.145 2796.150 ;
        RECT 1375.985 2795.720 1384.805 2796.150 ;
        RECT 1385.645 2795.720 1394.465 2796.150 ;
        RECT 1395.305 2795.720 1404.125 2796.150 ;
        RECT 1404.965 2795.720 1413.785 2796.150 ;
        RECT 1414.625 2795.720 1423.445 2796.150 ;
        RECT 1424.285 2795.720 1433.105 2796.150 ;
        RECT 1433.945 2795.720 1442.765 2796.150 ;
        RECT 1443.605 2795.720 1452.425 2796.150 ;
        RECT 1453.265 2795.720 1462.085 2796.150 ;
        RECT 1462.925 2795.720 1471.745 2796.150 ;
        RECT 1472.585 2795.720 1481.405 2796.150 ;
        RECT 1482.245 2795.720 1491.065 2796.150 ;
        RECT 1491.905 2795.720 1500.725 2796.150 ;
        RECT 1501.565 2795.720 1510.385 2796.150 ;
        RECT 1511.225 2795.720 1520.045 2796.150 ;
        RECT 1520.885 2795.720 1529.245 2796.150 ;
        RECT 1530.085 2795.720 1538.905 2796.150 ;
        RECT 1539.745 2795.720 1548.565 2796.150 ;
        RECT 1549.405 2795.720 1558.225 2796.150 ;
        RECT 1559.065 2795.720 1567.885 2796.150 ;
        RECT 1568.725 2795.720 1577.545 2796.150 ;
        RECT 1578.385 2795.720 1587.205 2796.150 ;
        RECT 1588.045 2795.720 1596.865 2796.150 ;
        RECT 1597.705 2795.720 1606.525 2796.150 ;
        RECT 1607.365 2795.720 1616.185 2796.150 ;
        RECT 1617.025 2795.720 1625.845 2796.150 ;
        RECT 1626.685 2795.720 1635.505 2796.150 ;
        RECT 1636.345 2795.720 1645.165 2796.150 ;
        RECT 1646.005 2795.720 1654.825 2796.150 ;
        RECT 1655.665 2795.720 1664.485 2796.150 ;
        RECT 1665.325 2795.720 1674.145 2796.150 ;
        RECT 1674.985 2795.720 1683.805 2796.150 ;
        RECT 1684.645 2795.720 1693.465 2796.150 ;
        RECT 1694.305 2795.720 1703.125 2796.150 ;
        RECT 1703.965 2795.720 1712.785 2796.150 ;
        RECT 1713.625 2795.720 1722.445 2796.150 ;
        RECT 1723.285 2795.720 1732.105 2796.150 ;
        RECT 1732.945 2795.720 1741.765 2796.150 ;
        RECT 1742.605 2795.720 1751.425 2796.150 ;
        RECT 1752.265 2795.720 1761.085 2796.150 ;
        RECT 1761.925 2795.720 1770.745 2796.150 ;
        RECT 1771.585 2795.720 1780.405 2796.150 ;
        RECT 1781.245 2795.720 1790.065 2796.150 ;
        RECT 1790.905 2795.720 1799.725 2796.150 ;
        RECT 1800.565 2795.720 1809.385 2796.150 ;
        RECT 1810.225 2795.720 1819.045 2796.150 ;
        RECT 1819.885 2795.720 1828.705 2796.150 ;
        RECT 1829.545 2795.720 1838.365 2796.150 ;
        RECT 1839.205 2795.720 1848.025 2796.150 ;
        RECT 1848.865 2795.720 1857.685 2796.150 ;
        RECT 1858.525 2795.720 1867.345 2796.150 ;
        RECT 1868.185 2795.720 1877.005 2796.150 ;
        RECT 1877.845 2795.720 1886.665 2796.150 ;
        RECT 1887.505 2795.720 1895.865 2796.150 ;
        RECT 1896.705 2795.720 1905.525 2796.150 ;
        RECT 1906.365 2795.720 1915.185 2796.150 ;
        RECT 1916.025 2795.720 1924.845 2796.150 ;
        RECT 1925.685 2795.720 1934.505 2796.150 ;
        RECT 1935.345 2795.720 1944.165 2796.150 ;
        RECT 1945.005 2795.720 1953.825 2796.150 ;
        RECT 1954.665 2795.720 1963.485 2796.150 ;
        RECT 1964.325 2795.720 1973.145 2796.150 ;
        RECT 1973.985 2795.720 1982.805 2796.150 ;
        RECT 1983.645 2795.720 1992.465 2796.150 ;
        RECT 1993.305 2795.720 2002.125 2796.150 ;
        RECT 2002.965 2795.720 2011.785 2796.150 ;
        RECT 2012.625 2795.720 2021.445 2796.150 ;
        RECT 2022.285 2795.720 2031.105 2796.150 ;
        RECT 2031.945 2795.720 2040.765 2796.150 ;
        RECT 2041.605 2795.720 2050.425 2796.150 ;
        RECT 2051.265 2795.720 2060.085 2796.150 ;
        RECT 2060.925 2795.720 2069.745 2796.150 ;
        RECT 2070.585 2795.720 2079.405 2796.150 ;
        RECT 2080.245 2795.720 2089.065 2796.150 ;
        RECT 2089.905 2795.720 2098.725 2796.150 ;
        RECT 2099.565 2795.720 2108.385 2796.150 ;
        RECT 2109.225 2795.720 2118.045 2796.150 ;
        RECT 2118.885 2795.720 2127.705 2796.150 ;
        RECT 2128.545 2795.720 2137.365 2796.150 ;
        RECT 2138.205 2795.720 2147.025 2796.150 ;
        RECT 2147.865 2795.720 2156.685 2796.150 ;
        RECT 2157.525 2795.720 2166.345 2796.150 ;
        RECT 2167.185 2795.720 2176.005 2796.150 ;
        RECT 2176.845 2795.720 2185.665 2796.150 ;
        RECT 2186.505 2795.720 2195.325 2796.150 ;
        RECT 2196.165 2795.720 2204.985 2796.150 ;
        RECT 2205.825 2795.720 2214.645 2796.150 ;
        RECT 2215.485 2795.720 2224.305 2796.150 ;
        RECT 2225.145 2795.720 2233.965 2796.150 ;
        RECT 2234.805 2795.720 2243.625 2796.150 ;
        RECT 2244.465 2795.720 2247.855 2796.150 ;
        RECT 1150.025 1704.280 2247.855 2795.720 ;
        RECT 1150.585 1704.000 1151.585 1704.280 ;
        RECT 1152.425 1704.000 1153.885 1704.280 ;
        RECT 1154.725 1704.000 1156.185 1704.280 ;
        RECT 1157.025 1704.000 1158.485 1704.280 ;
        RECT 1159.325 1704.000 1160.785 1704.280 ;
        RECT 1161.625 1704.000 1163.085 1704.280 ;
        RECT 1163.925 1704.000 1165.385 1704.280 ;
        RECT 1166.225 1704.000 1167.685 1704.280 ;
        RECT 1168.525 1704.000 1169.525 1704.280 ;
        RECT 1170.365 1704.000 1171.825 1704.280 ;
        RECT 1172.665 1704.000 1174.125 1704.280 ;
        RECT 1174.965 1704.000 1176.425 1704.280 ;
        RECT 1177.265 1704.000 1178.725 1704.280 ;
        RECT 1179.565 1704.000 1181.025 1704.280 ;
        RECT 1181.865 1704.000 1183.325 1704.280 ;
        RECT 1184.165 1704.000 1185.625 1704.280 ;
        RECT 1186.465 1704.000 1187.465 1704.280 ;
        RECT 1188.305 1704.000 1189.765 1704.280 ;
        RECT 1190.605 1704.000 1192.065 1704.280 ;
        RECT 1192.905 1704.000 1194.365 1704.280 ;
        RECT 1195.205 1704.000 1196.665 1704.280 ;
        RECT 1197.505 1704.000 1198.965 1704.280 ;
        RECT 1199.805 1704.000 1201.265 1704.280 ;
        RECT 1202.105 1704.000 1203.565 1704.280 ;
        RECT 1204.405 1704.000 1205.405 1704.280 ;
        RECT 1206.245 1704.000 1207.705 1704.280 ;
        RECT 1208.545 1704.000 1210.005 1704.280 ;
        RECT 1210.845 1704.000 1212.305 1704.280 ;
        RECT 1213.145 1704.000 1214.605 1704.280 ;
        RECT 1215.445 1704.000 1216.905 1704.280 ;
        RECT 1217.745 1704.000 1219.205 1704.280 ;
        RECT 1220.045 1704.000 1221.505 1704.280 ;
        RECT 1222.345 1704.000 1223.805 1704.280 ;
        RECT 1224.645 1704.000 1225.645 1704.280 ;
        RECT 1226.485 1704.000 1227.945 1704.280 ;
        RECT 1228.785 1704.000 1230.245 1704.280 ;
        RECT 1231.085 1704.000 1232.545 1704.280 ;
        RECT 1233.385 1704.000 1234.845 1704.280 ;
        RECT 1235.685 1704.000 1237.145 1704.280 ;
        RECT 1237.985 1704.000 1239.445 1704.280 ;
        RECT 1240.285 1704.000 1241.745 1704.280 ;
        RECT 1242.585 1704.000 1243.585 1704.280 ;
        RECT 1244.425 1704.000 1245.885 1704.280 ;
        RECT 1246.725 1704.000 1248.185 1704.280 ;
        RECT 1249.025 1704.000 1250.485 1704.280 ;
        RECT 1251.325 1704.000 1252.785 1704.280 ;
        RECT 1253.625 1704.000 1255.085 1704.280 ;
        RECT 1255.925 1704.000 1257.385 1704.280 ;
        RECT 1258.225 1704.000 1259.685 1704.280 ;
        RECT 1260.525 1704.000 1261.525 1704.280 ;
        RECT 1262.365 1704.000 1263.825 1704.280 ;
        RECT 1264.665 1704.000 1266.125 1704.280 ;
        RECT 1266.965 1704.000 1268.425 1704.280 ;
        RECT 1269.265 1704.000 1270.725 1704.280 ;
        RECT 1271.565 1704.000 1273.025 1704.280 ;
        RECT 1273.865 1704.000 1275.325 1704.280 ;
        RECT 1276.165 1704.000 1277.625 1704.280 ;
        RECT 1278.465 1704.000 1279.925 1704.280 ;
        RECT 1280.765 1704.000 1281.765 1704.280 ;
        RECT 1282.605 1704.000 1284.065 1704.280 ;
        RECT 1284.905 1704.000 1286.365 1704.280 ;
        RECT 1287.205 1704.000 1288.665 1704.280 ;
        RECT 1289.505 1704.000 1290.965 1704.280 ;
        RECT 1291.805 1704.000 1293.265 1704.280 ;
        RECT 1294.105 1704.000 1295.565 1704.280 ;
        RECT 1296.405 1704.000 1297.865 1704.280 ;
        RECT 1298.705 1704.000 1299.705 1704.280 ;
        RECT 1300.545 1704.000 1302.005 1704.280 ;
        RECT 1302.845 1704.000 1304.305 1704.280 ;
        RECT 1305.145 1704.000 1306.605 1704.280 ;
        RECT 1307.445 1704.000 1308.905 1704.280 ;
        RECT 1309.745 1704.000 1311.205 1704.280 ;
        RECT 1312.045 1704.000 1313.505 1704.280 ;
        RECT 1314.345 1704.000 1315.805 1704.280 ;
        RECT 1316.645 1704.000 1317.645 1704.280 ;
        RECT 1318.485 1704.000 1319.945 1704.280 ;
        RECT 1320.785 1704.000 1322.245 1704.280 ;
        RECT 1323.085 1704.000 1324.545 1704.280 ;
        RECT 1325.385 1704.000 1326.845 1704.280 ;
        RECT 1327.685 1704.000 1329.145 1704.280 ;
        RECT 1329.985 1704.000 1331.445 1704.280 ;
        RECT 1332.285 1704.000 1333.745 1704.280 ;
        RECT 1334.585 1704.000 1336.045 1704.280 ;
        RECT 1336.885 1704.000 1337.885 1704.280 ;
        RECT 1338.725 1704.000 1340.185 1704.280 ;
        RECT 1341.025 1704.000 1342.485 1704.280 ;
        RECT 1343.325 1704.000 1344.785 1704.280 ;
        RECT 1345.625 1704.000 1347.085 1704.280 ;
        RECT 1347.925 1704.000 1349.385 1704.280 ;
        RECT 1350.225 1704.000 1351.685 1704.280 ;
        RECT 1352.525 1704.000 1353.985 1704.280 ;
        RECT 1354.825 1704.000 1355.825 1704.280 ;
        RECT 1356.665 1704.000 1358.125 1704.280 ;
        RECT 1358.965 1704.000 1360.425 1704.280 ;
        RECT 1361.265 1704.000 1362.725 1704.280 ;
        RECT 1363.565 1704.000 1365.025 1704.280 ;
        RECT 1365.865 1704.000 1367.325 1704.280 ;
        RECT 1368.165 1704.000 1369.625 1704.280 ;
        RECT 1370.465 1704.000 1371.925 1704.280 ;
        RECT 1372.765 1704.000 1373.765 1704.280 ;
        RECT 1374.605 1704.000 1376.065 1704.280 ;
        RECT 1376.905 1704.000 1378.365 1704.280 ;
        RECT 1379.205 1704.000 1380.665 1704.280 ;
        RECT 1381.505 1704.000 1382.965 1704.280 ;
        RECT 1383.805 1704.000 1385.265 1704.280 ;
        RECT 1386.105 1704.000 1387.565 1704.280 ;
        RECT 1388.405 1704.000 1389.865 1704.280 ;
        RECT 1390.705 1704.000 1391.705 1704.280 ;
        RECT 1392.545 1704.000 1394.005 1704.280 ;
        RECT 1394.845 1704.000 1396.305 1704.280 ;
        RECT 1397.145 1704.000 1398.605 1704.280 ;
        RECT 1399.445 1704.000 1400.905 1704.280 ;
        RECT 1401.745 1704.000 1403.205 1704.280 ;
        RECT 1404.045 1704.000 1405.505 1704.280 ;
        RECT 1406.345 1704.000 1407.805 1704.280 ;
        RECT 1408.645 1704.000 1410.105 1704.280 ;
        RECT 1410.945 1704.000 1411.945 1704.280 ;
        RECT 1412.785 1704.000 1414.245 1704.280 ;
        RECT 1415.085 1704.000 1416.545 1704.280 ;
        RECT 1417.385 1704.000 1418.845 1704.280 ;
        RECT 1419.685 1704.000 1421.145 1704.280 ;
        RECT 1421.985 1704.000 1423.445 1704.280 ;
        RECT 1424.285 1704.000 1425.745 1704.280 ;
        RECT 1426.585 1704.000 1428.045 1704.280 ;
        RECT 1428.885 1704.000 1429.885 1704.280 ;
        RECT 1430.725 1704.000 1432.185 1704.280 ;
        RECT 1433.025 1704.000 1434.485 1704.280 ;
        RECT 1435.325 1704.000 1436.785 1704.280 ;
        RECT 1437.625 1704.000 1439.085 1704.280 ;
        RECT 1439.925 1704.000 1441.385 1704.280 ;
        RECT 1442.225 1704.000 1443.685 1704.280 ;
        RECT 1444.525 1704.000 1445.985 1704.280 ;
        RECT 1446.825 1704.000 1447.825 1704.280 ;
        RECT 1448.665 1704.000 1450.125 1704.280 ;
        RECT 1450.965 1704.000 1452.425 1704.280 ;
        RECT 1453.265 1704.000 1454.725 1704.280 ;
        RECT 1455.565 1704.000 1457.025 1704.280 ;
        RECT 1457.865 1704.000 1459.325 1704.280 ;
        RECT 1460.165 1704.000 1461.625 1704.280 ;
        RECT 1462.465 1704.000 1463.925 1704.280 ;
        RECT 1464.765 1704.000 1466.225 1704.280 ;
        RECT 1467.065 1704.000 1468.065 1704.280 ;
        RECT 1468.905 1704.000 1470.365 1704.280 ;
        RECT 1471.205 1704.000 1472.665 1704.280 ;
        RECT 1473.505 1704.000 1474.965 1704.280 ;
        RECT 1475.805 1704.000 1477.265 1704.280 ;
        RECT 1478.105 1704.000 1479.565 1704.280 ;
        RECT 1480.405 1704.000 1481.865 1704.280 ;
        RECT 1482.705 1704.000 1484.165 1704.280 ;
        RECT 1485.005 1704.000 1486.005 1704.280 ;
        RECT 1486.845 1704.000 1488.305 1704.280 ;
        RECT 1489.145 1704.000 1490.605 1704.280 ;
        RECT 1491.445 1704.000 1492.905 1704.280 ;
        RECT 1493.745 1704.000 1495.205 1704.280 ;
        RECT 1496.045 1704.000 1497.505 1704.280 ;
        RECT 1498.345 1704.000 1499.805 1704.280 ;
        RECT 1500.645 1704.000 1502.105 1704.280 ;
        RECT 1502.945 1704.000 1503.945 1704.280 ;
        RECT 1504.785 1704.000 1506.245 1704.280 ;
        RECT 1507.085 1704.000 1508.545 1704.280 ;
        RECT 1509.385 1704.000 1510.845 1704.280 ;
        RECT 1511.685 1704.000 1513.145 1704.280 ;
        RECT 1513.985 1704.000 1515.445 1704.280 ;
        RECT 1516.285 1704.000 1517.745 1704.280 ;
        RECT 1518.585 1704.000 1520.045 1704.280 ;
        RECT 1520.885 1704.000 1522.345 1704.280 ;
        RECT 1523.185 1704.000 1524.185 1704.280 ;
        RECT 1525.025 1704.000 1526.485 1704.280 ;
        RECT 1527.325 1704.000 1528.785 1704.280 ;
        RECT 1529.625 1704.000 1531.085 1704.280 ;
        RECT 1531.925 1704.000 1533.385 1704.280 ;
        RECT 1534.225 1704.000 1535.685 1704.280 ;
        RECT 1536.525 1704.000 1537.985 1704.280 ;
        RECT 1538.825 1704.000 1540.285 1704.280 ;
        RECT 1541.125 1704.000 1542.125 1704.280 ;
        RECT 1542.965 1704.000 1544.425 1704.280 ;
        RECT 1545.265 1704.000 1546.725 1704.280 ;
        RECT 1547.565 1704.000 1549.025 1704.280 ;
        RECT 1549.865 1704.000 1551.325 1704.280 ;
        RECT 1552.165 1704.000 1553.625 1704.280 ;
        RECT 1554.465 1704.000 1555.925 1704.280 ;
        RECT 1556.765 1704.000 1558.225 1704.280 ;
        RECT 1559.065 1704.000 1560.065 1704.280 ;
        RECT 1560.905 1704.000 1562.365 1704.280 ;
        RECT 1563.205 1704.000 1564.665 1704.280 ;
        RECT 1565.505 1704.000 1566.965 1704.280 ;
        RECT 1567.805 1704.000 1569.265 1704.280 ;
        RECT 1570.105 1704.000 1571.565 1704.280 ;
        RECT 1572.405 1704.000 1573.865 1704.280 ;
        RECT 1574.705 1704.000 1576.165 1704.280 ;
        RECT 1577.005 1704.000 1578.465 1704.280 ;
        RECT 1579.305 1704.000 1580.305 1704.280 ;
        RECT 1581.145 1704.000 1582.605 1704.280 ;
        RECT 1583.445 1704.000 1584.905 1704.280 ;
        RECT 1585.745 1704.000 1587.205 1704.280 ;
        RECT 1588.045 1704.000 1589.505 1704.280 ;
        RECT 1590.345 1704.000 1591.805 1704.280 ;
        RECT 1592.645 1704.000 1594.105 1704.280 ;
        RECT 1594.945 1704.000 1596.405 1704.280 ;
        RECT 1597.245 1704.000 1598.245 1704.280 ;
        RECT 1599.085 1704.000 1600.545 1704.280 ;
        RECT 1601.385 1704.000 1602.845 1704.280 ;
        RECT 1603.685 1704.000 1605.145 1704.280 ;
        RECT 1605.985 1704.000 1607.445 1704.280 ;
        RECT 1608.285 1704.000 1609.745 1704.280 ;
        RECT 1610.585 1704.000 1612.045 1704.280 ;
        RECT 1612.885 1704.000 1614.345 1704.280 ;
        RECT 1615.185 1704.000 1616.185 1704.280 ;
        RECT 1617.025 1704.000 1618.485 1704.280 ;
        RECT 1619.325 1704.000 1620.785 1704.280 ;
        RECT 1621.625 1704.000 1623.085 1704.280 ;
        RECT 1623.925 1704.000 1625.385 1704.280 ;
        RECT 1626.225 1704.000 1627.685 1704.280 ;
        RECT 1628.525 1704.000 1629.985 1704.280 ;
        RECT 1630.825 1704.000 1632.285 1704.280 ;
        RECT 1633.125 1704.000 1634.125 1704.280 ;
        RECT 1634.965 1704.000 1636.425 1704.280 ;
        RECT 1637.265 1704.000 1638.725 1704.280 ;
        RECT 1639.565 1704.000 1641.025 1704.280 ;
        RECT 1641.865 1704.000 1643.325 1704.280 ;
        RECT 1644.165 1704.000 1645.625 1704.280 ;
        RECT 1646.465 1704.000 1647.925 1704.280 ;
        RECT 1648.765 1704.000 1650.225 1704.280 ;
        RECT 1651.065 1704.000 1652.525 1704.280 ;
        RECT 1653.365 1704.000 1654.365 1704.280 ;
        RECT 1655.205 1704.000 1656.665 1704.280 ;
        RECT 1657.505 1704.000 1658.965 1704.280 ;
        RECT 1659.805 1704.000 1661.265 1704.280 ;
        RECT 1662.105 1704.000 1663.565 1704.280 ;
        RECT 1664.405 1704.000 1665.865 1704.280 ;
        RECT 1666.705 1704.000 1668.165 1704.280 ;
        RECT 1669.005 1704.000 1670.465 1704.280 ;
        RECT 1671.305 1704.000 1672.305 1704.280 ;
        RECT 1673.145 1704.000 1674.605 1704.280 ;
        RECT 1675.445 1704.000 1676.905 1704.280 ;
        RECT 1677.745 1704.000 1679.205 1704.280 ;
        RECT 1680.045 1704.000 1681.505 1704.280 ;
        RECT 1682.345 1704.000 1683.805 1704.280 ;
        RECT 1684.645 1704.000 1686.105 1704.280 ;
        RECT 1686.945 1704.000 1688.405 1704.280 ;
        RECT 1689.245 1704.000 1690.245 1704.280 ;
        RECT 1691.085 1704.000 1692.545 1704.280 ;
        RECT 1693.385 1704.000 1694.845 1704.280 ;
        RECT 1695.685 1704.000 1697.145 1704.280 ;
        RECT 1697.985 1704.000 1699.445 1704.280 ;
        RECT 1700.285 1704.000 1701.745 1704.280 ;
        RECT 1702.585 1704.000 1704.045 1704.280 ;
        RECT 1704.885 1704.000 1706.345 1704.280 ;
        RECT 1707.185 1704.000 1708.645 1704.280 ;
        RECT 1709.485 1704.000 1710.485 1704.280 ;
        RECT 1711.325 1704.000 1712.785 1704.280 ;
        RECT 1713.625 1704.000 1715.085 1704.280 ;
        RECT 1715.925 1704.000 1717.385 1704.280 ;
        RECT 1718.225 1704.000 1719.685 1704.280 ;
        RECT 1720.525 1704.000 1721.985 1704.280 ;
        RECT 1722.825 1704.000 1724.285 1704.280 ;
        RECT 1725.125 1704.000 1726.585 1704.280 ;
        RECT 1727.425 1704.000 1728.425 1704.280 ;
        RECT 1729.265 1704.000 1730.725 1704.280 ;
        RECT 1731.565 1704.000 1733.025 1704.280 ;
        RECT 1733.865 1704.000 1735.325 1704.280 ;
        RECT 1736.165 1704.000 1737.625 1704.280 ;
        RECT 1738.465 1704.000 1739.925 1704.280 ;
        RECT 1740.765 1704.000 1742.225 1704.280 ;
        RECT 1743.065 1704.000 1744.525 1704.280 ;
        RECT 1745.365 1704.000 1746.365 1704.280 ;
        RECT 1747.205 1704.000 1748.665 1704.280 ;
        RECT 1749.505 1704.000 1750.965 1704.280 ;
        RECT 1751.805 1704.000 1753.265 1704.280 ;
        RECT 1754.105 1704.000 1755.565 1704.280 ;
        RECT 1756.405 1704.000 1757.865 1704.280 ;
        RECT 1758.705 1704.000 1760.165 1704.280 ;
        RECT 1761.005 1704.000 1762.465 1704.280 ;
        RECT 1763.305 1704.000 1764.765 1704.280 ;
        RECT 1765.605 1704.000 1766.605 1704.280 ;
        RECT 1767.445 1704.000 1768.905 1704.280 ;
        RECT 1769.745 1704.000 1771.205 1704.280 ;
        RECT 1772.045 1704.000 1773.505 1704.280 ;
        RECT 1774.345 1704.000 1775.805 1704.280 ;
        RECT 1776.645 1704.000 1778.105 1704.280 ;
        RECT 1778.945 1704.000 1780.405 1704.280 ;
        RECT 1781.245 1704.000 1782.705 1704.280 ;
        RECT 1783.545 1704.000 1784.545 1704.280 ;
        RECT 1785.385 1704.000 1786.845 1704.280 ;
        RECT 1787.685 1704.000 1789.145 1704.280 ;
        RECT 1789.985 1704.000 1791.445 1704.280 ;
        RECT 1792.285 1704.000 1793.745 1704.280 ;
        RECT 1794.585 1704.000 1796.045 1704.280 ;
        RECT 1796.885 1704.000 1798.345 1704.280 ;
        RECT 1799.185 1704.000 1800.645 1704.280 ;
        RECT 1801.485 1704.000 1802.485 1704.280 ;
        RECT 1803.325 1704.000 1804.785 1704.280 ;
        RECT 1805.625 1704.000 1807.085 1704.280 ;
        RECT 1807.925 1704.000 1809.385 1704.280 ;
        RECT 1810.225 1704.000 1811.685 1704.280 ;
        RECT 1812.525 1704.000 1813.985 1704.280 ;
        RECT 1814.825 1704.000 1816.285 1704.280 ;
        RECT 1817.125 1704.000 1818.585 1704.280 ;
        RECT 1819.425 1704.000 1820.425 1704.280 ;
        RECT 1821.265 1704.000 1822.725 1704.280 ;
        RECT 1823.565 1704.000 1825.025 1704.280 ;
        RECT 1825.865 1704.000 1827.325 1704.280 ;
        RECT 1828.165 1704.000 1829.625 1704.280 ;
        RECT 1830.465 1704.000 1831.925 1704.280 ;
        RECT 1832.765 1704.000 1834.225 1704.280 ;
        RECT 1835.065 1704.000 1836.525 1704.280 ;
        RECT 1837.365 1704.000 1838.825 1704.280 ;
        RECT 1839.665 1704.000 1840.665 1704.280 ;
        RECT 1841.505 1704.000 1842.965 1704.280 ;
        RECT 1843.805 1704.000 1845.265 1704.280 ;
        RECT 1846.105 1704.000 1847.565 1704.280 ;
        RECT 1848.405 1704.000 1849.865 1704.280 ;
        RECT 1850.705 1704.000 1852.165 1704.280 ;
        RECT 1853.005 1704.000 1854.465 1704.280 ;
        RECT 1855.305 1704.000 1856.765 1704.280 ;
        RECT 1857.605 1704.000 1858.605 1704.280 ;
        RECT 1859.445 1704.000 1860.905 1704.280 ;
        RECT 1861.745 1704.000 1863.205 1704.280 ;
        RECT 1864.045 1704.000 1865.505 1704.280 ;
        RECT 1866.345 1704.000 1867.805 1704.280 ;
        RECT 1868.645 1704.000 1870.105 1704.280 ;
        RECT 1870.945 1704.000 1872.405 1704.280 ;
        RECT 1873.245 1704.000 1874.705 1704.280 ;
        RECT 1875.545 1704.000 1876.545 1704.280 ;
        RECT 1877.385 1704.000 1878.845 1704.280 ;
        RECT 1879.685 1704.000 1881.145 1704.280 ;
        RECT 1881.985 1704.000 1883.445 1704.280 ;
        RECT 1884.285 1704.000 1885.745 1704.280 ;
        RECT 1886.585 1704.000 1888.045 1704.280 ;
        RECT 1888.885 1704.000 1890.345 1704.280 ;
        RECT 1891.185 1704.000 1892.645 1704.280 ;
        RECT 1893.485 1704.000 1894.945 1704.280 ;
        RECT 1895.785 1704.000 1896.785 1704.280 ;
        RECT 1897.625 1704.000 1899.085 1704.280 ;
        RECT 1899.925 1704.000 1901.385 1704.280 ;
        RECT 1902.225 1704.000 1903.685 1704.280 ;
        RECT 1904.525 1704.000 1905.985 1704.280 ;
        RECT 1906.825 1704.000 1908.285 1704.280 ;
        RECT 1909.125 1704.000 1910.585 1704.280 ;
        RECT 1911.425 1704.000 1912.885 1704.280 ;
        RECT 1913.725 1704.000 1914.725 1704.280 ;
        RECT 1915.565 1704.000 1917.025 1704.280 ;
        RECT 1917.865 1704.000 1919.325 1704.280 ;
        RECT 1920.165 1704.000 1921.625 1704.280 ;
        RECT 1922.465 1704.000 1923.925 1704.280 ;
        RECT 1924.765 1704.000 1926.225 1704.280 ;
        RECT 1927.065 1704.000 1928.525 1704.280 ;
        RECT 1929.365 1704.000 1930.825 1704.280 ;
        RECT 1931.665 1704.000 1932.665 1704.280 ;
        RECT 1933.505 1704.000 1934.965 1704.280 ;
        RECT 1935.805 1704.000 1937.265 1704.280 ;
        RECT 1938.105 1704.000 1939.565 1704.280 ;
        RECT 1940.405 1704.000 1941.865 1704.280 ;
        RECT 1942.705 1704.000 1944.165 1704.280 ;
        RECT 1945.005 1704.000 1946.465 1704.280 ;
        RECT 1947.305 1704.000 1948.765 1704.280 ;
        RECT 1949.605 1704.000 1951.065 1704.280 ;
        RECT 1951.905 1704.000 1952.905 1704.280 ;
        RECT 1953.745 1704.000 1955.205 1704.280 ;
        RECT 1956.045 1704.000 1957.505 1704.280 ;
        RECT 1958.345 1704.000 1959.805 1704.280 ;
        RECT 1960.645 1704.000 1962.105 1704.280 ;
        RECT 1962.945 1704.000 1964.405 1704.280 ;
        RECT 1965.245 1704.000 1966.705 1704.280 ;
        RECT 1967.545 1704.000 1969.005 1704.280 ;
        RECT 1969.845 1704.000 1970.845 1704.280 ;
        RECT 1971.685 1704.000 1973.145 1704.280 ;
        RECT 1973.985 1704.000 1975.445 1704.280 ;
        RECT 1976.285 1704.000 1977.745 1704.280 ;
        RECT 1978.585 1704.000 1980.045 1704.280 ;
        RECT 1980.885 1704.000 1982.345 1704.280 ;
        RECT 1983.185 1704.000 1984.645 1704.280 ;
        RECT 1985.485 1704.000 1986.945 1704.280 ;
        RECT 1987.785 1704.000 1988.785 1704.280 ;
        RECT 1989.625 1704.000 1991.085 1704.280 ;
        RECT 1991.925 1704.000 1993.385 1704.280 ;
        RECT 1994.225 1704.000 1995.685 1704.280 ;
        RECT 1996.525 1704.000 1997.985 1704.280 ;
        RECT 1998.825 1704.000 2000.285 1704.280 ;
        RECT 2001.125 1704.000 2002.585 1704.280 ;
        RECT 2003.425 1704.000 2004.885 1704.280 ;
        RECT 2005.725 1704.000 2007.185 1704.280 ;
        RECT 2008.025 1704.000 2009.025 1704.280 ;
        RECT 2009.865 1704.000 2011.325 1704.280 ;
        RECT 2012.165 1704.000 2013.625 1704.280 ;
        RECT 2014.465 1704.000 2015.925 1704.280 ;
        RECT 2016.765 1704.000 2018.225 1704.280 ;
        RECT 2019.065 1704.000 2020.525 1704.280 ;
        RECT 2021.365 1704.000 2022.825 1704.280 ;
        RECT 2023.665 1704.000 2025.125 1704.280 ;
        RECT 2025.965 1704.000 2026.965 1704.280 ;
        RECT 2027.805 1704.000 2029.265 1704.280 ;
        RECT 2030.105 1704.000 2031.565 1704.280 ;
        RECT 2032.405 1704.000 2033.865 1704.280 ;
        RECT 2034.705 1704.000 2036.165 1704.280 ;
        RECT 2037.005 1704.000 2038.465 1704.280 ;
        RECT 2039.305 1704.000 2040.765 1704.280 ;
        RECT 2041.605 1704.000 2043.065 1704.280 ;
        RECT 2043.905 1704.000 2044.905 1704.280 ;
        RECT 2045.745 1704.000 2047.205 1704.280 ;
        RECT 2048.045 1704.000 2049.505 1704.280 ;
        RECT 2050.345 1704.000 2051.805 1704.280 ;
        RECT 2052.645 1704.000 2054.105 1704.280 ;
        RECT 2054.945 1704.000 2056.405 1704.280 ;
        RECT 2057.245 1704.000 2058.705 1704.280 ;
        RECT 2059.545 1704.000 2061.005 1704.280 ;
        RECT 2061.845 1704.000 2062.845 1704.280 ;
        RECT 2063.685 1704.000 2065.145 1704.280 ;
        RECT 2065.985 1704.000 2067.445 1704.280 ;
        RECT 2068.285 1704.000 2069.745 1704.280 ;
        RECT 2070.585 1704.000 2072.045 1704.280 ;
        RECT 2072.885 1704.000 2074.345 1704.280 ;
        RECT 2075.185 1704.000 2076.645 1704.280 ;
        RECT 2077.485 1704.000 2078.945 1704.280 ;
        RECT 2079.785 1704.000 2081.245 1704.280 ;
        RECT 2082.085 1704.000 2083.085 1704.280 ;
        RECT 2083.925 1704.000 2085.385 1704.280 ;
        RECT 2086.225 1704.000 2087.685 1704.280 ;
        RECT 2088.525 1704.000 2089.985 1704.280 ;
        RECT 2090.825 1704.000 2092.285 1704.280 ;
        RECT 2093.125 1704.000 2094.585 1704.280 ;
        RECT 2095.425 1704.000 2096.885 1704.280 ;
        RECT 2097.725 1704.000 2099.185 1704.280 ;
        RECT 2100.025 1704.000 2101.025 1704.280 ;
        RECT 2101.865 1704.000 2103.325 1704.280 ;
        RECT 2104.165 1704.000 2105.625 1704.280 ;
        RECT 2106.465 1704.000 2107.925 1704.280 ;
        RECT 2108.765 1704.000 2110.225 1704.280 ;
        RECT 2111.065 1704.000 2112.525 1704.280 ;
        RECT 2113.365 1704.000 2114.825 1704.280 ;
        RECT 2115.665 1704.000 2117.125 1704.280 ;
        RECT 2117.965 1704.000 2118.965 1704.280 ;
        RECT 2119.805 1704.000 2121.265 1704.280 ;
        RECT 2122.105 1704.000 2123.565 1704.280 ;
        RECT 2124.405 1704.000 2125.865 1704.280 ;
        RECT 2126.705 1704.000 2128.165 1704.280 ;
        RECT 2129.005 1704.000 2130.465 1704.280 ;
        RECT 2131.305 1704.000 2132.765 1704.280 ;
        RECT 2133.605 1704.000 2135.065 1704.280 ;
        RECT 2135.905 1704.000 2137.365 1704.280 ;
        RECT 2138.205 1704.000 2139.205 1704.280 ;
        RECT 2140.045 1704.000 2141.505 1704.280 ;
        RECT 2142.345 1704.000 2143.805 1704.280 ;
        RECT 2144.645 1704.000 2146.105 1704.280 ;
        RECT 2146.945 1704.000 2148.405 1704.280 ;
        RECT 2149.245 1704.000 2150.705 1704.280 ;
        RECT 2151.545 1704.000 2153.005 1704.280 ;
        RECT 2153.845 1704.000 2155.305 1704.280 ;
        RECT 2156.145 1704.000 2157.145 1704.280 ;
        RECT 2157.985 1704.000 2159.445 1704.280 ;
        RECT 2160.285 1704.000 2161.745 1704.280 ;
        RECT 2162.585 1704.000 2164.045 1704.280 ;
        RECT 2164.885 1704.000 2166.345 1704.280 ;
        RECT 2167.185 1704.000 2168.645 1704.280 ;
        RECT 2169.485 1704.000 2170.945 1704.280 ;
        RECT 2171.785 1704.000 2173.245 1704.280 ;
        RECT 2174.085 1704.000 2175.085 1704.280 ;
        RECT 2175.925 1704.000 2177.385 1704.280 ;
        RECT 2178.225 1704.000 2179.685 1704.280 ;
        RECT 2180.525 1704.000 2181.985 1704.280 ;
        RECT 2182.825 1704.000 2184.285 1704.280 ;
        RECT 2185.125 1704.000 2186.585 1704.280 ;
        RECT 2187.425 1704.000 2188.885 1704.280 ;
        RECT 2189.725 1704.000 2191.185 1704.280 ;
        RECT 2192.025 1704.000 2193.485 1704.280 ;
        RECT 2194.325 1704.000 2195.325 1704.280 ;
        RECT 2196.165 1704.000 2197.625 1704.280 ;
        RECT 2198.465 1704.000 2199.925 1704.280 ;
        RECT 2200.765 1704.000 2202.225 1704.280 ;
        RECT 2203.065 1704.000 2204.525 1704.280 ;
        RECT 2205.365 1704.000 2206.825 1704.280 ;
        RECT 2207.665 1704.000 2209.125 1704.280 ;
        RECT 2209.965 1704.000 2211.425 1704.280 ;
        RECT 2212.265 1704.000 2213.265 1704.280 ;
        RECT 2214.105 1704.000 2215.565 1704.280 ;
        RECT 2216.405 1704.000 2217.865 1704.280 ;
        RECT 2218.705 1704.000 2220.165 1704.280 ;
        RECT 2221.005 1704.000 2222.465 1704.280 ;
        RECT 2223.305 1704.000 2224.765 1704.280 ;
        RECT 2225.605 1704.000 2227.065 1704.280 ;
        RECT 2227.905 1704.000 2229.365 1704.280 ;
        RECT 2230.205 1704.000 2231.205 1704.280 ;
        RECT 2232.045 1704.000 2233.505 1704.280 ;
        RECT 2234.345 1704.000 2235.805 1704.280 ;
        RECT 2236.645 1704.000 2238.105 1704.280 ;
        RECT 2238.945 1704.000 2240.405 1704.280 ;
        RECT 2241.245 1704.000 2242.705 1704.280 ;
        RECT 2243.545 1704.000 2245.005 1704.280 ;
        RECT 2245.845 1704.000 2247.305 1704.280 ;
      LAYER met3 ;
        RECT 1150.000 1704.255 2229.030 2788.165 ;
      LAYER met4 ;
        RECT 1170.055 1710.640 1171.655 2788.240 ;
      LAYER met4 ;
        RECT 1195.310 1710.640 1210.020 2788.240 ;
        RECT 1213.020 1710.640 1228.020 2788.240 ;
        RECT 1231.020 1710.640 1246.455 2788.240 ;
      LAYER met4 ;
        RECT 1246.855 1710.640 1248.455 2788.240 ;
      LAYER met4 ;
        RECT 1248.855 1710.640 1264.020 2788.240 ;
        RECT 1267.020 1710.640 1282.020 2788.240 ;
        RECT 1285.020 1710.640 1300.020 2788.240 ;
        RECT 1303.020 1710.640 1318.020 2788.240 ;
        RECT 1321.020 1710.640 1354.020 2788.240 ;
        RECT 1357.020 1710.640 1372.020 2788.240 ;
        RECT 1375.020 1710.640 1390.020 2788.240 ;
        RECT 1393.020 1710.640 1408.020 2788.240 ;
        RECT 1411.020 1710.640 1444.020 2788.240 ;
        RECT 1447.020 1710.640 1462.020 2788.240 ;
        RECT 1465.020 1710.640 1480.020 2788.240 ;
        RECT 1483.020 1710.640 1498.020 2788.240 ;
        RECT 1501.020 1710.640 1534.020 2788.240 ;
        RECT 1537.020 1710.640 1552.020 2788.240 ;
        RECT 1555.020 1710.640 1570.020 2788.240 ;
        RECT 1573.020 1710.640 1588.020 2788.240 ;
        RECT 1591.020 1710.640 1624.020 2788.240 ;
        RECT 1627.020 1710.640 1642.020 2788.240 ;
        RECT 1645.020 1710.640 1660.020 2788.240 ;
        RECT 1663.020 1710.640 1678.020 2788.240 ;
        RECT 1681.020 1710.640 1714.020 2788.240 ;
        RECT 1717.020 1710.640 1732.020 2788.240 ;
        RECT 1735.020 1710.640 1750.020 2788.240 ;
        RECT 1753.020 1710.640 1768.020 2788.240 ;
        RECT 1771.020 1710.640 1804.020 2788.240 ;
        RECT 1807.020 1710.640 1822.020 2788.240 ;
        RECT 1825.020 1710.640 1840.020 2788.240 ;
        RECT 1843.020 1710.640 1858.020 2788.240 ;
        RECT 1861.020 1710.640 1894.020 2788.240 ;
        RECT 1897.020 1710.640 1912.020 2788.240 ;
        RECT 1915.020 1710.640 1930.020 2788.240 ;
        RECT 1933.020 1710.640 1948.020 2788.240 ;
        RECT 1951.020 1710.640 1984.020 2788.240 ;
        RECT 1987.020 1710.640 2002.020 2788.240 ;
        RECT 2005.020 1710.640 2020.020 2788.240 ;
        RECT 2023.020 1710.640 2038.020 2788.240 ;
        RECT 2041.020 1710.640 2074.020 2788.240 ;
        RECT 2077.020 1710.640 2092.020 2788.240 ;
        RECT 2095.020 1710.640 2110.020 2788.240 ;
        RECT 2113.020 1710.640 2128.020 2788.240 ;
        RECT 2131.020 1710.640 2164.020 2788.240 ;
        RECT 2167.020 1710.640 2182.020 2788.240 ;
        RECT 2185.020 1710.640 2200.020 2788.240 ;
        RECT 2203.020 1710.640 2218.020 2788.240 ;
  END
END user_project_wrapper
END LIBRARY

