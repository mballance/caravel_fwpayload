VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1197.700 BY 1200.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.160 1196.000 4.440 1200.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.720 1196.000 320.000 1200.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.460 1196.000 351.740 1200.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.740 1196.000 383.020 1200.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.480 1196.000 414.760 1200.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 446.220 1196.000 446.500 1200.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.500 1196.000 477.780 1200.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.240 1196.000 509.520 1200.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.980 1196.000 541.260 1200.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.260 1196.000 572.540 1200.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.000 1196.000 604.280 1200.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.440 1196.000 35.720 1200.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 635.740 1196.000 636.020 1200.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 667.020 1196.000 667.300 1200.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.760 1196.000 699.040 1200.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 730.500 1196.000 730.780 1200.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.780 1196.000 762.060 1200.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.520 1196.000 793.800 1200.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.260 1196.000 825.540 1200.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 856.540 1196.000 856.820 1200.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.280 1196.000 888.560 1200.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.020 1196.000 920.300 1200.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.180 1196.000 67.460 1200.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 951.300 1196.000 951.580 1200.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.040 1196.000 983.320 1200.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.780 1196.000 1015.060 1200.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.060 1196.000 1046.340 1200.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.800 1196.000 1078.080 1200.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.540 1196.000 1109.820 1200.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1140.820 1196.000 1141.100 1200.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1172.560 1196.000 1172.840 1200.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.460 1196.000 98.740 1200.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.200 1196.000 130.480 1200.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.940 1196.000 162.220 1200.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.220 1196.000 193.500 1200.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.960 1196.000 225.240 1200.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.700 1196.000 256.980 1200.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.980 1196.000 288.260 1200.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.280 1196.000 14.560 1200.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 330.300 1196.000 330.580 1200.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.040 1196.000 362.320 1200.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 393.320 1196.000 393.600 1200.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 425.060 1196.000 425.340 1200.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.800 1196.000 457.080 1200.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.080 1196.000 488.360 1200.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.820 1196.000 520.100 1200.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 551.560 1196.000 551.840 1200.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.840 1196.000 583.120 1200.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.580 1196.000 614.860 1200.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.020 1196.000 46.300 1200.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.320 1196.000 646.600 1200.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.600 1196.000 677.880 1200.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.340 1196.000 709.620 1200.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.080 1196.000 741.360 1200.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 772.360 1196.000 772.640 1200.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.100 1196.000 804.380 1200.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.380 1196.000 835.660 1200.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 867.120 1196.000 867.400 1200.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 898.860 1196.000 899.140 1200.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 930.140 1196.000 930.420 1200.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.760 1196.000 78.040 1200.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.880 1196.000 962.160 1200.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 993.620 1196.000 993.900 1200.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.900 1196.000 1025.180 1200.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1056.640 1196.000 1056.920 1200.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1088.380 1196.000 1088.660 1200.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1119.660 1196.000 1119.940 1200.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.400 1196.000 1151.680 1200.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1183.140 1196.000 1183.420 1200.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.040 1196.000 109.320 1200.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.780 1196.000 141.060 1200.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.520 1196.000 172.800 1200.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 203.800 1196.000 204.080 1200.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.540 1196.000 235.820 1200.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.280 1196.000 267.560 1200.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.560 1196.000 298.840 1200.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.860 1196.000 25.140 1200.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.880 1196.000 341.160 1200.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.620 1196.000 372.900 1200.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 403.900 1196.000 404.180 1200.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.640 1196.000 435.920 1200.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.920 1196.000 467.200 1200.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 498.660 1196.000 498.940 1200.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.400 1196.000 530.680 1200.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 561.680 1196.000 561.960 1200.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.420 1196.000 593.700 1200.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 625.160 1196.000 625.440 1200.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.600 1196.000 56.880 1200.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.440 1196.000 656.720 1200.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 688.180 1196.000 688.460 1200.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 719.920 1196.000 720.200 1200.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.200 1196.000 751.480 1200.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 782.940 1196.000 783.220 1200.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.680 1196.000 814.960 1200.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.960 1196.000 846.240 1200.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 877.700 1196.000 877.980 1200.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.440 1196.000 909.720 1200.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 940.720 1196.000 941.000 1200.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.340 1196.000 88.620 1200.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.460 1196.000 972.740 1200.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1004.200 1196.000 1004.480 1200.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1035.480 1196.000 1035.760 1200.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.220 1196.000 1067.500 1200.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1098.960 1196.000 1099.240 1200.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1130.240 1196.000 1130.520 1200.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1161.980 1196.000 1162.260 1200.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1193.720 1196.000 1194.000 1200.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.620 1196.000 119.900 1200.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.360 1196.000 151.640 1200.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.100 1196.000 183.380 1200.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 214.380 1196.000 214.660 1200.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.120 1196.000 246.400 1200.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.860 1196.000 278.140 1200.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.140 1196.000 309.420 1200.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 259.460 0.000 259.740 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.080 0.000 994.360 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.440 0.000 1001.720 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1008.800 0.000 1009.080 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.160 0.000 1016.440 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.520 0.000 1023.800 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.880 0.000 1031.160 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1038.240 0.000 1038.520 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.600 0.000 1045.880 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.960 0.000 1053.240 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.320 0.000 1060.600 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.060 0.000 333.340 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1067.680 0.000 1067.960 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.040 0.000 1075.320 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.400 0.000 1082.680 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1089.760 0.000 1090.040 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.120 0.000 1097.400 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1104.480 0.000 1104.760 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1111.840 0.000 1112.120 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1119.200 0.000 1119.480 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.560 0.000 1126.840 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.920 0.000 1134.200 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.420 0.000 340.700 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1141.280 0.000 1141.560 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1148.640 0.000 1148.920 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.000 0.000 1156.280 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1163.360 0.000 1163.640 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1170.720 0.000 1171.000 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.080 0.000 1178.360 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.440 0.000 1185.720 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1192.800 0.000 1193.080 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.780 0.000 348.060 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 355.140 0.000 355.420 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 362.500 0.000 362.780 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.400 0.000 369.680 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.760 0.000 377.040 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.120 0.000 384.400 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.480 0.000 391.760 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 398.840 0.000 399.120 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.820 0.000 267.100 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.200 0.000 406.480 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.560 0.000 413.840 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.920 0.000 421.200 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 428.280 0.000 428.560 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.640 0.000 435.920 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.000 0.000 443.280 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.360 0.000 450.640 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.720 0.000 458.000 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.080 0.000 465.360 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.440 0.000 472.720 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.180 0.000 274.460 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.800 0.000 480.080 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 487.160 0.000 487.440 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.520 0.000 494.800 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.880 0.000 502.160 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.240 0.000 509.520 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 516.600 0.000 516.880 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.960 0.000 524.240 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.320 0.000 531.600 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.680 0.000 538.960 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.040 0.000 546.320 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.540 0.000 281.820 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.400 0.000 553.680 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.760 0.000 561.040 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.120 0.000 568.400 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.480 0.000 575.760 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 582.840 0.000 583.120 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.200 0.000 590.480 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.560 0.000 597.840 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.920 0.000 605.200 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 612.280 0.000 612.560 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.640 0.000 619.920 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.900 0.000 289.180 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.000 0.000 627.280 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 634.360 0.000 634.640 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 641.720 0.000 642.000 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.620 0.000 648.900 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.980 0.000 656.260 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 663.340 0.000 663.620 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.700 0.000 670.980 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 678.060 0.000 678.340 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.420 0.000 685.700 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 692.780 0.000 693.060 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 296.260 0.000 296.540 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.140 0.000 700.420 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.500 0.000 707.780 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.860 0.000 715.140 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.220 0.000 722.500 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.580 0.000 729.860 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 736.940 0.000 737.220 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.300 0.000 744.580 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 751.660 0.000 751.940 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.020 0.000 759.300 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 766.380 0.000 766.660 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.620 0.000 303.900 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 773.740 0.000 774.020 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.100 0.000 781.380 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.460 0.000 788.740 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 795.820 0.000 796.100 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.180 0.000 803.460 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 810.540 0.000 810.820 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.900 0.000 818.180 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.260 0.000 825.540 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 832.620 0.000 832.900 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 839.980 0.000 840.260 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.980 0.000 311.260 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 847.340 0.000 847.620 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.700 0.000 854.980 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 862.060 0.000 862.340 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.420 0.000 869.700 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.780 0.000 877.060 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.140 0.000 884.420 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.500 0.000 891.780 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 898.860 0.000 899.140 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 906.220 0.000 906.500 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.580 0.000 913.860 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.340 0.000 318.620 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.940 0.000 921.220 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.840 0.000 928.120 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.200 0.000 935.480 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.560 0.000 942.840 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.920 0.000 950.200 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 957.280 0.000 957.560 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 964.640 0.000 964.920 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 972.000 0.000 972.280 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.360 0.000 979.640 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 986.720 0.000 987.000 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.700 0.000 325.980 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 261.760 0.000 262.040 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 996.840 0.000 997.120 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1004.200 0.000 1004.480 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1011.560 0.000 1011.840 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1018.460 0.000 1018.740 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1025.820 0.000 1026.100 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1033.180 0.000 1033.460 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1040.540 0.000 1040.820 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1047.900 0.000 1048.180 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1055.260 0.000 1055.540 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1062.620 0.000 1062.900 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.360 0.000 335.640 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1069.980 0.000 1070.260 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1077.340 0.000 1077.620 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.700 0.000 1084.980 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1092.060 0.000 1092.340 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1099.420 0.000 1099.700 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1106.780 0.000 1107.060 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1114.140 0.000 1114.420 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1121.500 0.000 1121.780 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1128.860 0.000 1129.140 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1136.220 0.000 1136.500 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 342.720 0.000 343.000 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1143.580 0.000 1143.860 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1150.940 0.000 1151.220 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1158.300 0.000 1158.580 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1165.660 0.000 1165.940 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.020 0.000 1173.300 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1180.380 0.000 1180.660 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1187.740 0.000 1188.020 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1195.100 0.000 1195.380 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 350.080 0.000 350.360 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.440 0.000 357.720 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.800 0.000 365.080 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.160 0.000 372.440 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.520 0.000 379.800 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 386.880 0.000 387.160 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.240 0.000 394.520 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.600 0.000 401.880 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.120 0.000 269.400 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.960 0.000 409.240 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 416.320 0.000 416.600 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.680 0.000 423.960 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.040 0.000 431.320 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.400 0.000 438.680 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.760 0.000 446.040 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.120 0.000 453.400 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 460.480 0.000 460.760 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.380 0.000 467.660 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 474.740 0.000 475.020 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.480 0.000 276.760 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.100 0.000 482.380 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.460 0.000 489.740 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.820 0.000 497.100 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 504.180 0.000 504.460 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.540 0.000 511.820 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 518.900 0.000 519.180 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.260 0.000 526.540 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.620 0.000 533.900 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.980 0.000 541.260 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 548.340 0.000 548.620 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.840 0.000 284.120 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.700 0.000 555.980 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.060 0.000 563.340 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.420 0.000 570.700 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 577.780 0.000 578.060 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.140 0.000 585.420 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.500 0.000 592.780 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 599.860 0.000 600.140 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 607.220 0.000 607.500 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.580 0.000 614.860 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.940 0.000 622.220 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.200 0.000 291.480 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 629.300 0.000 629.580 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 636.660 0.000 636.940 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.020 0.000 644.300 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 651.380 0.000 651.660 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 658.740 0.000 659.020 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 666.100 0.000 666.380 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.460 0.000 673.740 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 680.820 0.000 681.100 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 688.180 0.000 688.460 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 695.540 0.000 695.820 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.560 0.000 298.840 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 702.900 0.000 703.180 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.260 0.000 710.540 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 717.620 0.000 717.900 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.980 0.000 725.260 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 732.340 0.000 732.620 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 739.240 0.000 739.520 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.600 0.000 746.880 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.960 0.000 754.240 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 761.320 0.000 761.600 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.680 0.000 768.960 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.920 0.000 306.200 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 776.040 0.000 776.320 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.400 0.000 783.680 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 790.760 0.000 791.040 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 798.120 0.000 798.400 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.480 0.000 805.760 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 812.840 0.000 813.120 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 820.200 0.000 820.480 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 827.560 0.000 827.840 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 834.920 0.000 835.200 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 842.280 0.000 842.560 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.280 0.000 313.560 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 849.640 0.000 849.920 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 857.000 0.000 857.280 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 864.360 0.000 864.640 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 871.720 0.000 872.000 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.080 0.000 879.360 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.440 0.000 886.720 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.800 0.000 894.080 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 901.160 0.000 901.440 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 908.520 0.000 908.800 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.880 0.000 916.160 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.640 0.000 320.920 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 923.240 0.000 923.520 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 930.600 0.000 930.880 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.960 0.000 938.240 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 945.320 0.000 945.600 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 952.680 0.000 952.960 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.040 0.000 960.320 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.400 0.000 967.680 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.760 0.000 975.040 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 982.120 0.000 982.400 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.480 0.000 989.760 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.000 0.000 328.280 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.520 0.000 264.800 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 999.140 0.000 999.420 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.500 0.000 1006.780 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.860 0.000 1014.140 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.220 0.000 1021.500 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.580 0.000 1028.860 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.940 0.000 1036.220 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.300 0.000 1043.580 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.660 0.000 1050.940 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.020 0.000 1058.300 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.380 0.000 1065.660 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.660 0.000 337.940 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.740 0.000 1073.020 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.100 0.000 1080.380 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.460 0.000 1087.740 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.820 0.000 1095.100 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1102.180 0.000 1102.460 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.080 0.000 1109.360 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.440 0.000 1116.720 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1123.800 0.000 1124.080 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.160 0.000 1131.440 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1138.520 0.000 1138.800 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.020 0.000 345.300 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.880 0.000 1146.160 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1153.240 0.000 1153.520 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.600 0.000 1160.880 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1167.960 0.000 1168.240 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.320 0.000 1175.600 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1182.680 0.000 1182.960 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1190.040 0.000 1190.320 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.400 0.000 1197.680 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.380 0.000 352.660 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.740 0.000 360.020 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.100 0.000 367.380 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.460 0.000 374.740 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.820 0.000 382.100 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.180 0.000 389.460 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.540 0.000 396.820 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.900 0.000 404.180 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.880 0.000 272.160 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 411.260 0.000 411.540 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.620 0.000 418.900 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.980 0.000 426.260 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.340 0.000 433.620 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.700 0.000 440.980 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.060 0.000 448.340 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.420 0.000 455.700 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.780 0.000 463.060 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.140 0.000 470.420 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.500 0.000 477.780 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.780 0.000 279.060 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.860 0.000 485.140 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.220 0.000 492.500 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.580 0.000 499.860 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.940 0.000 507.220 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.300 0.000 514.580 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 521.660 0.000 521.940 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 529.020 0.000 529.300 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.380 0.000 536.660 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.740 0.000 544.020 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.100 0.000 551.380 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.140 0.000 286.420 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.000 0.000 558.280 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.360 0.000 565.640 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.720 0.000 573.000 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.080 0.000 580.360 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.440 0.000 587.720 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 594.800 0.000 595.080 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 602.160 0.000 602.440 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.520 0.000 609.800 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.880 0.000 617.160 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 624.240 0.000 624.520 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.500 0.000 293.780 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 631.600 0.000 631.880 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 638.960 0.000 639.240 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 646.320 0.000 646.600 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.680 0.000 653.960 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.040 0.000 661.320 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.400 0.000 668.680 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.760 0.000 676.040 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 683.120 0.000 683.400 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.480 0.000 690.760 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 697.840 0.000 698.120 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.860 0.000 301.140 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.200 0.000 705.480 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 712.560 0.000 712.840 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 719.920 0.000 720.200 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.280 0.000 727.560 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.640 0.000 734.920 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.000 0.000 742.280 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 749.360 0.000 749.640 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 756.720 0.000 757.000 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 764.080 0.000 764.360 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.440 0.000 771.720 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 308.220 0.000 308.500 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 778.800 0.000 779.080 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 786.160 0.000 786.440 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.520 0.000 793.800 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.880 0.000 801.160 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 808.240 0.000 808.520 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 815.600 0.000 815.880 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.960 0.000 823.240 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.320 0.000 830.600 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.220 0.000 837.500 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.580 0.000 844.860 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.580 0.000 315.860 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.940 0.000 852.220 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 859.300 0.000 859.580 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.660 0.000 866.940 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.020 0.000 874.300 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.380 0.000 881.660 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.740 0.000 889.020 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.100 0.000 896.380 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 903.460 0.000 903.740 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 910.820 0.000 911.100 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.180 0.000 918.460 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.940 0.000 323.220 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 925.540 0.000 925.820 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.900 0.000 933.180 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.260 0.000 940.540 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 947.620 0.000 947.900 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.980 0.000 955.260 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.340 0.000 962.620 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.700 0.000 969.980 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.060 0.000 977.340 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.420 0.000 984.700 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.780 0.000 992.060 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.300 0.000 330.580 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.320 0.000 2.600 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.620 0.000 4.900 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.280 0.000 14.560 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.540 0.000 97.820 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.900 0.000 105.180 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.260 0.000 112.540 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.620 0.000 119.900 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.980 0.000 127.260 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.340 0.000 134.620 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.700 0.000 141.980 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.060 0.000 149.340 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.420 0.000 156.700 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.780 0.000 164.060 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.400 0.000 24.680 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.140 0.000 171.420 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.500 0.000 178.780 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.860 0.000 186.140 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.220 0.000 193.500 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.580 0.000 200.860 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.940 0.000 208.220 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.300 0.000 215.580 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.660 0.000 222.940 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.020 0.000 230.300 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.380 0.000 237.660 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.060 0.000 34.340 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.740 0.000 245.020 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.100 0.000 252.380 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.840 0.000 54.120 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.200 0.000 61.480 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.560 0.000 68.840 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.920 0.000 76.200 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.280 0.000 83.560 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.640 0.000 90.920 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.920 0.000 7.200 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.040 0.000 17.320 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.300 0.000 100.580 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.660 0.000 107.940 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.020 0.000 115.300 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.380 0.000 122.660 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.740 0.000 130.020 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.100 0.000 137.380 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.460 0.000 144.740 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.820 0.000 152.100 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.180 0.000 159.460 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.540 0.000 166.820 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.700 0.000 26.980 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.900 0.000 174.180 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.260 0.000 181.540 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.160 0.000 188.440 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.520 0.000 195.800 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.880 0.000 203.160 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.240 0.000 210.520 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.600 0.000 217.880 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.960 0.000 225.240 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.320 0.000 232.600 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.680 0.000 239.960 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.360 0.000 36.640 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.040 0.000 247.320 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.400 0.000 254.680 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.480 0.000 46.760 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.140 0.000 56.420 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.500 0.000 63.780 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.860 0.000 71.140 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.220 0.000 78.500 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.580 0.000 85.860 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.940 0.000 93.220 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.340 0.000 19.620 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.600 0.000 102.880 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.960 0.000 110.240 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.320 0.000 117.600 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.680 0.000 124.960 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.040 0.000 132.320 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.400 0.000 139.680 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.760 0.000 147.040 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.120 0.000 154.400 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.480 0.000 161.760 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.840 0.000 169.120 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.000 0.000 29.280 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.200 0.000 176.480 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.560 0.000 183.840 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.920 0.000 191.200 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.280 0.000 198.560 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.640 0.000 205.920 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.000 0.000 213.280 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.360 0.000 220.640 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 227.720 0.000 228.000 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.080 0.000 235.360 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 242.440 0.000 242.720 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.120 0.000 39.400 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.800 0.000 250.080 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.160 0.000 257.440 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.780 0.000 49.060 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.440 0.000 58.720 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.800 0.000 66.080 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.160 0.000 73.440 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.520 0.000 80.800 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.880 0.000 88.160 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.240 0.000 95.520 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.640 0.000 21.920 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.760 0.000 32.040 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.420 0.000 41.700 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.080 0.000 51.360 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.680 0.000 9.960 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.980 0.000 12.260 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.050 10.640 21.650 1188.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.850 10.640 98.450 1188.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.530 10.795 1193.170 1188.725 ;
      LAYER met1 ;
        RECT 0.000 4.800 1197.700 1188.880 ;
      LAYER met2 ;
        RECT 0.030 1195.720 3.880 1196.000 ;
        RECT 4.720 1195.720 14.000 1196.000 ;
        RECT 14.840 1195.720 24.580 1196.000 ;
        RECT 25.420 1195.720 35.160 1196.000 ;
        RECT 36.000 1195.720 45.740 1196.000 ;
        RECT 46.580 1195.720 56.320 1196.000 ;
        RECT 57.160 1195.720 66.900 1196.000 ;
        RECT 67.740 1195.720 77.480 1196.000 ;
        RECT 78.320 1195.720 88.060 1196.000 ;
        RECT 88.900 1195.720 98.180 1196.000 ;
        RECT 99.020 1195.720 108.760 1196.000 ;
        RECT 109.600 1195.720 119.340 1196.000 ;
        RECT 120.180 1195.720 129.920 1196.000 ;
        RECT 130.760 1195.720 140.500 1196.000 ;
        RECT 141.340 1195.720 151.080 1196.000 ;
        RECT 151.920 1195.720 161.660 1196.000 ;
        RECT 162.500 1195.720 172.240 1196.000 ;
        RECT 173.080 1195.720 182.820 1196.000 ;
        RECT 183.660 1195.720 192.940 1196.000 ;
        RECT 193.780 1195.720 203.520 1196.000 ;
        RECT 204.360 1195.720 214.100 1196.000 ;
        RECT 214.940 1195.720 224.680 1196.000 ;
        RECT 225.520 1195.720 235.260 1196.000 ;
        RECT 236.100 1195.720 245.840 1196.000 ;
        RECT 246.680 1195.720 256.420 1196.000 ;
        RECT 257.260 1195.720 267.000 1196.000 ;
        RECT 267.840 1195.720 277.580 1196.000 ;
        RECT 278.420 1195.720 287.700 1196.000 ;
        RECT 288.540 1195.720 298.280 1196.000 ;
        RECT 299.120 1195.720 308.860 1196.000 ;
        RECT 309.700 1195.720 319.440 1196.000 ;
        RECT 320.280 1195.720 330.020 1196.000 ;
        RECT 330.860 1195.720 340.600 1196.000 ;
        RECT 341.440 1195.720 351.180 1196.000 ;
        RECT 352.020 1195.720 361.760 1196.000 ;
        RECT 362.600 1195.720 372.340 1196.000 ;
        RECT 373.180 1195.720 382.460 1196.000 ;
        RECT 383.300 1195.720 393.040 1196.000 ;
        RECT 393.880 1195.720 403.620 1196.000 ;
        RECT 404.460 1195.720 414.200 1196.000 ;
        RECT 415.040 1195.720 424.780 1196.000 ;
        RECT 425.620 1195.720 435.360 1196.000 ;
        RECT 436.200 1195.720 445.940 1196.000 ;
        RECT 446.780 1195.720 456.520 1196.000 ;
        RECT 457.360 1195.720 466.640 1196.000 ;
        RECT 467.480 1195.720 477.220 1196.000 ;
        RECT 478.060 1195.720 487.800 1196.000 ;
        RECT 488.640 1195.720 498.380 1196.000 ;
        RECT 499.220 1195.720 508.960 1196.000 ;
        RECT 509.800 1195.720 519.540 1196.000 ;
        RECT 520.380 1195.720 530.120 1196.000 ;
        RECT 530.960 1195.720 540.700 1196.000 ;
        RECT 541.540 1195.720 551.280 1196.000 ;
        RECT 552.120 1195.720 561.400 1196.000 ;
        RECT 562.240 1195.720 571.980 1196.000 ;
        RECT 572.820 1195.720 582.560 1196.000 ;
        RECT 583.400 1195.720 593.140 1196.000 ;
        RECT 593.980 1195.720 603.720 1196.000 ;
        RECT 604.560 1195.720 614.300 1196.000 ;
        RECT 615.140 1195.720 624.880 1196.000 ;
        RECT 625.720 1195.720 635.460 1196.000 ;
        RECT 636.300 1195.720 646.040 1196.000 ;
        RECT 646.880 1195.720 656.160 1196.000 ;
        RECT 657.000 1195.720 666.740 1196.000 ;
        RECT 667.580 1195.720 677.320 1196.000 ;
        RECT 678.160 1195.720 687.900 1196.000 ;
        RECT 688.740 1195.720 698.480 1196.000 ;
        RECT 699.320 1195.720 709.060 1196.000 ;
        RECT 709.900 1195.720 719.640 1196.000 ;
        RECT 720.480 1195.720 730.220 1196.000 ;
        RECT 731.060 1195.720 740.800 1196.000 ;
        RECT 741.640 1195.720 750.920 1196.000 ;
        RECT 751.760 1195.720 761.500 1196.000 ;
        RECT 762.340 1195.720 772.080 1196.000 ;
        RECT 772.920 1195.720 782.660 1196.000 ;
        RECT 783.500 1195.720 793.240 1196.000 ;
        RECT 794.080 1195.720 803.820 1196.000 ;
        RECT 804.660 1195.720 814.400 1196.000 ;
        RECT 815.240 1195.720 824.980 1196.000 ;
        RECT 825.820 1195.720 835.100 1196.000 ;
        RECT 835.940 1195.720 845.680 1196.000 ;
        RECT 846.520 1195.720 856.260 1196.000 ;
        RECT 857.100 1195.720 866.840 1196.000 ;
        RECT 867.680 1195.720 877.420 1196.000 ;
        RECT 878.260 1195.720 888.000 1196.000 ;
        RECT 888.840 1195.720 898.580 1196.000 ;
        RECT 899.420 1195.720 909.160 1196.000 ;
        RECT 910.000 1195.720 919.740 1196.000 ;
        RECT 920.580 1195.720 929.860 1196.000 ;
        RECT 930.700 1195.720 940.440 1196.000 ;
        RECT 941.280 1195.720 951.020 1196.000 ;
        RECT 951.860 1195.720 961.600 1196.000 ;
        RECT 962.440 1195.720 972.180 1196.000 ;
        RECT 973.020 1195.720 982.760 1196.000 ;
        RECT 983.600 1195.720 993.340 1196.000 ;
        RECT 994.180 1195.720 1003.920 1196.000 ;
        RECT 1004.760 1195.720 1014.500 1196.000 ;
        RECT 1015.340 1195.720 1024.620 1196.000 ;
        RECT 1025.460 1195.720 1035.200 1196.000 ;
        RECT 1036.040 1195.720 1045.780 1196.000 ;
        RECT 1046.620 1195.720 1056.360 1196.000 ;
        RECT 1057.200 1195.720 1066.940 1196.000 ;
        RECT 1067.780 1195.720 1077.520 1196.000 ;
        RECT 1078.360 1195.720 1088.100 1196.000 ;
        RECT 1088.940 1195.720 1098.680 1196.000 ;
        RECT 1099.520 1195.720 1109.260 1196.000 ;
        RECT 1110.100 1195.720 1119.380 1196.000 ;
        RECT 1120.220 1195.720 1129.960 1196.000 ;
        RECT 1130.800 1195.720 1140.540 1196.000 ;
        RECT 1141.380 1195.720 1151.120 1196.000 ;
        RECT 1151.960 1195.720 1161.700 1196.000 ;
        RECT 1162.540 1195.720 1172.280 1196.000 ;
        RECT 1173.120 1195.720 1182.860 1196.000 ;
        RECT 1183.700 1195.720 1193.440 1196.000 ;
        RECT 1194.280 1195.720 1197.670 1196.000 ;
        RECT 0.030 4.280 1197.670 1195.720 ;
        RECT 0.580 4.000 2.040 4.280 ;
        RECT 2.880 4.000 4.340 4.280 ;
        RECT 5.180 4.000 6.640 4.280 ;
        RECT 7.480 4.000 9.400 4.280 ;
        RECT 10.240 4.000 11.700 4.280 ;
        RECT 12.540 4.000 14.000 4.280 ;
        RECT 14.840 4.000 16.760 4.280 ;
        RECT 17.600 4.000 19.060 4.280 ;
        RECT 19.900 4.000 21.360 4.280 ;
        RECT 22.200 4.000 24.120 4.280 ;
        RECT 24.960 4.000 26.420 4.280 ;
        RECT 27.260 4.000 28.720 4.280 ;
        RECT 29.560 4.000 31.480 4.280 ;
        RECT 32.320 4.000 33.780 4.280 ;
        RECT 34.620 4.000 36.080 4.280 ;
        RECT 36.920 4.000 38.840 4.280 ;
        RECT 39.680 4.000 41.140 4.280 ;
        RECT 41.980 4.000 43.440 4.280 ;
        RECT 44.280 4.000 46.200 4.280 ;
        RECT 47.040 4.000 48.500 4.280 ;
        RECT 49.340 4.000 50.800 4.280 ;
        RECT 51.640 4.000 53.560 4.280 ;
        RECT 54.400 4.000 55.860 4.280 ;
        RECT 56.700 4.000 58.160 4.280 ;
        RECT 59.000 4.000 60.920 4.280 ;
        RECT 61.760 4.000 63.220 4.280 ;
        RECT 64.060 4.000 65.520 4.280 ;
        RECT 66.360 4.000 68.280 4.280 ;
        RECT 69.120 4.000 70.580 4.280 ;
        RECT 71.420 4.000 72.880 4.280 ;
        RECT 73.720 4.000 75.640 4.280 ;
        RECT 76.480 4.000 77.940 4.280 ;
        RECT 78.780 4.000 80.240 4.280 ;
        RECT 81.080 4.000 83.000 4.280 ;
        RECT 83.840 4.000 85.300 4.280 ;
        RECT 86.140 4.000 87.600 4.280 ;
        RECT 88.440 4.000 90.360 4.280 ;
        RECT 91.200 4.000 92.660 4.280 ;
        RECT 93.500 4.000 94.960 4.280 ;
        RECT 95.800 4.000 97.260 4.280 ;
        RECT 98.100 4.000 100.020 4.280 ;
        RECT 100.860 4.000 102.320 4.280 ;
        RECT 103.160 4.000 104.620 4.280 ;
        RECT 105.460 4.000 107.380 4.280 ;
        RECT 108.220 4.000 109.680 4.280 ;
        RECT 110.520 4.000 111.980 4.280 ;
        RECT 112.820 4.000 114.740 4.280 ;
        RECT 115.580 4.000 117.040 4.280 ;
        RECT 117.880 4.000 119.340 4.280 ;
        RECT 120.180 4.000 122.100 4.280 ;
        RECT 122.940 4.000 124.400 4.280 ;
        RECT 125.240 4.000 126.700 4.280 ;
        RECT 127.540 4.000 129.460 4.280 ;
        RECT 130.300 4.000 131.760 4.280 ;
        RECT 132.600 4.000 134.060 4.280 ;
        RECT 134.900 4.000 136.820 4.280 ;
        RECT 137.660 4.000 139.120 4.280 ;
        RECT 139.960 4.000 141.420 4.280 ;
        RECT 142.260 4.000 144.180 4.280 ;
        RECT 145.020 4.000 146.480 4.280 ;
        RECT 147.320 4.000 148.780 4.280 ;
        RECT 149.620 4.000 151.540 4.280 ;
        RECT 152.380 4.000 153.840 4.280 ;
        RECT 154.680 4.000 156.140 4.280 ;
        RECT 156.980 4.000 158.900 4.280 ;
        RECT 159.740 4.000 161.200 4.280 ;
        RECT 162.040 4.000 163.500 4.280 ;
        RECT 164.340 4.000 166.260 4.280 ;
        RECT 167.100 4.000 168.560 4.280 ;
        RECT 169.400 4.000 170.860 4.280 ;
        RECT 171.700 4.000 173.620 4.280 ;
        RECT 174.460 4.000 175.920 4.280 ;
        RECT 176.760 4.000 178.220 4.280 ;
        RECT 179.060 4.000 180.980 4.280 ;
        RECT 181.820 4.000 183.280 4.280 ;
        RECT 184.120 4.000 185.580 4.280 ;
        RECT 186.420 4.000 187.880 4.280 ;
        RECT 188.720 4.000 190.640 4.280 ;
        RECT 191.480 4.000 192.940 4.280 ;
        RECT 193.780 4.000 195.240 4.280 ;
        RECT 196.080 4.000 198.000 4.280 ;
        RECT 198.840 4.000 200.300 4.280 ;
        RECT 201.140 4.000 202.600 4.280 ;
        RECT 203.440 4.000 205.360 4.280 ;
        RECT 206.200 4.000 207.660 4.280 ;
        RECT 208.500 4.000 209.960 4.280 ;
        RECT 210.800 4.000 212.720 4.280 ;
        RECT 213.560 4.000 215.020 4.280 ;
        RECT 215.860 4.000 217.320 4.280 ;
        RECT 218.160 4.000 220.080 4.280 ;
        RECT 220.920 4.000 222.380 4.280 ;
        RECT 223.220 4.000 224.680 4.280 ;
        RECT 225.520 4.000 227.440 4.280 ;
        RECT 228.280 4.000 229.740 4.280 ;
        RECT 230.580 4.000 232.040 4.280 ;
        RECT 232.880 4.000 234.800 4.280 ;
        RECT 235.640 4.000 237.100 4.280 ;
        RECT 237.940 4.000 239.400 4.280 ;
        RECT 240.240 4.000 242.160 4.280 ;
        RECT 243.000 4.000 244.460 4.280 ;
        RECT 245.300 4.000 246.760 4.280 ;
        RECT 247.600 4.000 249.520 4.280 ;
        RECT 250.360 4.000 251.820 4.280 ;
        RECT 252.660 4.000 254.120 4.280 ;
        RECT 254.960 4.000 256.880 4.280 ;
        RECT 257.720 4.000 259.180 4.280 ;
        RECT 260.020 4.000 261.480 4.280 ;
        RECT 262.320 4.000 264.240 4.280 ;
        RECT 265.080 4.000 266.540 4.280 ;
        RECT 267.380 4.000 268.840 4.280 ;
        RECT 269.680 4.000 271.600 4.280 ;
        RECT 272.440 4.000 273.900 4.280 ;
        RECT 274.740 4.000 276.200 4.280 ;
        RECT 277.040 4.000 278.500 4.280 ;
        RECT 279.340 4.000 281.260 4.280 ;
        RECT 282.100 4.000 283.560 4.280 ;
        RECT 284.400 4.000 285.860 4.280 ;
        RECT 286.700 4.000 288.620 4.280 ;
        RECT 289.460 4.000 290.920 4.280 ;
        RECT 291.760 4.000 293.220 4.280 ;
        RECT 294.060 4.000 295.980 4.280 ;
        RECT 296.820 4.000 298.280 4.280 ;
        RECT 299.120 4.000 300.580 4.280 ;
        RECT 301.420 4.000 303.340 4.280 ;
        RECT 304.180 4.000 305.640 4.280 ;
        RECT 306.480 4.000 307.940 4.280 ;
        RECT 308.780 4.000 310.700 4.280 ;
        RECT 311.540 4.000 313.000 4.280 ;
        RECT 313.840 4.000 315.300 4.280 ;
        RECT 316.140 4.000 318.060 4.280 ;
        RECT 318.900 4.000 320.360 4.280 ;
        RECT 321.200 4.000 322.660 4.280 ;
        RECT 323.500 4.000 325.420 4.280 ;
        RECT 326.260 4.000 327.720 4.280 ;
        RECT 328.560 4.000 330.020 4.280 ;
        RECT 330.860 4.000 332.780 4.280 ;
        RECT 333.620 4.000 335.080 4.280 ;
        RECT 335.920 4.000 337.380 4.280 ;
        RECT 338.220 4.000 340.140 4.280 ;
        RECT 340.980 4.000 342.440 4.280 ;
        RECT 343.280 4.000 344.740 4.280 ;
        RECT 345.580 4.000 347.500 4.280 ;
        RECT 348.340 4.000 349.800 4.280 ;
        RECT 350.640 4.000 352.100 4.280 ;
        RECT 352.940 4.000 354.860 4.280 ;
        RECT 355.700 4.000 357.160 4.280 ;
        RECT 358.000 4.000 359.460 4.280 ;
        RECT 360.300 4.000 362.220 4.280 ;
        RECT 363.060 4.000 364.520 4.280 ;
        RECT 365.360 4.000 366.820 4.280 ;
        RECT 367.660 4.000 369.120 4.280 ;
        RECT 369.960 4.000 371.880 4.280 ;
        RECT 372.720 4.000 374.180 4.280 ;
        RECT 375.020 4.000 376.480 4.280 ;
        RECT 377.320 4.000 379.240 4.280 ;
        RECT 380.080 4.000 381.540 4.280 ;
        RECT 382.380 4.000 383.840 4.280 ;
        RECT 384.680 4.000 386.600 4.280 ;
        RECT 387.440 4.000 388.900 4.280 ;
        RECT 389.740 4.000 391.200 4.280 ;
        RECT 392.040 4.000 393.960 4.280 ;
        RECT 394.800 4.000 396.260 4.280 ;
        RECT 397.100 4.000 398.560 4.280 ;
        RECT 399.400 4.000 401.320 4.280 ;
        RECT 402.160 4.000 403.620 4.280 ;
        RECT 404.460 4.000 405.920 4.280 ;
        RECT 406.760 4.000 408.680 4.280 ;
        RECT 409.520 4.000 410.980 4.280 ;
        RECT 411.820 4.000 413.280 4.280 ;
        RECT 414.120 4.000 416.040 4.280 ;
        RECT 416.880 4.000 418.340 4.280 ;
        RECT 419.180 4.000 420.640 4.280 ;
        RECT 421.480 4.000 423.400 4.280 ;
        RECT 424.240 4.000 425.700 4.280 ;
        RECT 426.540 4.000 428.000 4.280 ;
        RECT 428.840 4.000 430.760 4.280 ;
        RECT 431.600 4.000 433.060 4.280 ;
        RECT 433.900 4.000 435.360 4.280 ;
        RECT 436.200 4.000 438.120 4.280 ;
        RECT 438.960 4.000 440.420 4.280 ;
        RECT 441.260 4.000 442.720 4.280 ;
        RECT 443.560 4.000 445.480 4.280 ;
        RECT 446.320 4.000 447.780 4.280 ;
        RECT 448.620 4.000 450.080 4.280 ;
        RECT 450.920 4.000 452.840 4.280 ;
        RECT 453.680 4.000 455.140 4.280 ;
        RECT 455.980 4.000 457.440 4.280 ;
        RECT 458.280 4.000 460.200 4.280 ;
        RECT 461.040 4.000 462.500 4.280 ;
        RECT 463.340 4.000 464.800 4.280 ;
        RECT 465.640 4.000 467.100 4.280 ;
        RECT 467.940 4.000 469.860 4.280 ;
        RECT 470.700 4.000 472.160 4.280 ;
        RECT 473.000 4.000 474.460 4.280 ;
        RECT 475.300 4.000 477.220 4.280 ;
        RECT 478.060 4.000 479.520 4.280 ;
        RECT 480.360 4.000 481.820 4.280 ;
        RECT 482.660 4.000 484.580 4.280 ;
        RECT 485.420 4.000 486.880 4.280 ;
        RECT 487.720 4.000 489.180 4.280 ;
        RECT 490.020 4.000 491.940 4.280 ;
        RECT 492.780 4.000 494.240 4.280 ;
        RECT 495.080 4.000 496.540 4.280 ;
        RECT 497.380 4.000 499.300 4.280 ;
        RECT 500.140 4.000 501.600 4.280 ;
        RECT 502.440 4.000 503.900 4.280 ;
        RECT 504.740 4.000 506.660 4.280 ;
        RECT 507.500 4.000 508.960 4.280 ;
        RECT 509.800 4.000 511.260 4.280 ;
        RECT 512.100 4.000 514.020 4.280 ;
        RECT 514.860 4.000 516.320 4.280 ;
        RECT 517.160 4.000 518.620 4.280 ;
        RECT 519.460 4.000 521.380 4.280 ;
        RECT 522.220 4.000 523.680 4.280 ;
        RECT 524.520 4.000 525.980 4.280 ;
        RECT 526.820 4.000 528.740 4.280 ;
        RECT 529.580 4.000 531.040 4.280 ;
        RECT 531.880 4.000 533.340 4.280 ;
        RECT 534.180 4.000 536.100 4.280 ;
        RECT 536.940 4.000 538.400 4.280 ;
        RECT 539.240 4.000 540.700 4.280 ;
        RECT 541.540 4.000 543.460 4.280 ;
        RECT 544.300 4.000 545.760 4.280 ;
        RECT 546.600 4.000 548.060 4.280 ;
        RECT 548.900 4.000 550.820 4.280 ;
        RECT 551.660 4.000 553.120 4.280 ;
        RECT 553.960 4.000 555.420 4.280 ;
        RECT 556.260 4.000 557.720 4.280 ;
        RECT 558.560 4.000 560.480 4.280 ;
        RECT 561.320 4.000 562.780 4.280 ;
        RECT 563.620 4.000 565.080 4.280 ;
        RECT 565.920 4.000 567.840 4.280 ;
        RECT 568.680 4.000 570.140 4.280 ;
        RECT 570.980 4.000 572.440 4.280 ;
        RECT 573.280 4.000 575.200 4.280 ;
        RECT 576.040 4.000 577.500 4.280 ;
        RECT 578.340 4.000 579.800 4.280 ;
        RECT 580.640 4.000 582.560 4.280 ;
        RECT 583.400 4.000 584.860 4.280 ;
        RECT 585.700 4.000 587.160 4.280 ;
        RECT 588.000 4.000 589.920 4.280 ;
        RECT 590.760 4.000 592.220 4.280 ;
        RECT 593.060 4.000 594.520 4.280 ;
        RECT 595.360 4.000 597.280 4.280 ;
        RECT 598.120 4.000 599.580 4.280 ;
        RECT 600.420 4.000 601.880 4.280 ;
        RECT 602.720 4.000 604.640 4.280 ;
        RECT 605.480 4.000 606.940 4.280 ;
        RECT 607.780 4.000 609.240 4.280 ;
        RECT 610.080 4.000 612.000 4.280 ;
        RECT 612.840 4.000 614.300 4.280 ;
        RECT 615.140 4.000 616.600 4.280 ;
        RECT 617.440 4.000 619.360 4.280 ;
        RECT 620.200 4.000 621.660 4.280 ;
        RECT 622.500 4.000 623.960 4.280 ;
        RECT 624.800 4.000 626.720 4.280 ;
        RECT 627.560 4.000 629.020 4.280 ;
        RECT 629.860 4.000 631.320 4.280 ;
        RECT 632.160 4.000 634.080 4.280 ;
        RECT 634.920 4.000 636.380 4.280 ;
        RECT 637.220 4.000 638.680 4.280 ;
        RECT 639.520 4.000 641.440 4.280 ;
        RECT 642.280 4.000 643.740 4.280 ;
        RECT 644.580 4.000 646.040 4.280 ;
        RECT 646.880 4.000 648.340 4.280 ;
        RECT 649.180 4.000 651.100 4.280 ;
        RECT 651.940 4.000 653.400 4.280 ;
        RECT 654.240 4.000 655.700 4.280 ;
        RECT 656.540 4.000 658.460 4.280 ;
        RECT 659.300 4.000 660.760 4.280 ;
        RECT 661.600 4.000 663.060 4.280 ;
        RECT 663.900 4.000 665.820 4.280 ;
        RECT 666.660 4.000 668.120 4.280 ;
        RECT 668.960 4.000 670.420 4.280 ;
        RECT 671.260 4.000 673.180 4.280 ;
        RECT 674.020 4.000 675.480 4.280 ;
        RECT 676.320 4.000 677.780 4.280 ;
        RECT 678.620 4.000 680.540 4.280 ;
        RECT 681.380 4.000 682.840 4.280 ;
        RECT 683.680 4.000 685.140 4.280 ;
        RECT 685.980 4.000 687.900 4.280 ;
        RECT 688.740 4.000 690.200 4.280 ;
        RECT 691.040 4.000 692.500 4.280 ;
        RECT 693.340 4.000 695.260 4.280 ;
        RECT 696.100 4.000 697.560 4.280 ;
        RECT 698.400 4.000 699.860 4.280 ;
        RECT 700.700 4.000 702.620 4.280 ;
        RECT 703.460 4.000 704.920 4.280 ;
        RECT 705.760 4.000 707.220 4.280 ;
        RECT 708.060 4.000 709.980 4.280 ;
        RECT 710.820 4.000 712.280 4.280 ;
        RECT 713.120 4.000 714.580 4.280 ;
        RECT 715.420 4.000 717.340 4.280 ;
        RECT 718.180 4.000 719.640 4.280 ;
        RECT 720.480 4.000 721.940 4.280 ;
        RECT 722.780 4.000 724.700 4.280 ;
        RECT 725.540 4.000 727.000 4.280 ;
        RECT 727.840 4.000 729.300 4.280 ;
        RECT 730.140 4.000 732.060 4.280 ;
        RECT 732.900 4.000 734.360 4.280 ;
        RECT 735.200 4.000 736.660 4.280 ;
        RECT 737.500 4.000 738.960 4.280 ;
        RECT 739.800 4.000 741.720 4.280 ;
        RECT 742.560 4.000 744.020 4.280 ;
        RECT 744.860 4.000 746.320 4.280 ;
        RECT 747.160 4.000 749.080 4.280 ;
        RECT 749.920 4.000 751.380 4.280 ;
        RECT 752.220 4.000 753.680 4.280 ;
        RECT 754.520 4.000 756.440 4.280 ;
        RECT 757.280 4.000 758.740 4.280 ;
        RECT 759.580 4.000 761.040 4.280 ;
        RECT 761.880 4.000 763.800 4.280 ;
        RECT 764.640 4.000 766.100 4.280 ;
        RECT 766.940 4.000 768.400 4.280 ;
        RECT 769.240 4.000 771.160 4.280 ;
        RECT 772.000 4.000 773.460 4.280 ;
        RECT 774.300 4.000 775.760 4.280 ;
        RECT 776.600 4.000 778.520 4.280 ;
        RECT 779.360 4.000 780.820 4.280 ;
        RECT 781.660 4.000 783.120 4.280 ;
        RECT 783.960 4.000 785.880 4.280 ;
        RECT 786.720 4.000 788.180 4.280 ;
        RECT 789.020 4.000 790.480 4.280 ;
        RECT 791.320 4.000 793.240 4.280 ;
        RECT 794.080 4.000 795.540 4.280 ;
        RECT 796.380 4.000 797.840 4.280 ;
        RECT 798.680 4.000 800.600 4.280 ;
        RECT 801.440 4.000 802.900 4.280 ;
        RECT 803.740 4.000 805.200 4.280 ;
        RECT 806.040 4.000 807.960 4.280 ;
        RECT 808.800 4.000 810.260 4.280 ;
        RECT 811.100 4.000 812.560 4.280 ;
        RECT 813.400 4.000 815.320 4.280 ;
        RECT 816.160 4.000 817.620 4.280 ;
        RECT 818.460 4.000 819.920 4.280 ;
        RECT 820.760 4.000 822.680 4.280 ;
        RECT 823.520 4.000 824.980 4.280 ;
        RECT 825.820 4.000 827.280 4.280 ;
        RECT 828.120 4.000 830.040 4.280 ;
        RECT 830.880 4.000 832.340 4.280 ;
        RECT 833.180 4.000 834.640 4.280 ;
        RECT 835.480 4.000 836.940 4.280 ;
        RECT 837.780 4.000 839.700 4.280 ;
        RECT 840.540 4.000 842.000 4.280 ;
        RECT 842.840 4.000 844.300 4.280 ;
        RECT 845.140 4.000 847.060 4.280 ;
        RECT 847.900 4.000 849.360 4.280 ;
        RECT 850.200 4.000 851.660 4.280 ;
        RECT 852.500 4.000 854.420 4.280 ;
        RECT 855.260 4.000 856.720 4.280 ;
        RECT 857.560 4.000 859.020 4.280 ;
        RECT 859.860 4.000 861.780 4.280 ;
        RECT 862.620 4.000 864.080 4.280 ;
        RECT 864.920 4.000 866.380 4.280 ;
        RECT 867.220 4.000 869.140 4.280 ;
        RECT 869.980 4.000 871.440 4.280 ;
        RECT 872.280 4.000 873.740 4.280 ;
        RECT 874.580 4.000 876.500 4.280 ;
        RECT 877.340 4.000 878.800 4.280 ;
        RECT 879.640 4.000 881.100 4.280 ;
        RECT 881.940 4.000 883.860 4.280 ;
        RECT 884.700 4.000 886.160 4.280 ;
        RECT 887.000 4.000 888.460 4.280 ;
        RECT 889.300 4.000 891.220 4.280 ;
        RECT 892.060 4.000 893.520 4.280 ;
        RECT 894.360 4.000 895.820 4.280 ;
        RECT 896.660 4.000 898.580 4.280 ;
        RECT 899.420 4.000 900.880 4.280 ;
        RECT 901.720 4.000 903.180 4.280 ;
        RECT 904.020 4.000 905.940 4.280 ;
        RECT 906.780 4.000 908.240 4.280 ;
        RECT 909.080 4.000 910.540 4.280 ;
        RECT 911.380 4.000 913.300 4.280 ;
        RECT 914.140 4.000 915.600 4.280 ;
        RECT 916.440 4.000 917.900 4.280 ;
        RECT 918.740 4.000 920.660 4.280 ;
        RECT 921.500 4.000 922.960 4.280 ;
        RECT 923.800 4.000 925.260 4.280 ;
        RECT 926.100 4.000 927.560 4.280 ;
        RECT 928.400 4.000 930.320 4.280 ;
        RECT 931.160 4.000 932.620 4.280 ;
        RECT 933.460 4.000 934.920 4.280 ;
        RECT 935.760 4.000 937.680 4.280 ;
        RECT 938.520 4.000 939.980 4.280 ;
        RECT 940.820 4.000 942.280 4.280 ;
        RECT 943.120 4.000 945.040 4.280 ;
        RECT 945.880 4.000 947.340 4.280 ;
        RECT 948.180 4.000 949.640 4.280 ;
        RECT 950.480 4.000 952.400 4.280 ;
        RECT 953.240 4.000 954.700 4.280 ;
        RECT 955.540 4.000 957.000 4.280 ;
        RECT 957.840 4.000 959.760 4.280 ;
        RECT 960.600 4.000 962.060 4.280 ;
        RECT 962.900 4.000 964.360 4.280 ;
        RECT 965.200 4.000 967.120 4.280 ;
        RECT 967.960 4.000 969.420 4.280 ;
        RECT 970.260 4.000 971.720 4.280 ;
        RECT 972.560 4.000 974.480 4.280 ;
        RECT 975.320 4.000 976.780 4.280 ;
        RECT 977.620 4.000 979.080 4.280 ;
        RECT 979.920 4.000 981.840 4.280 ;
        RECT 982.680 4.000 984.140 4.280 ;
        RECT 984.980 4.000 986.440 4.280 ;
        RECT 987.280 4.000 989.200 4.280 ;
        RECT 990.040 4.000 991.500 4.280 ;
        RECT 992.340 4.000 993.800 4.280 ;
        RECT 994.640 4.000 996.560 4.280 ;
        RECT 997.400 4.000 998.860 4.280 ;
        RECT 999.700 4.000 1001.160 4.280 ;
        RECT 1002.000 4.000 1003.920 4.280 ;
        RECT 1004.760 4.000 1006.220 4.280 ;
        RECT 1007.060 4.000 1008.520 4.280 ;
        RECT 1009.360 4.000 1011.280 4.280 ;
        RECT 1012.120 4.000 1013.580 4.280 ;
        RECT 1014.420 4.000 1015.880 4.280 ;
        RECT 1016.720 4.000 1018.180 4.280 ;
        RECT 1019.020 4.000 1020.940 4.280 ;
        RECT 1021.780 4.000 1023.240 4.280 ;
        RECT 1024.080 4.000 1025.540 4.280 ;
        RECT 1026.380 4.000 1028.300 4.280 ;
        RECT 1029.140 4.000 1030.600 4.280 ;
        RECT 1031.440 4.000 1032.900 4.280 ;
        RECT 1033.740 4.000 1035.660 4.280 ;
        RECT 1036.500 4.000 1037.960 4.280 ;
        RECT 1038.800 4.000 1040.260 4.280 ;
        RECT 1041.100 4.000 1043.020 4.280 ;
        RECT 1043.860 4.000 1045.320 4.280 ;
        RECT 1046.160 4.000 1047.620 4.280 ;
        RECT 1048.460 4.000 1050.380 4.280 ;
        RECT 1051.220 4.000 1052.680 4.280 ;
        RECT 1053.520 4.000 1054.980 4.280 ;
        RECT 1055.820 4.000 1057.740 4.280 ;
        RECT 1058.580 4.000 1060.040 4.280 ;
        RECT 1060.880 4.000 1062.340 4.280 ;
        RECT 1063.180 4.000 1065.100 4.280 ;
        RECT 1065.940 4.000 1067.400 4.280 ;
        RECT 1068.240 4.000 1069.700 4.280 ;
        RECT 1070.540 4.000 1072.460 4.280 ;
        RECT 1073.300 4.000 1074.760 4.280 ;
        RECT 1075.600 4.000 1077.060 4.280 ;
        RECT 1077.900 4.000 1079.820 4.280 ;
        RECT 1080.660 4.000 1082.120 4.280 ;
        RECT 1082.960 4.000 1084.420 4.280 ;
        RECT 1085.260 4.000 1087.180 4.280 ;
        RECT 1088.020 4.000 1089.480 4.280 ;
        RECT 1090.320 4.000 1091.780 4.280 ;
        RECT 1092.620 4.000 1094.540 4.280 ;
        RECT 1095.380 4.000 1096.840 4.280 ;
        RECT 1097.680 4.000 1099.140 4.280 ;
        RECT 1099.980 4.000 1101.900 4.280 ;
        RECT 1102.740 4.000 1104.200 4.280 ;
        RECT 1105.040 4.000 1106.500 4.280 ;
        RECT 1107.340 4.000 1108.800 4.280 ;
        RECT 1109.640 4.000 1111.560 4.280 ;
        RECT 1112.400 4.000 1113.860 4.280 ;
        RECT 1114.700 4.000 1116.160 4.280 ;
        RECT 1117.000 4.000 1118.920 4.280 ;
        RECT 1119.760 4.000 1121.220 4.280 ;
        RECT 1122.060 4.000 1123.520 4.280 ;
        RECT 1124.360 4.000 1126.280 4.280 ;
        RECT 1127.120 4.000 1128.580 4.280 ;
        RECT 1129.420 4.000 1130.880 4.280 ;
        RECT 1131.720 4.000 1133.640 4.280 ;
        RECT 1134.480 4.000 1135.940 4.280 ;
        RECT 1136.780 4.000 1138.240 4.280 ;
        RECT 1139.080 4.000 1141.000 4.280 ;
        RECT 1141.840 4.000 1143.300 4.280 ;
        RECT 1144.140 4.000 1145.600 4.280 ;
        RECT 1146.440 4.000 1148.360 4.280 ;
        RECT 1149.200 4.000 1150.660 4.280 ;
        RECT 1151.500 4.000 1152.960 4.280 ;
        RECT 1153.800 4.000 1155.720 4.280 ;
        RECT 1156.560 4.000 1158.020 4.280 ;
        RECT 1158.860 4.000 1160.320 4.280 ;
        RECT 1161.160 4.000 1163.080 4.280 ;
        RECT 1163.920 4.000 1165.380 4.280 ;
        RECT 1166.220 4.000 1167.680 4.280 ;
        RECT 1168.520 4.000 1170.440 4.280 ;
        RECT 1171.280 4.000 1172.740 4.280 ;
        RECT 1173.580 4.000 1175.040 4.280 ;
        RECT 1175.880 4.000 1177.800 4.280 ;
        RECT 1178.640 4.000 1180.100 4.280 ;
        RECT 1180.940 4.000 1182.400 4.280 ;
        RECT 1183.240 4.000 1185.160 4.280 ;
        RECT 1186.000 4.000 1187.460 4.280 ;
        RECT 1188.300 4.000 1189.760 4.280 ;
        RECT 1190.600 4.000 1192.520 4.280 ;
        RECT 1193.360 4.000 1194.820 4.280 ;
        RECT 1195.660 4.000 1197.120 4.280 ;
      LAYER met3 ;
        RECT 2.295 4.255 1183.905 1188.805 ;
      LAYER met4 ;
        RECT 67.385 10.640 96.450 1188.880 ;
        RECT 98.850 10.640 1173.650 1188.880 ;
  END
END user_proj_example
END LIBRARY

