magic
tech sky130A
magscale 1 2
timestamp 1607998175
<< locali >>
rect 364533 676243 364567 685797
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 364533 608651 364567 618205
rect 429393 601715 429427 608549
rect 559113 601715 559147 608549
rect 364625 589339 364659 598893
rect 429577 589339 429611 598893
rect 559297 589339 559331 598893
rect 247969 578595 248003 579309
rect 254225 578663 254259 579309
rect 292129 579139 292163 579309
rect 415685 578527 415719 579309
rect 428381 578459 428415 579309
rect 441077 578391 441111 579309
rect 453589 578323 453623 579309
rect 455797 578255 455831 579309
rect 87003 338045 87245 338079
rect 87095 337909 87245 337943
rect 87095 337773 87245 337807
rect 229109 337739 229143 338113
rect 230489 337705 230707 337739
rect 87095 337637 87429 337671
rect 115707 337569 115857 337603
rect 135027 337569 135177 337603
rect 154347 337569 154497 337603
rect 173667 337569 173817 337603
rect 192987 337569 193137 337603
rect 212307 337569 212457 337603
rect 220955 337569 221105 337603
rect 230489 337535 230523 337705
rect 230673 337671 230707 337705
rect 238677 337671 238711 338113
rect 230673 337637 231225 337671
rect 238769 337671 238803 338657
rect 318935 338045 319085 338079
rect 302191 337773 302283 337807
rect 302249 337739 302283 337773
rect 230581 337535 230615 337637
rect 234445 337467 234479 337637
rect 87095 337433 87153 337467
rect 220955 337433 221105 337467
rect 259745 337399 259779 337637
rect 220955 337297 221105 337331
rect 86969 336991 87003 337093
rect 103437 336991 103471 337229
rect 113189 336787 113223 337229
rect 220863 337229 221013 337263
rect 122757 336787 122791 337229
rect 303997 337195 304031 337773
rect 315497 337331 315531 338045
rect 318935 337909 318993 337943
rect 318843 337773 318993 337807
rect 327089 337739 327123 338113
rect 318935 337569 318993 337603
rect 318843 337433 319085 337467
rect 326353 337195 326387 337297
rect 334725 336787 334759 337365
rect 335829 337059 335863 337501
rect 335921 337399 335955 337841
rect 336013 337671 336047 337841
rect 336657 337739 336691 338113
rect 346409 337739 346443 338657
rect 344201 337637 344661 337671
rect 344201 337535 344235 337637
rect 336197 336923 336231 337365
rect 340797 337127 340831 337365
rect 340613 336787 340647 337025
rect 340889 336855 340923 337365
rect 341717 337263 341751 337501
rect 342821 337195 342855 337501
rect 345581 336923 345615 337365
rect 345857 336991 345891 337161
rect 354045 336991 354079 337365
rect 364993 337195 365027 337637
rect 365177 337603 365211 338113
rect 374653 337603 374687 338045
rect 376769 337671 376803 338045
rect 466377 338011 466411 338113
rect 412557 337603 412591 337841
rect 365119 337501 365269 337535
rect 414121 337467 414155 337705
rect 369869 337195 369903 337365
rect 374653 337195 374687 337433
rect 422953 337263 422987 337433
rect 427921 336923 427955 337161
rect 432245 336991 432279 337705
rect 437431 337569 437581 337603
rect 436753 337127 436787 337365
rect 441629 336855 441663 337909
rect 446413 337535 446447 337773
rect 448529 337535 448563 337773
rect 449173 337399 449207 337705
rect 345523 336821 345765 336855
rect 451105 336855 451139 337909
rect 451289 336787 451323 337909
rect 451473 337875 451507 337977
rect 451381 337399 451415 337705
rect 456073 337399 456107 337501
rect 456993 337331 457027 337569
rect 340613 336753 340797 336787
rect 341015 336753 341165 336787
rect 457177 336787 457211 337229
rect 459109 336855 459143 337569
rect 461409 337535 461443 337841
rect 461593 337807 461627 337977
rect 460397 337263 460431 337501
rect 461593 336855 461627 337297
rect 466285 336719 466319 337977
rect 466469 336923 466503 337297
rect 469229 337263 469263 337909
rect 470793 336923 470827 337365
rect 480913 336923 480947 337365
rect 489929 337127 489963 337365
rect 500233 337127 500267 337365
rect 250177 327131 250211 334441
rect 236469 318835 236503 321657
rect 259837 318835 259871 328389
rect 265265 325703 265299 335257
rect 284401 335223 284435 336685
rect 270785 328491 270819 334305
rect 272257 328491 272291 334305
rect 273545 321555 273579 327029
rect 285965 317543 285999 327029
rect 288817 318631 288851 336685
rect 302617 318835 302651 328389
rect 327273 327131 327307 336685
rect 337393 328423 337427 336685
rect 330125 318835 330159 327029
rect 337393 318835 337427 321589
rect 339785 318835 339819 336685
rect 341349 318835 341383 328389
rect 389465 318835 389499 328389
rect 470609 318835 470643 328389
rect 232329 298163 232363 307717
rect 239137 299523 239171 309077
rect 250177 307819 250211 317373
rect 251557 307819 251591 317373
rect 284585 306391 284619 311865
rect 285965 306459 285999 311865
rect 232237 288439 232271 297993
rect 236285 288439 236319 298061
rect 245945 298027 245979 302413
rect 250177 289799 250211 298061
rect 251373 288439 251407 298061
rect 272165 283611 272199 289765
rect 273637 287079 273671 296633
rect 288725 290003 288759 308397
rect 290105 306323 290139 313225
rect 299765 299523 299799 317373
rect 306757 316047 306791 317441
rect 310897 307887 310931 311933
rect 325893 307819 325927 317373
rect 372721 309179 372755 318733
rect 306849 296735 306883 299489
rect 310713 298163 310747 307717
rect 310897 282795 310931 293029
rect 323317 288439 323351 299421
rect 324697 289867 324731 299421
rect 337025 298231 337059 307717
rect 339877 299931 339911 309077
rect 341165 299523 341199 309077
rect 367017 299523 367051 309077
rect 389281 299523 389315 309009
rect 421205 307819 421239 317373
rect 470609 299523 470643 309077
rect 325985 288439 326019 298061
rect 327181 288439 327215 298061
rect 337209 292451 337243 298061
rect 372721 289867 372755 299421
rect 330309 287079 330343 288405
rect 270693 275315 270727 280109
rect 273545 270555 273579 280109
rect 337117 278783 337151 282897
rect 341165 280211 341199 289765
rect 367017 280211 367051 289765
rect 389373 280211 389407 289765
rect 421205 288439 421239 298061
rect 470609 280211 470643 289765
rect 232237 269127 232271 270521
rect 310897 263483 310931 278681
rect 324513 269127 324547 278681
rect 330125 263211 330159 277253
rect 270693 256003 270727 260797
rect 250085 249815 250119 253929
rect 273545 251243 273579 260797
rect 259653 242675 259687 251141
rect 270693 241587 270727 244273
rect 251373 240159 251407 241485
rect 244381 230503 244415 234821
rect 250177 230503 250211 234617
rect 270693 232067 270727 241417
rect 284677 240159 284711 249713
rect 290013 248455 290047 258009
rect 294245 248455 294279 258009
rect 306849 249815 306883 262905
rect 337117 259471 337151 263585
rect 341165 260899 341199 270453
rect 362233 263483 362267 277321
rect 372721 270555 372755 280109
rect 375849 270555 375883 280109
rect 377137 270555 377171 280109
rect 424609 270555 424643 280109
rect 367017 260899 367051 270453
rect 389373 260899 389407 270453
rect 470609 260899 470643 270453
rect 310897 251311 310931 256037
rect 285965 234515 285999 244953
rect 291485 240091 291519 248353
rect 310713 241519 310747 251141
rect 323409 241519 323443 252705
rect 372721 251243 372755 260797
rect 375849 251243 375883 260797
rect 377137 251243 377171 260797
rect 424517 251243 424551 260797
rect 463709 251243 463743 260797
rect 325893 249815 325927 251141
rect 266737 230503 266771 231897
rect 299489 231863 299523 241417
rect 327181 240227 327215 249713
rect 367017 241519 367051 251141
rect 470609 241519 470643 251141
rect 302617 230503 302651 231965
rect 323409 231795 323443 234685
rect 270693 222275 270727 224961
rect 310805 222207 310839 231761
rect 327181 230571 327215 240057
rect 362233 230503 362267 241417
rect 375849 231863 375883 241417
rect 389281 234651 389315 241417
rect 367017 222207 367051 231761
rect 232237 209831 232271 211225
rect 244473 200175 244507 217957
rect 270693 212755 270727 222105
rect 299489 212551 299523 222105
rect 272165 211191 272199 212517
rect 265265 202759 265299 211089
rect 310805 202895 310839 212449
rect 330125 209831 330159 219385
rect 341165 215271 341199 220745
rect 362141 211191 362175 215305
rect 375849 212551 375883 222105
rect 330217 202827 330251 209729
rect 244381 180863 244415 186949
rect 267749 183583 267783 186337
rect 270693 183583 270727 186337
rect 284677 183515 284711 198645
rect 291485 190519 291519 200073
rect 299489 193239 299523 202793
rect 336933 193239 336967 202793
rect 358645 191879 358679 201433
rect 362233 193239 362267 198033
rect 375849 193239 375883 202793
rect 299857 183583 299891 188445
rect 306849 183583 306883 188445
rect 367017 183583 367051 193137
rect 259653 172567 259687 173893
rect 232329 144959 232363 154513
rect 245853 154479 245887 162809
rect 265173 161483 265207 179333
rect 284677 162911 284711 180761
rect 285965 175967 285999 180761
rect 288725 177871 288759 180761
rect 337117 178755 337151 183481
rect 245945 143599 245979 153153
rect 250361 151827 250395 161381
rect 272073 154547 272107 162809
rect 289093 160123 289127 169677
rect 324605 162911 324639 172465
rect 359013 169779 359047 179333
rect 375849 173927 375883 183481
rect 424057 176579 424091 183413
rect 302525 153255 302559 162809
rect 360301 161483 360335 171037
rect 362233 161483 362267 171037
rect 266645 144891 266679 153153
rect 232329 125715 232363 143497
rect 244473 137955 244507 143497
rect 249993 132515 250027 142069
rect 251465 133943 251499 137989
rect 259653 132515 259687 142069
rect 270969 135099 271003 143497
rect 273545 137955 273579 144857
rect 286057 132515 286091 142069
rect 288817 140811 288851 150365
rect 310805 147611 310839 153153
rect 337117 143599 337151 153153
rect 359105 151827 359139 161381
rect 372813 157335 372847 164169
rect 375849 154615 375883 164169
rect 421205 153255 421239 162809
rect 232329 114563 232363 124117
rect 249993 114563 250027 124117
rect 272165 114563 272199 124117
rect 273545 115991 273579 125545
rect 284677 122859 284711 132413
rect 291577 120139 291611 137921
rect 295717 131155 295751 140709
rect 296913 132515 296947 142069
rect 306757 129931 306791 132413
rect 310805 128299 310839 138669
rect 327273 135235 327307 143497
rect 267841 113135 267875 114461
rect 232329 95251 232363 104805
rect 268025 103615 268059 113101
rect 251465 96679 251499 99365
rect 232237 75939 232271 85493
rect 251465 77299 251499 86921
rect 266645 85595 266679 95149
rect 267841 93891 267875 103445
rect 272441 93891 272475 103445
rect 273545 99331 273579 106233
rect 291485 103547 291519 115209
rect 306849 111843 306883 121261
rect 310805 114631 310839 125477
rect 337209 124219 337243 133841
rect 357449 128231 357483 135201
rect 358737 133943 358771 143497
rect 367017 135303 367051 144857
rect 372721 135303 372755 138125
rect 375849 135303 375883 144857
rect 421205 133943 421239 143497
rect 310805 104907 310839 114461
rect 324605 113203 324639 120581
rect 330585 111775 330619 120037
rect 339785 115991 339819 118745
rect 341165 118643 341199 125545
rect 358737 114563 358771 124117
rect 367017 115991 367051 125545
rect 389465 122859 389499 133841
rect 284769 93891 284803 95149
rect 288725 92531 288759 102085
rect 302617 95251 302651 104805
rect 323409 95251 323443 104805
rect 324605 95251 324639 104805
rect 327181 98719 327215 103445
rect 330217 102187 330251 106709
rect 377045 106335 377079 115889
rect 421205 114563 421239 124117
rect 358737 104975 358771 106301
rect 291393 88995 291427 93789
rect 310805 85595 310839 95149
rect 266737 74579 266771 84133
rect 267749 74579 267783 84133
rect 272165 67643 272199 72437
rect 232237 48331 232271 66181
rect 236285 57987 236319 67541
rect 250085 60707 250119 66181
rect 250085 48331 250119 50949
rect 234997 37315 235031 46869
rect 236285 37315 236319 48229
rect 265265 46971 265299 66181
rect 266645 48331 266679 61421
rect 267749 55267 267783 64821
rect 273637 57987 273671 67541
rect 284677 66283 284711 84133
rect 285965 66283 285999 84133
rect 288725 75803 288759 84133
rect 289921 74579 289955 84133
rect 297005 74579 297039 84133
rect 301237 75871 301271 77333
rect 306757 75803 306791 84133
rect 317705 75939 317739 85493
rect 330125 82943 330159 97257
rect 337209 95251 337243 104805
rect 339417 95251 339451 103445
rect 358645 95251 358679 104805
rect 375849 97835 375883 106233
rect 377137 99331 377171 106233
rect 424517 104907 424551 114461
rect 341073 77299 341107 86921
rect 362325 85595 362359 95149
rect 367017 87023 367051 96577
rect 389373 87907 389407 99161
rect 421205 87023 421239 104805
rect 296821 64923 296855 74409
rect 310805 66351 310839 75837
rect 330217 69955 330251 75837
rect 341073 70295 341107 77129
rect 360209 75939 360243 85493
rect 357633 66283 357667 70465
rect 389373 67643 389407 77197
rect 421021 75939 421055 85493
rect 284677 48331 284711 57001
rect 267841 45611 267875 45917
rect 239137 37315 239171 41293
rect 244381 28067 244415 37213
rect 245853 27659 245887 37213
rect 265265 35955 265299 45509
rect 273545 38675 273579 48229
rect 286057 46971 286091 56525
rect 294245 55267 294279 64821
rect 310805 60027 310839 66181
rect 301053 51799 301087 57885
rect 306757 52003 306791 59993
rect 323317 48331 323351 61421
rect 325985 48195 326019 66181
rect 327181 56627 327215 66181
rect 336933 56627 336967 66181
rect 337301 46971 337335 56525
rect 339785 48331 339819 57885
rect 359105 56559 359139 64821
rect 362233 55267 362267 64821
rect 367017 48331 367051 57885
rect 389189 48331 389223 57885
rect 421113 56695 421147 66181
rect 421021 46971 421055 56525
rect 424517 48331 424551 53805
rect 470609 48331 470643 57885
rect 296821 38607 296855 45509
rect 301329 35955 301363 45509
rect 303813 32419 303847 40137
rect 307033 35955 307067 45509
rect 327273 37315 327307 46869
rect 330125 37315 330159 46869
rect 336933 37315 336967 46869
rect 341257 37315 341291 46869
rect 358645 37315 358679 46869
rect 359105 37315 359139 46869
rect 362233 38607 362267 41429
rect 377137 38743 377171 41293
rect 236285 18003 236319 27557
rect 244197 16643 244231 26197
rect 245853 16643 245887 26197
rect 265265 19295 265299 27557
rect 267749 10659 267783 26197
rect 284585 18003 284619 27557
rect 285965 18003 285999 27557
rect 288817 19295 288851 29801
rect 337117 27659 337151 37213
rect 367017 29087 367051 38573
rect 273453 10931 273487 17901
rect 299765 16643 299799 26197
rect 295625 12223 295659 12461
rect 330217 7803 330251 9605
rect 336933 8075 336967 9605
rect 227545 6987 227579 7633
rect 321569 4947 321603 5049
rect 327181 4947 327215 5049
rect 321569 4913 321753 4947
rect 327031 4913 327215 4947
rect 224233 4811 224267 4913
rect 224141 4267 224175 4777
rect 337117 4607 337151 11169
rect 341257 9707 341291 26197
rect 358553 9707 358587 27557
rect 367017 19363 367051 28917
rect 389465 19363 389499 28917
rect 421205 27659 421239 42041
rect 424517 29019 424551 38573
rect 362233 8347 362267 18037
rect 366925 10115 366959 19261
rect 376769 8347 376803 17901
rect 421205 9707 421239 22729
rect 45477 3179 45511 3349
rect 82921 2975 82955 3145
rect 93869 2839 93903 2941
rect 264621 1139 264655 4029
rect 278053 3859 278087 4097
rect 282929 3723 282963 4029
rect 287621 3995 287655 4165
rect 354873 4131 354907 4369
rect 287713 3723 287747 3961
rect 332333 3927 332367 4097
rect 273269 3043 273303 3213
rect 282837 3043 282871 3349
rect 288633 3315 288667 3825
rect 292497 3315 292531 3689
rect 320649 3451 320683 3621
rect 320833 3587 320867 3893
rect 326353 3723 326387 3893
rect 332241 3791 332275 3893
rect 332149 3587 332183 3757
rect 335369 3587 335403 4097
rect 336197 3723 336231 3893
rect 322765 3111 322799 3553
rect 335921 3043 335955 3553
rect 335461 3009 335679 3043
rect 336013 3145 336105 3179
rect 340647 3145 340831 3179
rect 335461 2839 335495 3009
rect 335645 2975 335679 3009
rect 336013 2975 336047 3145
rect 335645 2941 336047 2975
rect 335553 2839 335587 2941
rect 340797 2907 340831 3145
rect 341257 2839 341291 4097
rect 341441 2975 341475 3349
rect 341349 2839 341383 2941
rect 345581 2839 345615 3213
rect 345673 3179 345707 3349
rect 349169 3247 349203 4097
rect 356069 4131 356103 4369
rect 352021 2907 352055 4097
rect 352205 3655 352239 3961
rect 352113 2907 352147 3621
rect 352389 3247 352423 4029
rect 376769 3927 376803 5049
rect 355057 3689 355551 3723
rect 355057 3655 355091 3689
rect 355517 3655 355551 3689
rect 355425 3451 355459 3621
rect 376861 3519 376895 4913
rect 376803 3485 376895 3519
rect 352941 3247 352975 3349
rect 370329 3315 370363 3417
rect 369903 3281 370363 3315
rect 364993 3111 365027 3281
rect 355517 2771 355551 3077
rect 355609 2907 355643 3077
rect 360301 2975 360335 3009
rect 360301 2941 360485 2975
rect 389465 595 389499 9605
rect 461225 4879 461259 5117
rect 466101 4947 466135 5253
rect 471345 4811 471379 5049
rect 471437 4811 471471 5525
rect 414029 3791 414063 4097
rect 413201 3043 413235 3485
rect 422861 2839 422895 3689
rect 425253 3655 425287 3961
rect 431233 3043 431267 3621
rect 422953 2907 422987 3009
rect 431877 2839 431911 3689
rect 433901 3247 433935 3349
rect 441629 3247 441663 3689
rect 441721 3655 441755 3893
rect 445493 3859 445527 4097
rect 443101 3655 443135 3757
rect 446321 3247 446355 4029
rect 446505 3383 446539 3621
rect 446413 2839 446447 3349
rect 446689 3315 446723 3757
rect 451933 2975 451967 3825
rect 466101 3825 466377 3859
rect 451231 2873 451381 2907
rect 451841 2839 451875 2941
rect 456809 2907 456843 3689
rect 457177 2907 457211 3621
rect 466101 3587 466135 3825
rect 466227 3485 466319 3519
rect 461593 2907 461627 3009
rect 466285 2907 466319 3485
rect 466285 2873 466377 2907
rect 471529 595 471563 5593
rect 518173 3043 518207 3213
<< viali >>
rect 364533 685797 364567 685831
rect 364533 676209 364567 676243
rect 429577 684437 429611 684471
rect 559297 684437 559331 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 364533 618205 364567 618239
rect 364533 608617 364567 608651
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 364625 598893 364659 598927
rect 364625 589305 364659 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 247969 579309 248003 579343
rect 254225 579309 254259 579343
rect 292129 579309 292163 579343
rect 292129 579105 292163 579139
rect 415685 579309 415719 579343
rect 254225 578629 254259 578663
rect 247969 578561 248003 578595
rect 415685 578493 415719 578527
rect 428381 579309 428415 579343
rect 428381 578425 428415 578459
rect 441077 579309 441111 579343
rect 441077 578357 441111 578391
rect 453589 579309 453623 579343
rect 453589 578289 453623 578323
rect 455797 579309 455831 579343
rect 455797 578221 455831 578255
rect 238769 338657 238803 338691
rect 229109 338113 229143 338147
rect 86969 338045 87003 338079
rect 87245 338045 87279 338079
rect 87061 337909 87095 337943
rect 87245 337909 87279 337943
rect 87061 337773 87095 337807
rect 87245 337773 87279 337807
rect 238677 338113 238711 338147
rect 229109 337705 229143 337739
rect 87061 337637 87095 337671
rect 87429 337637 87463 337671
rect 115673 337569 115707 337603
rect 115857 337569 115891 337603
rect 134993 337569 135027 337603
rect 135177 337569 135211 337603
rect 154313 337569 154347 337603
rect 154497 337569 154531 337603
rect 173633 337569 173667 337603
rect 173817 337569 173851 337603
rect 192953 337569 192987 337603
rect 193137 337569 193171 337603
rect 212273 337569 212307 337603
rect 212457 337569 212491 337603
rect 220921 337569 220955 337603
rect 221105 337569 221139 337603
rect 230489 337501 230523 337535
rect 230581 337637 230615 337671
rect 231225 337637 231259 337671
rect 234445 337637 234479 337671
rect 238677 337637 238711 337671
rect 346409 338657 346443 338691
rect 327089 338113 327123 338147
rect 315497 338045 315531 338079
rect 318901 338045 318935 338079
rect 319085 338045 319119 338079
rect 302157 337773 302191 337807
rect 302249 337705 302283 337739
rect 303997 337773 304031 337807
rect 238769 337637 238803 337671
rect 259745 337637 259779 337671
rect 230581 337501 230615 337535
rect 87061 337433 87095 337467
rect 87153 337433 87187 337467
rect 220921 337433 220955 337467
rect 221105 337433 221139 337467
rect 234445 337433 234479 337467
rect 259745 337365 259779 337399
rect 220921 337297 220955 337331
rect 221105 337297 221139 337331
rect 103437 337229 103471 337263
rect 86969 337093 87003 337127
rect 86969 336957 87003 336991
rect 103437 336957 103471 336991
rect 113189 337229 113223 337263
rect 113189 336753 113223 336787
rect 122757 337229 122791 337263
rect 220829 337229 220863 337263
rect 221013 337229 221047 337263
rect 318901 337909 318935 337943
rect 318993 337909 319027 337943
rect 318809 337773 318843 337807
rect 318993 337773 319027 337807
rect 336657 338113 336691 338147
rect 327089 337705 327123 337739
rect 335921 337841 335955 337875
rect 318901 337569 318935 337603
rect 318993 337569 319027 337603
rect 335829 337501 335863 337535
rect 318809 337433 318843 337467
rect 319085 337433 319119 337467
rect 334725 337365 334759 337399
rect 315497 337297 315531 337331
rect 326353 337297 326387 337331
rect 303997 337161 304031 337195
rect 326353 337161 326387 337195
rect 122757 336753 122791 336787
rect 336013 337841 336047 337875
rect 336657 337705 336691 337739
rect 346409 337705 346443 337739
rect 365177 338113 365211 338147
rect 336013 337637 336047 337671
rect 344661 337637 344695 337671
rect 364993 337637 365027 337671
rect 341717 337501 341751 337535
rect 335921 337365 335955 337399
rect 336197 337365 336231 337399
rect 335829 337025 335863 337059
rect 340797 337365 340831 337399
rect 340797 337093 340831 337127
rect 340889 337365 340923 337399
rect 336197 336889 336231 336923
rect 340613 337025 340647 337059
rect 334725 336753 334759 336787
rect 341717 337229 341751 337263
rect 342821 337501 342855 337535
rect 344201 337501 344235 337535
rect 342821 337161 342855 337195
rect 345581 337365 345615 337399
rect 354045 337365 354079 337399
rect 345857 337161 345891 337195
rect 345857 336957 345891 336991
rect 466377 338113 466411 338147
rect 365177 337569 365211 337603
rect 374653 338045 374687 338079
rect 376769 338045 376803 338079
rect 451473 337977 451507 338011
rect 441629 337909 441663 337943
rect 376769 337637 376803 337671
rect 412557 337841 412591 337875
rect 374653 337569 374687 337603
rect 412557 337569 412591 337603
rect 414121 337705 414155 337739
rect 365085 337501 365119 337535
rect 365269 337501 365303 337535
rect 432245 337705 432279 337739
rect 374653 337433 374687 337467
rect 414121 337433 414155 337467
rect 422953 337433 422987 337467
rect 364993 337161 365027 337195
rect 369869 337365 369903 337399
rect 369869 337161 369903 337195
rect 422953 337229 422987 337263
rect 374653 337161 374687 337195
rect 427921 337161 427955 337195
rect 354045 336957 354079 336991
rect 345581 336889 345615 336923
rect 437397 337569 437431 337603
rect 437581 337569 437615 337603
rect 436753 337365 436787 337399
rect 436753 337093 436787 337127
rect 432245 336957 432279 336991
rect 427921 336889 427955 336923
rect 451105 337909 451139 337943
rect 446413 337773 446447 337807
rect 446413 337501 446447 337535
rect 448529 337773 448563 337807
rect 448529 337501 448563 337535
rect 449173 337705 449207 337739
rect 449173 337365 449207 337399
rect 340889 336821 340923 336855
rect 345489 336821 345523 336855
rect 345765 336821 345799 336855
rect 441629 336821 441663 336855
rect 451105 336821 451139 336855
rect 451289 337909 451323 337943
rect 461593 337977 461627 338011
rect 451473 337841 451507 337875
rect 461409 337841 461443 337875
rect 451381 337705 451415 337739
rect 456993 337569 457027 337603
rect 451381 337365 451415 337399
rect 456073 337501 456107 337535
rect 456073 337365 456107 337399
rect 456993 337297 457027 337331
rect 459109 337569 459143 337603
rect 340797 336753 340831 336787
rect 340981 336753 341015 336787
rect 341165 336753 341199 336787
rect 451289 336753 451323 336787
rect 457177 337229 457211 337263
rect 461593 337773 461627 337807
rect 466285 337977 466319 338011
rect 466377 337977 466411 338011
rect 460397 337501 460431 337535
rect 461409 337501 461443 337535
rect 460397 337229 460431 337263
rect 461593 337297 461627 337331
rect 459109 336821 459143 336855
rect 461593 336821 461627 336855
rect 457177 336753 457211 336787
rect 469229 337909 469263 337943
rect 466469 337297 466503 337331
rect 469229 337229 469263 337263
rect 470793 337365 470827 337399
rect 466469 336889 466503 336923
rect 470793 336889 470827 336923
rect 480913 337365 480947 337399
rect 489929 337365 489963 337399
rect 489929 337093 489963 337127
rect 500233 337365 500267 337399
rect 500233 337093 500267 337127
rect 480913 336889 480947 336923
rect 284401 336685 284435 336719
rect 265265 335257 265299 335291
rect 250177 334441 250211 334475
rect 250177 327097 250211 327131
rect 259837 328389 259871 328423
rect 236469 321657 236503 321691
rect 236469 318801 236503 318835
rect 284401 335189 284435 335223
rect 288817 336685 288851 336719
rect 270785 334305 270819 334339
rect 270785 328457 270819 328491
rect 272257 334305 272291 334339
rect 272257 328457 272291 328491
rect 265265 325669 265299 325703
rect 273545 327029 273579 327063
rect 273545 321521 273579 321555
rect 285965 327029 285999 327063
rect 259837 318801 259871 318835
rect 327273 336685 327307 336719
rect 302617 328389 302651 328423
rect 337393 336685 337427 336719
rect 337393 328389 337427 328423
rect 339785 336685 339819 336719
rect 466285 336685 466319 336719
rect 327273 327097 327307 327131
rect 302617 318801 302651 318835
rect 330125 327029 330159 327063
rect 330125 318801 330159 318835
rect 337393 321589 337427 321623
rect 337393 318801 337427 318835
rect 339785 318801 339819 318835
rect 341349 328389 341383 328423
rect 341349 318801 341383 318835
rect 389465 328389 389499 328423
rect 389465 318801 389499 318835
rect 470609 328389 470643 328423
rect 470609 318801 470643 318835
rect 288817 318597 288851 318631
rect 372721 318733 372755 318767
rect 285965 317509 285999 317543
rect 306757 317441 306791 317475
rect 250177 317373 250211 317407
rect 239137 309077 239171 309111
rect 232329 307717 232363 307751
rect 250177 307785 250211 307819
rect 251557 317373 251591 317407
rect 299765 317373 299799 317407
rect 290105 313225 290139 313259
rect 251557 307785 251591 307819
rect 284585 311865 284619 311899
rect 285965 311865 285999 311899
rect 285965 306425 285999 306459
rect 288725 308397 288759 308431
rect 284585 306357 284619 306391
rect 239137 299489 239171 299523
rect 245945 302413 245979 302447
rect 232329 298129 232363 298163
rect 236285 298061 236319 298095
rect 232237 297993 232271 298027
rect 232237 288405 232271 288439
rect 245945 297993 245979 298027
rect 250177 298061 250211 298095
rect 250177 289765 250211 289799
rect 251373 298061 251407 298095
rect 236285 288405 236319 288439
rect 273637 296633 273671 296667
rect 251373 288405 251407 288439
rect 272165 289765 272199 289799
rect 290105 306289 290139 306323
rect 306757 316013 306791 316047
rect 325893 317373 325927 317407
rect 310897 311933 310931 311967
rect 310897 307853 310931 307887
rect 372721 309145 372755 309179
rect 421205 317373 421239 317407
rect 325893 307785 325927 307819
rect 339877 309077 339911 309111
rect 310713 307717 310747 307751
rect 299765 299489 299799 299523
rect 306849 299489 306883 299523
rect 337025 307717 337059 307751
rect 310713 298129 310747 298163
rect 323317 299421 323351 299455
rect 306849 296701 306883 296735
rect 288725 289969 288759 290003
rect 310897 293029 310931 293063
rect 273637 287045 273671 287079
rect 272165 283577 272199 283611
rect 324697 299421 324731 299455
rect 339877 299897 339911 299931
rect 341165 309077 341199 309111
rect 341165 299489 341199 299523
rect 367017 309077 367051 309111
rect 367017 299489 367051 299523
rect 389281 309009 389315 309043
rect 421205 307785 421239 307819
rect 470609 309077 470643 309111
rect 389281 299489 389315 299523
rect 470609 299489 470643 299523
rect 337025 298197 337059 298231
rect 372721 299421 372755 299455
rect 324697 289833 324731 289867
rect 325985 298061 326019 298095
rect 323317 288405 323351 288439
rect 325985 288405 326019 288439
rect 327181 298061 327215 298095
rect 337209 298061 337243 298095
rect 337209 292417 337243 292451
rect 372721 289833 372755 289867
rect 421205 298061 421239 298095
rect 341165 289765 341199 289799
rect 327181 288405 327215 288439
rect 330309 288405 330343 288439
rect 330309 287045 330343 287079
rect 310897 282761 310931 282795
rect 337117 282897 337151 282931
rect 270693 280109 270727 280143
rect 270693 275281 270727 275315
rect 273545 280109 273579 280143
rect 341165 280177 341199 280211
rect 367017 289765 367051 289799
rect 367017 280177 367051 280211
rect 389373 289765 389407 289799
rect 421205 288405 421239 288439
rect 470609 289765 470643 289799
rect 389373 280177 389407 280211
rect 470609 280177 470643 280211
rect 337117 278749 337151 278783
rect 372721 280109 372755 280143
rect 232237 270521 232271 270555
rect 273545 270521 273579 270555
rect 310897 278681 310931 278715
rect 232237 269093 232271 269127
rect 324513 278681 324547 278715
rect 362233 277321 362267 277355
rect 324513 269093 324547 269127
rect 330125 277253 330159 277287
rect 310897 263449 310931 263483
rect 341165 270453 341199 270487
rect 330125 263177 330159 263211
rect 337117 263585 337151 263619
rect 306849 262905 306883 262939
rect 270693 260797 270727 260831
rect 270693 255969 270727 256003
rect 273545 260797 273579 260831
rect 250085 253929 250119 253963
rect 273545 251209 273579 251243
rect 290013 258009 290047 258043
rect 250085 249781 250119 249815
rect 259653 251141 259687 251175
rect 284677 249713 284711 249747
rect 259653 242641 259687 242675
rect 270693 244273 270727 244307
rect 270693 241553 270727 241587
rect 251373 241485 251407 241519
rect 251373 240125 251407 240159
rect 270693 241417 270727 241451
rect 244381 234821 244415 234855
rect 244381 230469 244415 230503
rect 250177 234617 250211 234651
rect 290013 248421 290047 248455
rect 294245 258009 294279 258043
rect 372721 270521 372755 270555
rect 375849 280109 375883 280143
rect 375849 270521 375883 270555
rect 377137 280109 377171 280143
rect 377137 270521 377171 270555
rect 424609 280109 424643 280143
rect 424609 270521 424643 270555
rect 362233 263449 362267 263483
rect 367017 270453 367051 270487
rect 341165 260865 341199 260899
rect 367017 260865 367051 260899
rect 389373 270453 389407 270487
rect 389373 260865 389407 260899
rect 470609 270453 470643 270487
rect 470609 260865 470643 260899
rect 337117 259437 337151 259471
rect 372721 260797 372755 260831
rect 310897 256037 310931 256071
rect 310897 251277 310931 251311
rect 323409 252705 323443 252739
rect 306849 249781 306883 249815
rect 310713 251141 310747 251175
rect 294245 248421 294279 248455
rect 291485 248353 291519 248387
rect 284677 240125 284711 240159
rect 285965 244953 285999 244987
rect 310713 241485 310747 241519
rect 372721 251209 372755 251243
rect 375849 260797 375883 260831
rect 375849 251209 375883 251243
rect 377137 260797 377171 260831
rect 377137 251209 377171 251243
rect 424517 260797 424551 260831
rect 424517 251209 424551 251243
rect 463709 260797 463743 260831
rect 463709 251209 463743 251243
rect 325893 251141 325927 251175
rect 325893 249781 325927 249815
rect 367017 251141 367051 251175
rect 323409 241485 323443 241519
rect 327181 249713 327215 249747
rect 291485 240057 291519 240091
rect 299489 241417 299523 241451
rect 285965 234481 285999 234515
rect 270693 232033 270727 232067
rect 250177 230469 250211 230503
rect 266737 231897 266771 231931
rect 367017 241485 367051 241519
rect 470609 251141 470643 251175
rect 470609 241485 470643 241519
rect 327181 240193 327215 240227
rect 362233 241417 362267 241451
rect 327181 240057 327215 240091
rect 323409 234685 323443 234719
rect 299489 231829 299523 231863
rect 302617 231965 302651 231999
rect 266737 230469 266771 230503
rect 302617 230469 302651 230503
rect 310805 231761 310839 231795
rect 323409 231761 323443 231795
rect 270693 224961 270727 224995
rect 270693 222241 270727 222275
rect 327181 230537 327215 230571
rect 375849 241417 375883 241451
rect 389281 241417 389315 241451
rect 389281 234617 389315 234651
rect 375849 231829 375883 231863
rect 362233 230469 362267 230503
rect 367017 231761 367051 231795
rect 310805 222173 310839 222207
rect 367017 222173 367051 222207
rect 270693 222105 270727 222139
rect 244473 217957 244507 217991
rect 232237 211225 232271 211259
rect 232237 209797 232271 209831
rect 270693 212721 270727 212755
rect 299489 222105 299523 222139
rect 375849 222105 375883 222139
rect 341165 220745 341199 220779
rect 272165 212517 272199 212551
rect 299489 212517 299523 212551
rect 330125 219385 330159 219419
rect 272165 211157 272199 211191
rect 310805 212449 310839 212483
rect 265265 211089 265299 211123
rect 341165 215237 341199 215271
rect 362141 215305 362175 215339
rect 375849 212517 375883 212551
rect 362141 211157 362175 211191
rect 330125 209797 330159 209831
rect 310805 202861 310839 202895
rect 330217 209729 330251 209763
rect 265265 202725 265299 202759
rect 299489 202793 299523 202827
rect 330217 202793 330251 202827
rect 336933 202793 336967 202827
rect 244473 200141 244507 200175
rect 291485 200073 291519 200107
rect 284677 198645 284711 198679
rect 244381 186949 244415 186983
rect 267749 186337 267783 186371
rect 267749 183549 267783 183583
rect 270693 186337 270727 186371
rect 270693 183549 270727 183583
rect 299489 193205 299523 193239
rect 375849 202793 375883 202827
rect 336933 193205 336967 193239
rect 358645 201433 358679 201467
rect 362233 198033 362267 198067
rect 362233 193205 362267 193239
rect 375849 193205 375883 193239
rect 358645 191845 358679 191879
rect 367017 193137 367051 193171
rect 291485 190485 291519 190519
rect 299857 188445 299891 188479
rect 299857 183549 299891 183583
rect 306849 188445 306883 188479
rect 306849 183549 306883 183583
rect 367017 183549 367051 183583
rect 284677 183481 284711 183515
rect 337117 183481 337151 183515
rect 244381 180829 244415 180863
rect 284677 180761 284711 180795
rect 265173 179333 265207 179367
rect 259653 173893 259687 173927
rect 259653 172533 259687 172567
rect 245853 162809 245887 162843
rect 232329 154513 232363 154547
rect 285965 180761 285999 180795
rect 288725 180761 288759 180795
rect 375849 183481 375883 183515
rect 337117 178721 337151 178755
rect 359013 179333 359047 179367
rect 288725 177837 288759 177871
rect 285965 175933 285999 175967
rect 324605 172465 324639 172499
rect 284677 162877 284711 162911
rect 289093 169677 289127 169711
rect 265173 161449 265207 161483
rect 272073 162809 272107 162843
rect 245853 154445 245887 154479
rect 250361 161381 250395 161415
rect 232329 144925 232363 144959
rect 245945 153153 245979 153187
rect 424057 183413 424091 183447
rect 424057 176545 424091 176579
rect 375849 173893 375883 173927
rect 359013 169745 359047 169779
rect 360301 171037 360335 171071
rect 324605 162877 324639 162911
rect 289093 160089 289127 160123
rect 302525 162809 302559 162843
rect 272073 154513 272107 154547
rect 360301 161449 360335 161483
rect 362233 171037 362267 171071
rect 362233 161449 362267 161483
rect 372813 164169 372847 164203
rect 302525 153221 302559 153255
rect 359105 161381 359139 161415
rect 250361 151793 250395 151827
rect 266645 153153 266679 153187
rect 310805 153153 310839 153187
rect 288817 150365 288851 150399
rect 266645 144857 266679 144891
rect 273545 144857 273579 144891
rect 245945 143565 245979 143599
rect 232329 143497 232363 143531
rect 244473 143497 244507 143531
rect 270969 143497 271003 143531
rect 244473 137921 244507 137955
rect 249993 142069 250027 142103
rect 259653 142069 259687 142103
rect 251465 137989 251499 138023
rect 251465 133909 251499 133943
rect 249993 132481 250027 132515
rect 273545 137921 273579 137955
rect 286057 142069 286091 142103
rect 270969 135065 271003 135099
rect 259653 132481 259687 132515
rect 310805 147577 310839 147611
rect 337117 153153 337151 153187
rect 372813 157301 372847 157335
rect 375849 164169 375883 164203
rect 375849 154581 375883 154615
rect 421205 162809 421239 162843
rect 421205 153221 421239 153255
rect 359105 151793 359139 151827
rect 337117 143565 337151 143599
rect 367017 144857 367051 144891
rect 327273 143497 327307 143531
rect 288817 140777 288851 140811
rect 296913 142069 296947 142103
rect 295717 140709 295751 140743
rect 286057 132481 286091 132515
rect 291577 137921 291611 137955
rect 232329 125681 232363 125715
rect 284677 132413 284711 132447
rect 273545 125545 273579 125579
rect 232329 124117 232363 124151
rect 232329 114529 232363 114563
rect 249993 124117 250027 124151
rect 249993 114529 250027 114563
rect 272165 124117 272199 124151
rect 284677 122825 284711 122859
rect 296913 132481 296947 132515
rect 310805 138669 310839 138703
rect 295717 131121 295751 131155
rect 306757 132413 306791 132447
rect 306757 129897 306791 129931
rect 358737 143497 358771 143531
rect 327273 135201 327307 135235
rect 357449 135201 357483 135235
rect 310805 128265 310839 128299
rect 337209 133841 337243 133875
rect 310805 125477 310839 125511
rect 291577 120105 291611 120139
rect 306849 121261 306883 121295
rect 273545 115957 273579 115991
rect 272165 114529 272199 114563
rect 291485 115209 291519 115243
rect 267841 114461 267875 114495
rect 267841 113101 267875 113135
rect 268025 113101 268059 113135
rect 232329 104805 232363 104839
rect 268025 103581 268059 103615
rect 273545 106233 273579 106267
rect 267841 103445 267875 103479
rect 251465 99365 251499 99399
rect 251465 96645 251499 96679
rect 232329 95217 232363 95251
rect 266645 95149 266679 95183
rect 251465 86921 251499 86955
rect 232237 85493 232271 85527
rect 267841 93857 267875 93891
rect 272441 103445 272475 103479
rect 375849 144857 375883 144891
rect 367017 135269 367051 135303
rect 372721 138125 372755 138159
rect 372721 135269 372755 135303
rect 375849 135269 375883 135303
rect 421205 143497 421239 143531
rect 358737 133909 358771 133943
rect 421205 133909 421239 133943
rect 357449 128197 357483 128231
rect 389465 133841 389499 133875
rect 337209 124185 337243 124219
rect 341165 125545 341199 125579
rect 310805 114597 310839 114631
rect 324605 120581 324639 120615
rect 306849 111809 306883 111843
rect 310805 114461 310839 114495
rect 324605 113169 324639 113203
rect 330585 120037 330619 120071
rect 339785 118745 339819 118779
rect 367017 125545 367051 125579
rect 341165 118609 341199 118643
rect 358737 124117 358771 124151
rect 339785 115957 339819 115991
rect 389465 122825 389499 122859
rect 421205 124117 421239 124151
rect 367017 115957 367051 115991
rect 358737 114529 358771 114563
rect 377045 115889 377079 115923
rect 330585 111741 330619 111775
rect 310805 104873 310839 104907
rect 330217 106709 330251 106743
rect 291485 103513 291519 103547
rect 302617 104805 302651 104839
rect 273545 99297 273579 99331
rect 288725 102085 288759 102119
rect 272441 93857 272475 93891
rect 284769 95149 284803 95183
rect 284769 93857 284803 93891
rect 302617 95217 302651 95251
rect 323409 104805 323443 104839
rect 323409 95217 323443 95251
rect 324605 104805 324639 104839
rect 327181 103445 327215 103479
rect 421205 114529 421239 114563
rect 358737 106301 358771 106335
rect 377045 106301 377079 106335
rect 424517 114461 424551 114495
rect 358737 104941 358771 104975
rect 375849 106233 375883 106267
rect 330217 102153 330251 102187
rect 337209 104805 337243 104839
rect 327181 98685 327215 98719
rect 324605 95217 324639 95251
rect 330125 97257 330159 97291
rect 310805 95149 310839 95183
rect 288725 92497 288759 92531
rect 291393 93789 291427 93823
rect 291393 88961 291427 88995
rect 266645 85561 266679 85595
rect 310805 85561 310839 85595
rect 317705 85493 317739 85527
rect 251465 77265 251499 77299
rect 266737 84133 266771 84167
rect 232237 75905 232271 75939
rect 266737 74545 266771 74579
rect 267749 84133 267783 84167
rect 267749 74545 267783 74579
rect 284677 84133 284711 84167
rect 272165 72437 272199 72471
rect 272165 67609 272199 67643
rect 236285 67541 236319 67575
rect 232237 66181 232271 66215
rect 273637 67541 273671 67575
rect 250085 66181 250119 66215
rect 250085 60673 250119 60707
rect 265265 66181 265299 66215
rect 236285 57953 236319 57987
rect 232237 48297 232271 48331
rect 250085 50949 250119 50983
rect 250085 48297 250119 48331
rect 236285 48229 236319 48263
rect 234997 46869 235031 46903
rect 234997 37281 235031 37315
rect 267749 64821 267783 64855
rect 266645 61421 266679 61455
rect 284677 66249 284711 66283
rect 285965 84133 285999 84167
rect 288725 84133 288759 84167
rect 288725 75769 288759 75803
rect 289921 84133 289955 84167
rect 289921 74545 289955 74579
rect 297005 84133 297039 84167
rect 306757 84133 306791 84167
rect 301237 77333 301271 77367
rect 301237 75837 301271 75871
rect 358645 104805 358679 104839
rect 337209 95217 337243 95251
rect 339417 103445 339451 103479
rect 339417 95217 339451 95251
rect 377137 106233 377171 106267
rect 424517 104873 424551 104907
rect 377137 99297 377171 99331
rect 421205 104805 421239 104839
rect 375849 97801 375883 97835
rect 389373 99161 389407 99195
rect 358645 95217 358679 95251
rect 367017 96577 367051 96611
rect 362325 95149 362359 95183
rect 330125 82909 330159 82943
rect 341073 86921 341107 86955
rect 389373 87873 389407 87907
rect 367017 86989 367051 87023
rect 421205 86989 421239 87023
rect 362325 85561 362359 85595
rect 341073 77265 341107 77299
rect 360209 85493 360243 85527
rect 317705 75905 317739 75939
rect 341073 77129 341107 77163
rect 306757 75769 306791 75803
rect 310805 75837 310839 75871
rect 297005 74545 297039 74579
rect 285965 66249 285999 66283
rect 296821 74409 296855 74443
rect 330217 75837 330251 75871
rect 421021 85493 421055 85527
rect 360209 75905 360243 75939
rect 389373 77197 389407 77231
rect 341073 70261 341107 70295
rect 357633 70465 357667 70499
rect 330217 69921 330251 69955
rect 310805 66317 310839 66351
rect 421021 75905 421055 75939
rect 389373 67609 389407 67643
rect 357633 66249 357667 66283
rect 296821 64889 296855 64923
rect 310805 66181 310839 66215
rect 273637 57953 273671 57987
rect 294245 64821 294279 64855
rect 267749 55233 267783 55267
rect 284677 57001 284711 57035
rect 266645 48297 266679 48331
rect 284677 48297 284711 48331
rect 286057 56525 286091 56559
rect 265265 46937 265299 46971
rect 273545 48229 273579 48263
rect 267841 45917 267875 45951
rect 267841 45577 267875 45611
rect 265265 45509 265299 45543
rect 236285 37281 236319 37315
rect 239137 41293 239171 41327
rect 239137 37281 239171 37315
rect 244381 37213 244415 37247
rect 244381 28033 244415 28067
rect 245853 37213 245887 37247
rect 325985 66181 326019 66215
rect 306757 59993 306791 60027
rect 310805 59993 310839 60027
rect 323317 61421 323351 61455
rect 294245 55233 294279 55267
rect 301053 57885 301087 57919
rect 306757 51969 306791 52003
rect 301053 51765 301087 51799
rect 323317 48297 323351 48331
rect 327181 66181 327215 66215
rect 327181 56593 327215 56627
rect 336933 66181 336967 66215
rect 421113 66181 421147 66215
rect 359105 64821 359139 64855
rect 336933 56593 336967 56627
rect 339785 57885 339819 57919
rect 325985 48161 326019 48195
rect 337301 56525 337335 56559
rect 286057 46937 286091 46971
rect 359105 56525 359139 56559
rect 362233 64821 362267 64855
rect 362233 55233 362267 55267
rect 367017 57885 367051 57919
rect 339785 48297 339819 48331
rect 367017 48297 367051 48331
rect 389189 57885 389223 57919
rect 421113 56661 421147 56695
rect 470609 57885 470643 57919
rect 389189 48297 389223 48331
rect 421021 56525 421055 56559
rect 337301 46937 337335 46971
rect 424517 53805 424551 53839
rect 424517 48297 424551 48331
rect 470609 48297 470643 48331
rect 421021 46937 421055 46971
rect 327273 46869 327307 46903
rect 273545 38641 273579 38675
rect 296821 45509 296855 45543
rect 296821 38573 296855 38607
rect 301329 45509 301363 45543
rect 265265 35921 265299 35955
rect 307033 45509 307067 45543
rect 301329 35921 301363 35955
rect 303813 40137 303847 40171
rect 327273 37281 327307 37315
rect 330125 46869 330159 46903
rect 330125 37281 330159 37315
rect 336933 46869 336967 46903
rect 336933 37281 336967 37315
rect 341257 46869 341291 46903
rect 341257 37281 341291 37315
rect 358645 46869 358679 46903
rect 358645 37281 358679 37315
rect 359105 46869 359139 46903
rect 421205 42041 421239 42075
rect 362233 41429 362267 41463
rect 377137 41293 377171 41327
rect 377137 38709 377171 38743
rect 362233 38573 362267 38607
rect 367017 38573 367051 38607
rect 359105 37281 359139 37315
rect 307033 35921 307067 35955
rect 337117 37213 337151 37247
rect 303813 32385 303847 32419
rect 245853 27625 245887 27659
rect 288817 29801 288851 29835
rect 236285 27557 236319 27591
rect 265265 27557 265299 27591
rect 236285 17969 236319 18003
rect 244197 26197 244231 26231
rect 244197 16609 244231 16643
rect 245853 26197 245887 26231
rect 284585 27557 284619 27591
rect 265265 19261 265299 19295
rect 267749 26197 267783 26231
rect 245853 16609 245887 16643
rect 284585 17969 284619 18003
rect 285965 27557 285999 27591
rect 367017 29053 367051 29087
rect 337117 27625 337151 27659
rect 367017 28917 367051 28951
rect 358553 27557 358587 27591
rect 288817 19261 288851 19295
rect 299765 26197 299799 26231
rect 285965 17969 285999 18003
rect 273453 17901 273487 17935
rect 299765 16609 299799 16643
rect 341257 26197 341291 26231
rect 295625 12461 295659 12495
rect 295625 12189 295659 12223
rect 273453 10897 273487 10931
rect 337117 11169 337151 11203
rect 267749 10625 267783 10659
rect 330217 9605 330251 9639
rect 336933 9605 336967 9639
rect 336933 8041 336967 8075
rect 330217 7769 330251 7803
rect 227545 7633 227579 7667
rect 227545 6953 227579 6987
rect 321569 5049 321603 5083
rect 327181 5049 327215 5083
rect 224233 4913 224267 4947
rect 321753 4913 321787 4947
rect 326997 4913 327031 4947
rect 224141 4777 224175 4811
rect 224233 4777 224267 4811
rect 341257 9673 341291 9707
rect 367017 19329 367051 19363
rect 389465 28917 389499 28951
rect 424517 38573 424551 38607
rect 424517 28985 424551 29019
rect 421205 27625 421239 27659
rect 389465 19329 389499 19363
rect 421205 22729 421239 22763
rect 366925 19261 366959 19295
rect 358553 9673 358587 9707
rect 362233 18037 362267 18071
rect 366925 10081 366959 10115
rect 376769 17901 376803 17935
rect 362233 8313 362267 8347
rect 421205 9673 421239 9707
rect 376769 8313 376803 8347
rect 389465 9605 389499 9639
rect 337117 4573 337151 4607
rect 376769 5049 376803 5083
rect 224141 4233 224175 4267
rect 354873 4369 354907 4403
rect 287621 4165 287655 4199
rect 278053 4097 278087 4131
rect 264621 4029 264655 4063
rect 45477 3349 45511 3383
rect 45477 3145 45511 3179
rect 82921 3145 82955 3179
rect 82921 2941 82955 2975
rect 93869 2941 93903 2975
rect 93869 2805 93903 2839
rect 278053 3825 278087 3859
rect 282929 4029 282963 4063
rect 332333 4097 332367 4131
rect 287621 3961 287655 3995
rect 287713 3961 287747 3995
rect 282929 3689 282963 3723
rect 320833 3893 320867 3927
rect 287713 3689 287747 3723
rect 288633 3825 288667 3859
rect 282837 3349 282871 3383
rect 273269 3213 273303 3247
rect 273269 3009 273303 3043
rect 288633 3281 288667 3315
rect 292497 3689 292531 3723
rect 320649 3621 320683 3655
rect 326353 3893 326387 3927
rect 332241 3893 332275 3927
rect 332333 3893 332367 3927
rect 335369 4097 335403 4131
rect 326353 3689 326387 3723
rect 332149 3757 332183 3791
rect 332241 3757 332275 3791
rect 320833 3553 320867 3587
rect 322765 3553 322799 3587
rect 332149 3553 332183 3587
rect 341257 4097 341291 4131
rect 336197 3893 336231 3927
rect 336197 3689 336231 3723
rect 335369 3553 335403 3587
rect 335921 3553 335955 3587
rect 320649 3417 320683 3451
rect 292497 3281 292531 3315
rect 322765 3077 322799 3111
rect 282837 3009 282871 3043
rect 335921 3009 335955 3043
rect 336105 3145 336139 3179
rect 340613 3145 340647 3179
rect 335461 2805 335495 2839
rect 335553 2941 335587 2975
rect 340797 2873 340831 2907
rect 335553 2805 335587 2839
rect 349169 4097 349203 4131
rect 341441 3349 341475 3383
rect 345673 3349 345707 3383
rect 341257 2805 341291 2839
rect 341349 2941 341383 2975
rect 341441 2941 341475 2975
rect 345581 3213 345615 3247
rect 341349 2805 341383 2839
rect 349169 3213 349203 3247
rect 352021 4097 352055 4131
rect 354873 4097 354907 4131
rect 356069 4369 356103 4403
rect 356069 4097 356103 4131
rect 345673 3145 345707 3179
rect 352389 4029 352423 4063
rect 352205 3961 352239 3995
rect 352021 2873 352055 2907
rect 352113 3621 352147 3655
rect 352205 3621 352239 3655
rect 376769 3893 376803 3927
rect 376861 4913 376895 4947
rect 355057 3621 355091 3655
rect 355425 3621 355459 3655
rect 355517 3621 355551 3655
rect 376769 3485 376803 3519
rect 355425 3417 355459 3451
rect 370329 3417 370363 3451
rect 352389 3213 352423 3247
rect 352941 3349 352975 3383
rect 352941 3213 352975 3247
rect 364993 3281 365027 3315
rect 369869 3281 369903 3315
rect 352113 2873 352147 2907
rect 355517 3077 355551 3111
rect 345581 2805 345615 2839
rect 355609 3077 355643 3111
rect 364993 3077 365027 3111
rect 360301 3009 360335 3043
rect 360485 2941 360519 2975
rect 355609 2873 355643 2907
rect 355517 2737 355551 2771
rect 264621 1105 264655 1139
rect 471529 5593 471563 5627
rect 471437 5525 471471 5559
rect 466101 5253 466135 5287
rect 461225 5117 461259 5151
rect 466101 4913 466135 4947
rect 471345 5049 471379 5083
rect 461225 4845 461259 4879
rect 471345 4777 471379 4811
rect 471437 4777 471471 4811
rect 414029 4097 414063 4131
rect 445493 4097 445527 4131
rect 414029 3757 414063 3791
rect 425253 3961 425287 3995
rect 422861 3689 422895 3723
rect 413201 3485 413235 3519
rect 413201 3009 413235 3043
rect 441721 3893 441755 3927
rect 431877 3689 431911 3723
rect 425253 3621 425287 3655
rect 431233 3621 431267 3655
rect 422953 3009 422987 3043
rect 431233 3009 431267 3043
rect 422953 2873 422987 2907
rect 422861 2805 422895 2839
rect 441629 3689 441663 3723
rect 433901 3349 433935 3383
rect 433901 3213 433935 3247
rect 445493 3825 445527 3859
rect 446321 4029 446355 4063
rect 441721 3621 441755 3655
rect 443101 3757 443135 3791
rect 443101 3621 443135 3655
rect 441629 3213 441663 3247
rect 451933 3825 451967 3859
rect 446689 3757 446723 3791
rect 446505 3621 446539 3655
rect 446321 3213 446355 3247
rect 446413 3349 446447 3383
rect 446505 3349 446539 3383
rect 431877 2805 431911 2839
rect 446689 3281 446723 3315
rect 466377 3825 466411 3859
rect 451841 2941 451875 2975
rect 451933 2941 451967 2975
rect 456809 3689 456843 3723
rect 451197 2873 451231 2907
rect 451381 2873 451415 2907
rect 446413 2805 446447 2839
rect 456809 2873 456843 2907
rect 457177 3621 457211 3655
rect 466101 3553 466135 3587
rect 466193 3485 466227 3519
rect 457177 2873 457211 2907
rect 461593 3009 461627 3043
rect 461593 2873 461627 2907
rect 466377 2873 466411 2907
rect 451841 2805 451875 2839
rect 389465 561 389499 595
rect 518173 3213 518207 3247
rect 518173 3009 518207 3043
rect 471529 561 471563 595
<< metal1 >>
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 358814 700992 358820 701004
rect 202840 700964 358820 700992
rect 202840 700952 202846 700964
rect 358814 700952 358820 700964
rect 358872 700952 358878 701004
rect 170306 700884 170312 700936
rect 170364 700924 170370 700936
rect 362954 700924 362960 700936
rect 170364 700896 362960 700924
rect 170364 700884 170370 700896
rect 362954 700884 362960 700896
rect 363012 700884 363018 700936
rect 328362 700816 328368 700868
rect 328420 700856 328426 700868
rect 527174 700856 527180 700868
rect 328420 700828 527180 700856
rect 328420 700816 328426 700828
rect 527174 700816 527180 700828
rect 527232 700816 527238 700868
rect 329742 700748 329748 700800
rect 329800 700788 329806 700800
rect 543458 700788 543464 700800
rect 329800 700760 543464 700788
rect 329800 700748 329806 700760
rect 543458 700748 543464 700760
rect 543516 700748 543522 700800
rect 154114 700680 154120 700732
rect 154172 700720 154178 700732
rect 367094 700720 367100 700732
rect 154172 700692 367100 700720
rect 154172 700680 154178 700692
rect 367094 700680 367100 700692
rect 367152 700680 367158 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 364334 700652 364340 700664
rect 137888 700624 364340 700652
rect 137888 700612 137894 700624
rect 364334 700612 364340 700624
rect 364392 700612 364398 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 368474 700584 368480 700596
rect 105504 700556 368480 700584
rect 105504 700544 105510 700556
rect 368474 700544 368480 700556
rect 368532 700544 368538 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 373994 700516 374000 700528
rect 89220 700488 374000 700516
rect 89220 700476 89226 700488
rect 373994 700476 374000 700488
rect 374052 700476 374058 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 371234 700448 371240 700460
rect 73028 700420 371240 700448
rect 73028 700408 73034 700420
rect 371234 700408 371240 700420
rect 371292 700408 371298 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 375374 700380 375380 700392
rect 40552 700352 375380 700380
rect 40552 700340 40558 700352
rect 375374 700340 375380 700352
rect 375432 700340 375438 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 379514 700312 379520 700324
rect 24360 700284 379520 700312
rect 24360 700272 24366 700284
rect 379514 700272 379520 700284
rect 379572 700272 379578 700324
rect 218974 700204 218980 700256
rect 219032 700244 219038 700256
rect 360194 700244 360200 700256
rect 219032 700216 360200 700244
rect 219032 700204 219038 700216
rect 360194 700204 360200 700216
rect 360252 700204 360258 700256
rect 336642 700136 336648 700188
rect 336700 700176 336706 700188
rect 478506 700176 478512 700188
rect 336700 700148 478512 700176
rect 336700 700136 336706 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 335262 700068 335268 700120
rect 335320 700108 335326 700120
rect 462314 700108 462320 700120
rect 335320 700080 462320 700108
rect 335320 700068 335326 700080
rect 462314 700068 462320 700080
rect 462372 700068 462378 700120
rect 235166 700000 235172 700052
rect 235224 700040 235230 700052
rect 356054 700040 356060 700052
rect 235224 700012 356060 700040
rect 235224 700000 235230 700012
rect 356054 700000 356060 700012
rect 356112 700000 356118 700052
rect 267642 699932 267648 699984
rect 267700 699972 267706 699984
rect 351914 699972 351920 699984
rect 267700 699944 351920 699972
rect 267700 699932 267706 699944
rect 351914 699932 351920 699944
rect 351972 699932 351978 699984
rect 283834 699864 283840 699916
rect 283892 699904 283898 699916
rect 354674 699904 354680 699916
rect 283892 699876 354680 699904
rect 283892 699864 283898 699876
rect 354674 699864 354680 699876
rect 354732 699864 354738 699916
rect 343542 699796 343548 699848
rect 343600 699836 343606 699848
rect 413646 699836 413652 699848
rect 343600 699808 413652 699836
rect 343600 699796 343606 699808
rect 413646 699796 413652 699808
rect 413704 699796 413710 699848
rect 340782 699728 340788 699780
rect 340840 699768 340846 699780
rect 397454 699768 397460 699780
rect 340840 699740 397460 699768
rect 340840 699728 340846 699740
rect 397454 699728 397460 699740
rect 397512 699728 397518 699780
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 332502 699660 332508 699712
rect 332560 699700 332566 699712
rect 346394 699700 346400 699712
rect 332560 699672 346400 699700
rect 332560 699660 332566 699672
rect 346394 699660 346400 699672
rect 346452 699660 346458 699712
rect 347774 699660 347780 699712
rect 347832 699700 347838 699712
rect 348786 699700 348792 699712
rect 347832 699672 348792 699700
rect 347832 699660 347838 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 321462 696940 321468 696992
rect 321520 696980 321526 696992
rect 580166 696980 580172 696992
rect 321520 696952 580172 696980
rect 321520 696940 321526 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 364610 687760 364616 687812
rect 364668 687800 364674 687812
rect 365162 687800 365168 687812
rect 364668 687772 365168 687800
rect 364668 687760 364674 687772
rect 365162 687760 365168 687772
rect 365220 687760 365226 687812
rect 429212 685936 429976 685964
rect 324222 685856 324228 685908
rect 324280 685896 324286 685908
rect 429212 685896 429240 685936
rect 324280 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 324280 685856 324286 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 364521 685831 364579 685837
rect 364521 685797 364533 685831
rect 364567 685828 364579 685831
rect 364610 685828 364616 685840
rect 364567 685800 364616 685828
rect 364567 685797 364579 685800
rect 364521 685791 364579 685797
rect 364610 685788 364616 685800
rect 364668 685788 364674 685840
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 382274 681748 382280 681760
rect 3568 681720 382280 681748
rect 3568 681708 3574 681720
rect 382274 681708 382280 681720
rect 382332 681708 382338 681760
rect 364518 676240 364524 676252
rect 364479 676212 364524 676240
rect 364518 676200 364524 676212
rect 364576 676200 364582 676252
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 320082 673480 320088 673532
rect 320140 673520 320146 673532
rect 580166 673520 580172 673532
rect 320140 673492 580172 673520
rect 320140 673480 320146 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 386414 667944 386420 667956
rect 3476 667916 386420 667944
rect 3476 667904 3482 667916
rect 386414 667904 386420 667916
rect 386472 667904 386478 667956
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 383654 652780 383660 652792
rect 3108 652752 383660 652780
rect 3108 652740 3114 652752
rect 383654 652740 383660 652752
rect 383712 652740 383718 652792
rect 315942 650020 315948 650072
rect 316000 650060 316006 650072
rect 580166 650060 580172 650072
rect 316000 650032 580172 650060
rect 316000 650020 316006 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 317322 638936 317328 638988
rect 317380 638976 317386 638988
rect 580166 638976 580172 638988
rect 317380 638948 580172 638976
rect 317380 638936 317386 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 313182 626560 313188 626612
rect 313240 626600 313246 626612
rect 580166 626600 580172 626612
rect 313240 626572 580172 626600
rect 313240 626560 313246 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 387794 623812 387800 623824
rect 3476 623784 387800 623812
rect 3476 623772 3482 623784
rect 387794 623772 387800 623784
rect 387852 623772 387858 623824
rect 364521 618239 364579 618245
rect 364521 618205 364533 618239
rect 364567 618236 364579 618239
rect 364610 618236 364616 618248
rect 364567 618208 364616 618236
rect 364567 618205 364579 618208
rect 364521 618199 364579 618205
rect 364610 618196 364616 618208
rect 364668 618196 364674 618248
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 391934 610008 391940 610020
rect 3476 609980 391940 610008
rect 3476 609968 3482 609980
rect 391934 609968 391940 609980
rect 391992 609968 391998 610020
rect 364518 608648 364524 608660
rect 364479 608620 364524 608648
rect 364518 608608 364524 608620
rect 364576 608608 364582 608660
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 309042 603100 309048 603152
rect 309100 603140 309106 603152
rect 580166 603140 580172 603152
rect 309100 603112 580172 603140
rect 309100 603100 309106 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 364610 598924 364616 598936
rect 364571 598896 364616 598924
rect 364610 598884 364616 598896
rect 364668 598884 364674 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 390554 594844 390560 594856
rect 3292 594816 390560 594844
rect 3292 594804 3298 594816
rect 390554 594804 390560 594816
rect 390612 594804 390618 594856
rect 311802 592016 311808 592068
rect 311860 592056 311866 592068
rect 580166 592056 580172 592068
rect 311860 592028 580172 592056
rect 311860 592016 311866 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 364613 589339 364671 589345
rect 364613 589305 364625 589339
rect 364659 589336 364671 589339
rect 364702 589336 364708 589348
rect 364659 589308 364708 589336
rect 364659 589305 364671 589308
rect 364613 589299 364671 589305
rect 364702 589296 364708 589308
rect 364760 589296 364766 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 344462 584672 344468 584724
rect 344520 584712 344526 584724
rect 364702 584712 364708 584724
rect 344520 584684 364708 584712
rect 344520 584672 344526 584684
rect 364702 584672 364708 584684
rect 364760 584672 364766 584724
rect 300762 584604 300768 584656
rect 300820 584644 300826 584656
rect 350810 584644 350816 584656
rect 300820 584616 350816 584644
rect 300820 584604 300826 584616
rect 350810 584604 350816 584616
rect 350868 584604 350874 584656
rect 338206 584536 338212 584588
rect 338264 584576 338270 584588
rect 429654 584576 429660 584588
rect 338264 584548 429660 584576
rect 338264 584536 338270 584548
rect 429654 584536 429660 584548
rect 429712 584536 429718 584588
rect 331858 584468 331864 584520
rect 331916 584508 331922 584520
rect 494238 584508 494244 584520
rect 331916 584480 494244 584508
rect 331916 584468 331922 584480
rect 494238 584468 494244 584480
rect 494296 584468 494302 584520
rect 325510 584400 325516 584452
rect 325568 584440 325574 584452
rect 559374 584440 559380 584452
rect 325568 584412 559380 584440
rect 325568 584400 325574 584412
rect 559374 584400 559380 584412
rect 559432 584400 559438 584452
rect 304534 583652 304540 583704
rect 304592 583692 304598 583704
rect 471330 583692 471336 583704
rect 304592 583664 471336 583692
rect 304592 583652 304598 583664
rect 471330 583652 471336 583664
rect 471388 583652 471394 583704
rect 298186 583584 298192 583636
rect 298244 583624 298250 583636
rect 471238 583624 471244 583636
rect 298244 583596 471244 583624
rect 298244 583584 298250 583596
rect 471238 583584 471244 583596
rect 471296 583584 471302 583636
rect 256050 583516 256056 583568
rect 256108 583556 256114 583568
rect 580626 583556 580632 583568
rect 256108 583528 580632 583556
rect 256108 583516 256114 583528
rect 580626 583516 580632 583528
rect 580684 583516 580690 583568
rect 251818 583448 251824 583500
rect 251876 583488 251882 583500
rect 580534 583488 580540 583500
rect 251876 583460 580540 583488
rect 251876 583448 251882 583460
rect 580534 583448 580540 583460
rect 580592 583448 580598 583500
rect 245562 583380 245568 583432
rect 245620 583420 245626 583432
rect 580350 583420 580356 583432
rect 245620 583392 580356 583420
rect 245620 583380 245626 583392
rect 580350 583380 580356 583392
rect 580408 583380 580414 583432
rect 4706 583312 4712 583364
rect 4764 583352 4770 583364
rect 399202 583352 399208 583364
rect 4764 583324 399208 583352
rect 4764 583312 4770 583324
rect 399202 583312 399208 583324
rect 399260 583312 399266 583364
rect 5442 583244 5448 583296
rect 5500 583284 5506 583296
rect 405550 583284 405556 583296
rect 5500 583256 405556 583284
rect 5500 583244 5506 583256
rect 405550 583244 405556 583256
rect 405608 583244 405614 583296
rect 10318 583176 10324 583228
rect 10376 583216 10382 583228
rect 411898 583216 411904 583228
rect 10376 583188 411904 583216
rect 10376 583176 10382 583188
rect 411898 583176 411904 583188
rect 411956 583176 411962 583228
rect 6270 583108 6276 583160
rect 6328 583148 6334 583160
rect 409782 583148 409788 583160
rect 6328 583120 409788 583148
rect 6328 583108 6334 583120
rect 409782 583108 409788 583120
rect 409840 583108 409846 583160
rect 3142 583040 3148 583092
rect 3200 583080 3206 583092
rect 407666 583080 407672 583092
rect 3200 583052 407672 583080
rect 3200 583040 3206 583052
rect 407666 583040 407672 583052
rect 407724 583040 407730 583092
rect 13078 582972 13084 583024
rect 13136 583012 13142 583024
rect 418154 583012 418160 583024
rect 13136 582984 418160 583012
rect 13136 582972 13142 582984
rect 418154 582972 418160 582984
rect 418212 582972 418218 583024
rect 14458 582904 14464 582956
rect 14516 582944 14522 582956
rect 424502 582944 424508 582956
rect 14516 582916 424508 582944
rect 14516 582904 14522 582916
rect 424502 582904 424508 582916
rect 424560 582904 424566 582956
rect 3234 582836 3240 582888
rect 3292 582876 3298 582888
rect 414014 582876 414020 582888
rect 3292 582848 414020 582876
rect 3292 582836 3298 582848
rect 414014 582836 414020 582848
rect 414072 582836 414078 582888
rect 5350 582768 5356 582820
rect 5408 582808 5414 582820
rect 422386 582808 422392 582820
rect 5408 582780 422392 582808
rect 5408 582768 5414 582780
rect 422386 582768 422392 582780
rect 422444 582768 422450 582820
rect 15838 582700 15844 582752
rect 15896 582740 15902 582752
rect 437106 582740 437112 582752
rect 15896 582712 437112 582740
rect 15896 582700 15902 582712
rect 437106 582700 437112 582712
rect 437164 582700 437170 582752
rect 4062 582632 4068 582684
rect 4120 582672 4126 582684
rect 430850 582672 430856 582684
rect 4120 582644 430856 582672
rect 4120 582632 4126 582644
rect 430850 582632 430856 582644
rect 430908 582632 430914 582684
rect 5258 582564 5264 582616
rect 5316 582604 5322 582616
rect 432966 582604 432972 582616
rect 5316 582576 432972 582604
rect 5316 582564 5322 582576
rect 432966 582564 432972 582576
rect 433024 582564 433030 582616
rect 3878 582496 3884 582548
rect 3936 582536 3942 582548
rect 434990 582536 434996 582548
rect 3936 582508 434996 582536
rect 3936 582496 3942 582508
rect 434990 582496 434996 582508
rect 435048 582496 435054 582548
rect 5166 582428 5172 582480
rect 5224 582468 5230 582480
rect 445570 582468 445576 582480
rect 5224 582440 445576 582468
rect 5224 582428 5230 582440
rect 445570 582428 445576 582440
rect 445628 582428 445634 582480
rect 3694 582360 3700 582412
rect 3752 582400 3758 582412
rect 443454 582400 443460 582412
rect 3752 582372 443460 582400
rect 3752 582360 3758 582372
rect 443454 582360 443460 582372
rect 443512 582360 443518 582412
rect 302418 581476 302424 581528
rect 302476 581516 302482 581528
rect 469582 581516 469588 581528
rect 302476 581488 469588 581516
rect 302476 581476 302482 581488
rect 469582 581476 469588 581488
rect 469640 581476 469646 581528
rect 296070 581408 296076 581460
rect 296128 581448 296134 581460
rect 469674 581448 469680 581460
rect 296128 581420 469680 581448
rect 296128 581408 296134 581420
rect 469674 581408 469680 581420
rect 469732 581408 469738 581460
rect 289722 581340 289728 581392
rect 289780 581380 289786 581392
rect 469766 581380 469772 581392
rect 289780 581352 469772 581380
rect 289780 581340 289786 581352
rect 469766 581340 469772 581352
rect 469824 581340 469830 581392
rect 287606 581272 287612 581324
rect 287664 581312 287670 581324
rect 470502 581312 470508 581324
rect 287664 581284 470508 581312
rect 287664 581272 287670 581284
rect 470502 581272 470508 581284
rect 470560 581272 470566 581324
rect 283466 581204 283472 581256
rect 283524 581244 283530 581256
rect 470410 581244 470416 581256
rect 283524 581216 470416 581244
rect 283524 581204 283530 581216
rect 470410 581204 470416 581216
rect 470468 581204 470474 581256
rect 281350 581136 281356 581188
rect 281408 581176 281414 581188
rect 470226 581176 470232 581188
rect 281408 581148 470232 581176
rect 281408 581136 281414 581148
rect 470226 581136 470232 581148
rect 470284 581136 470290 581188
rect 275002 581068 275008 581120
rect 275060 581108 275066 581120
rect 470134 581108 470140 581120
rect 275060 581080 470140 581108
rect 275060 581068 275066 581080
rect 470134 581068 470140 581080
rect 470192 581068 470198 581120
rect 264514 581000 264520 581052
rect 264572 581040 264578 581052
rect 580074 581040 580080 581052
rect 264572 581012 580080 581040
rect 264572 581000 264578 581012
rect 580074 581000 580080 581012
rect 580132 581000 580138 581052
rect 268654 580320 268660 580372
rect 268712 580360 268718 580372
rect 469950 580360 469956 580372
rect 268712 580332 469956 580360
rect 268712 580320 268718 580332
rect 469950 580320 469956 580332
rect 470008 580320 470014 580372
rect 262398 580252 262404 580304
rect 262456 580292 262462 580304
rect 469858 580292 469864 580304
rect 262456 580264 469864 580292
rect 262456 580252 262462 580264
rect 469858 580252 469864 580264
rect 469916 580252 469922 580304
rect 306558 580184 306564 580236
rect 306616 580224 306622 580236
rect 580166 580224 580172 580236
rect 306616 580196 580172 580224
rect 306616 580184 306622 580196
rect 580166 580184 580172 580196
rect 580224 580184 580230 580236
rect 6638 580116 6644 580168
rect 6696 580156 6702 580168
rect 395062 580156 395068 580168
rect 6696 580128 395068 580156
rect 6696 580116 6702 580128
rect 395062 580116 395068 580128
rect 395120 580116 395126 580168
rect 6546 580048 6552 580100
rect 6604 580088 6610 580100
rect 397086 580088 397092 580100
rect 6604 580060 397092 580088
rect 6604 580048 6610 580060
rect 397086 580048 397092 580060
rect 397144 580048 397150 580100
rect 6454 579980 6460 580032
rect 6512 580020 6518 580032
rect 400950 580020 400956 580032
rect 6512 579992 400956 580020
rect 6512 579980 6518 579992
rect 400950 579980 400956 579992
rect 401008 579980 401014 580032
rect 6362 579912 6368 579964
rect 6420 579952 6426 579964
rect 403158 579952 403164 579964
rect 6420 579924 403164 579952
rect 6420 579912 6426 579924
rect 403158 579912 403164 579924
rect 403216 579912 403222 579964
rect 3786 579844 3792 579896
rect 3844 579884 3850 579896
rect 438854 579884 438860 579896
rect 3844 579856 438860 579884
rect 3844 579844 3850 579856
rect 438854 579844 438860 579856
rect 438912 579844 438918 579896
rect 4982 579776 4988 579828
rect 5040 579816 5046 579828
rect 451550 579816 451556 579828
rect 5040 579788 451556 579816
rect 5040 579776 5046 579788
rect 451550 579776 451556 579788
rect 451608 579776 451614 579828
rect 4890 579708 4896 579760
rect 4948 579748 4954 579760
rect 458266 579748 458272 579760
rect 4948 579720 458272 579748
rect 4948 579708 4954 579720
rect 458266 579708 458272 579720
rect 458324 579708 458330 579760
rect 6178 579640 6184 579692
rect 6236 579680 6242 579692
rect 464246 579680 464252 579692
rect 6236 579652 464252 579680
rect 6236 579640 6242 579652
rect 464246 579640 464252 579652
rect 464304 579640 464310 579692
rect 271138 579368 271144 579420
rect 271196 579408 271202 579420
rect 271196 579380 282224 579408
rect 271196 579368 271202 579380
rect 247954 579340 247960 579352
rect 247915 579312 247960 579340
rect 247954 579300 247960 579312
rect 248012 579300 248018 579352
rect 254210 579340 254216 579352
rect 254171 579312 254216 579340
rect 254210 579300 254216 579312
rect 254268 579300 254274 579352
rect 258442 579300 258448 579352
rect 258500 579300 258506 579352
rect 260650 579300 260656 579352
rect 260708 579300 260714 579352
rect 266906 579300 266912 579352
rect 266964 579300 266970 579352
rect 273162 579300 273168 579352
rect 273220 579300 273226 579352
rect 277302 579300 277308 579352
rect 277360 579300 277366 579352
rect 279602 579300 279608 579352
rect 279660 579300 279666 579352
rect 258460 578728 258488 579300
rect 260668 578796 260696 579300
rect 266924 578864 266952 579300
rect 273180 578932 273208 579300
rect 277320 579000 277348 579300
rect 279620 579068 279648 579300
rect 282196 579204 282224 579380
rect 285766 579300 285772 579352
rect 285824 579300 285830 579352
rect 292114 579340 292120 579352
rect 292075 579312 292120 579340
rect 292114 579300 292120 579312
rect 292172 579300 292178 579352
rect 415670 579340 415676 579352
rect 415631 579312 415676 579340
rect 415670 579300 415676 579312
rect 415728 579300 415734 579352
rect 428366 579340 428372 579352
rect 428327 579312 428372 579340
rect 428366 579300 428372 579312
rect 428424 579300 428430 579352
rect 441062 579340 441068 579352
rect 441023 579312 441068 579340
rect 441062 579300 441068 579312
rect 441120 579300 441126 579352
rect 453574 579340 453580 579352
rect 453535 579312 453580 579340
rect 453574 579300 453580 579312
rect 453632 579300 453638 579352
rect 455782 579340 455788 579352
rect 455743 579312 455788 579340
rect 455782 579300 455788 579312
rect 455840 579300 455846 579352
rect 285784 579272 285812 579300
rect 470318 579272 470324 579284
rect 285784 579244 470324 579272
rect 470318 579232 470324 579244
rect 470376 579232 470382 579284
rect 470042 579204 470048 579216
rect 282196 579176 470048 579204
rect 470042 579164 470048 579176
rect 470100 579164 470106 579216
rect 292117 579139 292175 579145
rect 292117 579105 292129 579139
rect 292163 579136 292175 579139
rect 579798 579136 579804 579148
rect 292163 579108 579804 579136
rect 292163 579105 292175 579108
rect 292117 579099 292175 579105
rect 579798 579096 579804 579108
rect 579856 579096 579862 579148
rect 579982 579068 579988 579080
rect 279620 579040 579988 579068
rect 579982 579028 579988 579040
rect 580040 579028 580046 579080
rect 579890 579000 579896 579012
rect 277320 578972 579896 579000
rect 579890 578960 579896 578972
rect 579948 578960 579954 579012
rect 580074 578932 580080 578944
rect 273180 578904 580080 578932
rect 580074 578892 580080 578904
rect 580132 578892 580138 578944
rect 580902 578864 580908 578876
rect 266924 578836 580908 578864
rect 580902 578824 580908 578836
rect 580960 578824 580966 578876
rect 580718 578796 580724 578808
rect 260668 578768 580724 578796
rect 580718 578756 580724 578768
rect 580776 578756 580782 578808
rect 580810 578728 580816 578740
rect 258460 578700 580816 578728
rect 580810 578688 580816 578700
rect 580868 578688 580874 578740
rect 254213 578663 254271 578669
rect 254213 578629 254225 578663
rect 254259 578660 254271 578663
rect 580442 578660 580448 578672
rect 254259 578632 580448 578660
rect 254259 578629 254271 578632
rect 254213 578623 254271 578629
rect 580442 578620 580448 578632
rect 580500 578620 580506 578672
rect 247957 578595 248015 578601
rect 247957 578561 247969 578595
rect 248003 578592 248015 578595
rect 580258 578592 580264 578604
rect 248003 578564 580264 578592
rect 248003 578561 248015 578564
rect 247957 578555 248015 578561
rect 580258 578552 580264 578564
rect 580316 578552 580322 578604
rect 3326 578484 3332 578536
rect 3384 578524 3390 578536
rect 415673 578527 415731 578533
rect 415673 578524 415685 578527
rect 3384 578496 415685 578524
rect 3384 578484 3390 578496
rect 415673 578493 415685 578496
rect 415719 578493 415731 578527
rect 415673 578487 415731 578493
rect 3970 578416 3976 578468
rect 4028 578456 4034 578468
rect 428369 578459 428427 578465
rect 428369 578456 428381 578459
rect 4028 578428 428381 578456
rect 4028 578416 4034 578428
rect 428369 578425 428381 578428
rect 428415 578425 428427 578459
rect 428369 578419 428427 578425
rect 3602 578348 3608 578400
rect 3660 578388 3666 578400
rect 441065 578391 441123 578397
rect 441065 578388 441077 578391
rect 3660 578360 441077 578388
rect 3660 578348 3666 578360
rect 441065 578357 441077 578360
rect 441111 578357 441123 578391
rect 441065 578351 441123 578357
rect 3418 578280 3424 578332
rect 3476 578320 3482 578332
rect 453577 578323 453635 578329
rect 453577 578320 453589 578323
rect 3476 578292 453589 578320
rect 3476 578280 3482 578292
rect 453577 578289 453589 578292
rect 453623 578289 453635 578323
rect 453577 578283 453635 578289
rect 3510 578212 3516 578264
rect 3568 578252 3574 578264
rect 455785 578255 455843 578261
rect 455785 578252 455797 578255
rect 3568 578224 455797 578252
rect 3568 578212 3574 578224
rect 455785 578221 455797 578224
rect 455831 578221 455843 578255
rect 455785 578215 455843 578221
rect 3050 567332 3056 567384
rect 3108 567372 3114 567384
rect 6638 567372 6644 567384
rect 3108 567344 6644 567372
rect 3108 567332 3114 567344
rect 6638 567332 6644 567344
rect 6696 567332 6702 567384
rect 469582 557472 469588 557524
rect 469640 557512 469646 557524
rect 579706 557512 579712 557524
rect 469640 557484 579712 557512
rect 469640 557472 469646 557484
rect 579706 557472 579712 557484
rect 579764 557472 579770 557524
rect 2774 553052 2780 553104
rect 2832 553092 2838 553104
rect 4706 553092 4712 553104
rect 2832 553064 4712 553092
rect 2832 553052 2838 553064
rect 4706 553052 4712 553064
rect 4764 553052 4770 553104
rect 471330 546388 471336 546440
rect 471388 546428 471394 546440
rect 579706 546428 579712 546440
rect 471388 546400 579712 546428
rect 471388 546388 471394 546400
rect 579706 546388 579712 546400
rect 579764 546388 579770 546440
rect 3050 538636 3056 538688
rect 3108 538676 3114 538688
rect 6546 538676 6552 538688
rect 3108 538648 6552 538676
rect 3108 538636 3114 538648
rect 6546 538636 6552 538648
rect 6604 538636 6610 538688
rect 469674 510552 469680 510604
rect 469732 510592 469738 510604
rect 579706 510592 579712 510604
rect 469732 510564 579712 510592
rect 469732 510552 469738 510564
rect 579706 510552 579712 510564
rect 579764 510552 579770 510604
rect 3050 510212 3056 510264
rect 3108 510252 3114 510264
rect 6454 510252 6460 510264
rect 3108 510224 6460 510252
rect 3108 510212 3114 510224
rect 6454 510212 6460 510224
rect 6512 510212 6518 510264
rect 471238 499468 471244 499520
rect 471296 499508 471302 499520
rect 579706 499508 579712 499520
rect 471296 499480 579712 499508
rect 471296 499468 471302 499480
rect 579706 499468 579712 499480
rect 579764 499468 579770 499520
rect 2774 496680 2780 496732
rect 2832 496720 2838 496732
rect 5442 496720 5448 496732
rect 2832 496692 5448 496720
rect 2832 496680 2838 496692
rect 5442 496680 5448 496692
rect 5500 496680 5506 496732
rect 2958 481108 2964 481160
rect 3016 481148 3022 481160
rect 6362 481148 6368 481160
rect 3016 481120 6368 481148
rect 3016 481108 3022 481120
rect 6362 481108 6368 481120
rect 6420 481108 6426 481160
rect 469766 463632 469772 463684
rect 469824 463672 469830 463684
rect 579706 463672 579712 463684
rect 469824 463644 579712 463672
rect 469824 463632 469830 463644
rect 579706 463632 579712 463644
rect 579764 463632 579770 463684
rect 470502 440172 470508 440224
rect 470560 440212 470566 440224
rect 579798 440212 579804 440224
rect 470560 440184 579804 440212
rect 470560 440172 470566 440184
rect 579798 440172 579804 440184
rect 579856 440172 579862 440224
rect 3142 438812 3148 438864
rect 3200 438852 3206 438864
rect 10318 438852 10324 438864
rect 3200 438824 10324 438852
rect 3200 438812 3206 438824
rect 10318 438812 10324 438824
rect 10376 438812 10382 438864
rect 3142 424056 3148 424108
rect 3200 424096 3206 424108
rect 6270 424096 6276 424108
rect 3200 424068 6276 424096
rect 3200 424056 3206 424068
rect 6270 424056 6276 424068
rect 6328 424056 6334 424108
rect 470410 416712 470416 416764
rect 470468 416752 470474 416764
rect 579798 416752 579804 416764
rect 470468 416724 579804 416752
rect 470468 416712 470474 416724
rect 579798 416712 579804 416724
rect 579856 416712 579862 416764
rect 470318 405628 470324 405680
rect 470376 405668 470382 405680
rect 579798 405668 579804 405680
rect 470376 405640 579804 405668
rect 470376 405628 470382 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 470226 393252 470232 393304
rect 470284 393292 470290 393304
rect 579798 393292 579804 393304
rect 470284 393264 579804 393292
rect 470284 393252 470290 393264
rect 579798 393252 579804 393264
rect 579856 393252 579862 393304
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 13078 380848 13084 380860
rect 3292 380820 13084 380848
rect 3292 380808 3298 380820
rect 13078 380808 13084 380820
rect 13136 380808 13142 380860
rect 470134 346332 470140 346384
rect 470192 346372 470198 346384
rect 579982 346372 579988 346384
rect 470192 346344 579988 346372
rect 470192 346332 470198 346344
rect 579982 346332 579988 346344
rect 580040 346332 580046 346384
rect 238757 338691 238815 338697
rect 238757 338657 238769 338691
rect 238803 338688 238815 338691
rect 244642 338688 244648 338700
rect 238803 338660 244648 338688
rect 238803 338657 238815 338660
rect 238757 338651 238815 338657
rect 244642 338648 244648 338660
rect 244700 338648 244706 338700
rect 346397 338691 346455 338697
rect 346397 338657 346409 338691
rect 346443 338688 346455 338691
rect 348510 338688 348516 338700
rect 346443 338660 348516 338688
rect 346443 338657 346455 338660
rect 346397 338651 346455 338657
rect 348510 338648 348516 338660
rect 348568 338648 348574 338700
rect 229097 338147 229155 338153
rect 229097 338113 229109 338147
rect 229143 338144 229155 338147
rect 238665 338147 238723 338153
rect 238665 338144 238677 338147
rect 229143 338116 238677 338144
rect 229143 338113 229155 338116
rect 229097 338107 229155 338113
rect 238665 338113 238677 338116
rect 238711 338113 238723 338147
rect 238665 338107 238723 338113
rect 316126 338104 316132 338156
rect 316184 338144 316190 338156
rect 316310 338144 316316 338156
rect 316184 338116 316316 338144
rect 316184 338104 316190 338116
rect 316310 338104 316316 338116
rect 316368 338104 316374 338156
rect 318794 338104 318800 338156
rect 318852 338144 318858 338156
rect 319806 338144 319812 338156
rect 318852 338116 319812 338144
rect 318852 338104 318858 338116
rect 319806 338104 319812 338116
rect 319864 338104 319870 338156
rect 327077 338147 327135 338153
rect 327077 338113 327089 338147
rect 327123 338144 327135 338147
rect 336645 338147 336703 338153
rect 336645 338144 336657 338147
rect 327123 338116 336657 338144
rect 327123 338113 327135 338116
rect 327077 338107 327135 338113
rect 336645 338113 336657 338116
rect 336691 338113 336703 338147
rect 336645 338107 336703 338113
rect 337378 338104 337384 338156
rect 337436 338144 337442 338156
rect 337746 338144 337752 338156
rect 337436 338116 337752 338144
rect 337436 338104 337442 338116
rect 337746 338104 337752 338116
rect 337804 338104 337810 338156
rect 340322 338104 340328 338156
rect 340380 338144 340386 338156
rect 340690 338144 340696 338156
rect 340380 338116 340696 338144
rect 340380 338104 340386 338116
rect 340690 338104 340696 338116
rect 340748 338104 340754 338156
rect 365165 338147 365223 338153
rect 365165 338113 365177 338147
rect 365211 338144 365223 338147
rect 372062 338144 372068 338156
rect 365211 338116 372068 338144
rect 365211 338113 365223 338116
rect 365165 338107 365223 338113
rect 372062 338104 372068 338116
rect 372120 338104 372126 338156
rect 460842 338104 460848 338156
rect 460900 338144 460906 338156
rect 466365 338147 466423 338153
rect 466365 338144 466377 338147
rect 460900 338116 466377 338144
rect 460900 338104 460906 338116
rect 466365 338113 466377 338116
rect 466411 338113 466423 338147
rect 466365 338107 466423 338113
rect 71038 338036 71044 338088
rect 71096 338076 71102 338088
rect 86957 338079 87015 338085
rect 86957 338076 86969 338079
rect 71096 338048 86969 338076
rect 71096 338036 71102 338048
rect 86957 338045 86969 338048
rect 87003 338045 87015 338079
rect 86957 338039 87015 338045
rect 87233 338079 87291 338085
rect 87233 338045 87245 338079
rect 87279 338076 87291 338079
rect 254946 338076 254952 338088
rect 87279 338048 254952 338076
rect 87279 338045 87291 338048
rect 87233 338039 87291 338045
rect 254946 338036 254952 338048
rect 255004 338036 255010 338088
rect 314654 338036 314660 338088
rect 314712 338076 314718 338088
rect 315390 338076 315396 338088
rect 314712 338048 315396 338076
rect 314712 338036 314718 338048
rect 315390 338036 315396 338048
rect 315448 338036 315454 338088
rect 315485 338079 315543 338085
rect 315485 338045 315497 338079
rect 315531 338076 315543 338079
rect 318889 338079 318947 338085
rect 318889 338076 318901 338079
rect 315531 338048 318901 338076
rect 315531 338045 315543 338048
rect 315485 338039 315543 338045
rect 318889 338045 318901 338048
rect 318935 338045 318947 338079
rect 318889 338039 318947 338045
rect 319073 338079 319131 338085
rect 319073 338045 319085 338079
rect 319119 338076 319131 338079
rect 354398 338076 354404 338088
rect 319119 338048 354404 338076
rect 319119 338045 319131 338048
rect 319073 338039 319131 338045
rect 354398 338036 354404 338048
rect 354456 338036 354462 338088
rect 358078 338036 358084 338088
rect 358136 338076 358142 338088
rect 371510 338076 371516 338088
rect 358136 338048 371516 338076
rect 358136 338036 358142 338048
rect 371510 338036 371516 338048
rect 371568 338036 371574 338088
rect 374641 338079 374699 338085
rect 374641 338045 374653 338079
rect 374687 338076 374699 338079
rect 376757 338079 376815 338085
rect 376757 338076 376769 338079
rect 374687 338048 376769 338076
rect 374687 338045 374699 338048
rect 374641 338039 374699 338045
rect 376757 338045 376769 338048
rect 376803 338045 376815 338079
rect 376757 338039 376815 338045
rect 406286 338036 406292 338088
rect 406344 338076 406350 338088
rect 417418 338076 417424 338088
rect 406344 338048 417424 338076
rect 406344 338036 406350 338048
rect 417418 338036 417424 338048
rect 417476 338036 417482 338088
rect 419074 338036 419080 338088
rect 419132 338076 419138 338088
rect 431402 338076 431408 338088
rect 419132 338048 431408 338076
rect 419132 338036 419138 338048
rect 431402 338036 431408 338048
rect 431460 338036 431466 338088
rect 435726 338036 435732 338088
rect 435784 338076 435790 338088
rect 499574 338076 499580 338088
rect 435784 338048 499580 338076
rect 435784 338036 435790 338048
rect 499574 338036 499580 338048
rect 499632 338036 499638 338088
rect 66898 337968 66904 338020
rect 66956 338008 66962 338020
rect 252002 338008 252008 338020
rect 66956 337980 252008 338008
rect 66956 337968 66962 337980
rect 252002 337968 252008 337980
rect 252060 337968 252066 338020
rect 306190 337968 306196 338020
rect 306248 338008 306254 338020
rect 355870 338008 355876 338020
rect 306248 337980 355876 338008
rect 306248 337968 306254 337980
rect 355870 337968 355876 337980
rect 355928 337968 355934 338020
rect 364242 337968 364248 338020
rect 364300 338008 364306 338020
rect 379330 338008 379336 338020
rect 364300 337980 379336 338008
rect 364300 337968 364306 337980
rect 379330 337968 379336 337980
rect 379388 337968 379394 338020
rect 382274 338008 382280 338020
rect 379440 337980 382280 338008
rect 61378 337900 61384 337952
rect 61436 337940 61442 337952
rect 87049 337943 87107 337949
rect 87049 337940 87061 337943
rect 61436 337912 87061 337940
rect 61436 337900 61442 337912
rect 87049 337909 87061 337912
rect 87095 337909 87107 337943
rect 87049 337903 87107 337909
rect 87233 337943 87291 337949
rect 87233 337909 87245 337943
rect 87279 337940 87291 337943
rect 247586 337940 247592 337952
rect 87279 337912 247592 337940
rect 87279 337909 87291 337912
rect 87233 337903 87291 337909
rect 247586 337900 247592 337912
rect 247644 337900 247650 337952
rect 303154 337900 303160 337952
rect 303212 337940 303218 337952
rect 318889 337943 318947 337949
rect 318889 337940 318901 337943
rect 303212 337912 318901 337940
rect 303212 337900 303218 337912
rect 318889 337909 318901 337912
rect 318935 337909 318947 337943
rect 318889 337903 318947 337909
rect 318981 337943 319039 337949
rect 318981 337909 318993 337943
rect 319027 337940 319039 337943
rect 352926 337940 352932 337952
rect 319027 337912 352932 337940
rect 319027 337909 319039 337912
rect 318981 337903 319039 337909
rect 352926 337900 352932 337912
rect 352984 337900 352990 337952
rect 355318 337900 355324 337952
rect 355376 337940 355382 337952
rect 370038 337940 370044 337952
rect 355376 337912 370044 337940
rect 355376 337900 355382 337912
rect 370038 337900 370044 337912
rect 370096 337900 370102 337952
rect 371142 337900 371148 337952
rect 371200 337940 371206 337952
rect 379440 337940 379468 337980
rect 382274 337968 382280 337980
rect 382332 337968 382338 338020
rect 397454 337968 397460 338020
rect 397512 338008 397518 338020
rect 403618 338008 403624 338020
rect 397512 337980 403624 338008
rect 397512 337968 397518 337980
rect 403618 337968 403624 337980
rect 403676 337968 403682 338020
rect 414658 337968 414664 338020
rect 414716 338008 414722 338020
rect 429746 338008 429752 338020
rect 414716 337980 429752 338008
rect 414716 337968 414722 337980
rect 429746 337968 429752 337980
rect 429804 337968 429810 338020
rect 437198 337968 437204 338020
rect 437256 338008 437262 338020
rect 442350 338008 442356 338020
rect 437256 337980 442356 338008
rect 437256 337968 437262 337980
rect 442350 337968 442356 337980
rect 442408 337968 442414 338020
rect 446030 337968 446036 338020
rect 446088 338008 446094 338020
rect 451461 338011 451519 338017
rect 451461 338008 451473 338011
rect 446088 337980 451473 338008
rect 446088 337968 446094 337980
rect 451461 337977 451473 337980
rect 451507 337977 451519 338011
rect 451461 337971 451519 337977
rect 454770 337968 454776 338020
rect 454828 338008 454834 338020
rect 461581 338011 461639 338017
rect 461581 338008 461593 338011
rect 454828 337980 461593 338008
rect 454828 337968 454834 337980
rect 461581 337977 461593 337980
rect 461627 337977 461639 338011
rect 461581 337971 461639 337977
rect 461670 337968 461676 338020
rect 461728 338008 461734 338020
rect 466273 338011 466331 338017
rect 466273 338008 466285 338011
rect 461728 337980 466285 338008
rect 461728 337968 461734 337980
rect 466273 337977 466285 337980
rect 466319 337977 466331 338011
rect 466273 337971 466331 337977
rect 466365 338011 466423 338017
rect 466365 337977 466377 338011
rect 466411 338008 466423 338011
rect 525058 338008 525064 338020
rect 466411 337980 525064 338008
rect 466411 337977 466423 337980
rect 466365 337971 466423 337977
rect 525058 337968 525064 337980
rect 525116 337968 525122 338020
rect 371200 337912 379468 337940
rect 371200 337900 371206 337912
rect 400398 337900 400404 337952
rect 400456 337940 400462 337952
rect 413278 337940 413284 337952
rect 400456 337912 413284 337940
rect 400456 337900 400462 337912
rect 413278 337900 413284 337912
rect 413336 337900 413342 337952
rect 413646 337900 413652 337952
rect 413704 337940 413710 337952
rect 420178 337940 420184 337952
rect 413704 337912 420184 337940
rect 413704 337900 413710 337912
rect 420178 337900 420184 337912
rect 420236 337900 420242 337952
rect 420546 337900 420552 337952
rect 420604 337940 420610 337952
rect 441617 337943 441675 337949
rect 441617 337940 441629 337943
rect 420604 337912 441629 337940
rect 420604 337900 420610 337912
rect 441617 337909 441629 337912
rect 441663 337909 441675 337943
rect 441617 337903 441675 337909
rect 451093 337943 451151 337949
rect 451093 337909 451105 337943
rect 451139 337940 451151 337943
rect 451277 337943 451335 337949
rect 451277 337940 451289 337943
rect 451139 337912 451289 337940
rect 451139 337909 451151 337912
rect 451093 337903 451151 337909
rect 451277 337909 451289 337912
rect 451323 337909 451335 337943
rect 455598 337940 455604 337952
rect 451277 337903 451335 337909
rect 451384 337912 455604 337940
rect 57238 337832 57244 337884
rect 57296 337872 57302 337884
rect 247126 337872 247132 337884
rect 57296 337844 247132 337872
rect 57296 337832 57302 337844
rect 247126 337832 247132 337844
rect 247184 337832 247190 337884
rect 290458 337832 290464 337884
rect 290516 337872 290522 337884
rect 335909 337875 335967 337881
rect 335909 337872 335921 337875
rect 290516 337844 335921 337872
rect 290516 337832 290522 337844
rect 335909 337841 335921 337844
rect 335955 337841 335967 337875
rect 335909 337835 335967 337841
rect 336001 337875 336059 337881
rect 336001 337841 336013 337875
rect 336047 337872 336059 337875
rect 347038 337872 347044 337884
rect 336047 337844 347044 337872
rect 336047 337841 336059 337844
rect 336001 337835 336059 337841
rect 347038 337832 347044 337844
rect 347096 337832 347102 337884
rect 348418 337832 348424 337884
rect 348476 337872 348482 337884
rect 365622 337872 365628 337884
rect 348476 337844 365628 337872
rect 348476 337832 348482 337844
rect 365622 337832 365628 337844
rect 365680 337832 365686 337884
rect 378870 337872 378876 337884
rect 370332 337844 378876 337872
rect 50338 337764 50344 337816
rect 50396 337804 50402 337816
rect 87049 337807 87107 337813
rect 87049 337804 87061 337807
rect 50396 337776 87061 337804
rect 50396 337764 50402 337776
rect 87049 337773 87061 337776
rect 87095 337773 87107 337807
rect 87049 337767 87107 337773
rect 87233 337807 87291 337813
rect 87233 337773 87245 337807
rect 87279 337804 87291 337807
rect 244182 337804 244188 337816
rect 87279 337776 244188 337804
rect 87279 337773 87291 337776
rect 87233 337767 87291 337773
rect 244182 337764 244188 337776
rect 244240 337764 244246 337816
rect 259638 337764 259644 337816
rect 259696 337804 259702 337816
rect 260098 337804 260104 337816
rect 259696 337776 260104 337804
rect 259696 337764 259702 337776
rect 260098 337764 260104 337776
rect 260156 337764 260162 337816
rect 288250 337764 288256 337816
rect 288308 337804 288314 337816
rect 302145 337807 302203 337813
rect 302145 337804 302157 337807
rect 288308 337776 302157 337804
rect 288308 337764 288314 337776
rect 302145 337773 302157 337776
rect 302191 337773 302203 337807
rect 302145 337767 302203 337773
rect 303985 337807 304043 337813
rect 303985 337773 303997 337807
rect 304031 337804 304043 337807
rect 318797 337807 318855 337813
rect 318797 337804 318809 337807
rect 304031 337776 318809 337804
rect 304031 337773 304043 337776
rect 303985 337767 304043 337773
rect 318797 337773 318809 337776
rect 318843 337773 318855 337807
rect 318797 337767 318855 337773
rect 318981 337807 319039 337813
rect 318981 337773 318993 337807
rect 319027 337804 319039 337807
rect 351914 337804 351920 337816
rect 319027 337776 351920 337804
rect 319027 337773 319039 337776
rect 318981 337767 319039 337773
rect 351914 337764 351920 337776
rect 351972 337764 351978 337816
rect 362862 337764 362868 337816
rect 362920 337804 362926 337816
rect 370332 337804 370360 337844
rect 378870 337832 378876 337844
rect 378928 337832 378934 337884
rect 388438 337832 388444 337884
rect 388496 337872 388502 337884
rect 389174 337872 389180 337884
rect 388496 337844 389180 337872
rect 388496 337832 388502 337844
rect 389174 337832 389180 337844
rect 389232 337832 389238 337884
rect 404814 337832 404820 337884
rect 404872 337872 404878 337884
rect 412545 337875 412603 337881
rect 412545 337872 412557 337875
rect 404872 337844 412557 337872
rect 404872 337832 404878 337844
rect 412545 337841 412557 337844
rect 412591 337841 412603 337875
rect 412545 337835 412603 337841
rect 413848 337844 416820 337872
rect 377398 337804 377404 337816
rect 362920 337776 370360 337804
rect 370424 337776 377404 337804
rect 362920 337764 362926 337776
rect 39298 337696 39304 337748
rect 39356 337736 39362 337748
rect 57974 337736 57980 337748
rect 39356 337708 57980 337736
rect 39356 337696 39362 337708
rect 57974 337696 57980 337708
rect 58032 337696 58038 337748
rect 67542 337696 67548 337748
rect 67600 337736 67606 337748
rect 77294 337736 77300 337748
rect 67600 337708 77300 337736
rect 67600 337696 67606 337708
rect 77294 337696 77300 337708
rect 77352 337696 77358 337748
rect 86862 337696 86868 337748
rect 86920 337736 86926 337748
rect 95234 337736 95240 337748
rect 86920 337708 95240 337736
rect 86920 337696 86926 337708
rect 95234 337696 95240 337708
rect 95292 337696 95298 337748
rect 104802 337696 104808 337748
rect 104860 337736 104866 337748
rect 114554 337736 114560 337748
rect 104860 337708 114560 337736
rect 104860 337696 104866 337708
rect 114554 337696 114560 337708
rect 114612 337696 114618 337748
rect 124122 337696 124128 337748
rect 124180 337736 124186 337748
rect 133874 337736 133880 337748
rect 124180 337708 133880 337736
rect 124180 337696 124186 337708
rect 133874 337696 133880 337708
rect 133932 337696 133938 337748
rect 143442 337696 143448 337748
rect 143500 337736 143506 337748
rect 153194 337736 153200 337748
rect 143500 337708 153200 337736
rect 143500 337696 143506 337708
rect 153194 337696 153200 337708
rect 153252 337696 153258 337748
rect 162762 337696 162768 337748
rect 162820 337736 162826 337748
rect 172514 337736 172520 337748
rect 162820 337708 172520 337736
rect 162820 337696 162826 337708
rect 172514 337696 172520 337708
rect 172572 337696 172578 337748
rect 182082 337696 182088 337748
rect 182140 337736 182146 337748
rect 191834 337736 191840 337748
rect 182140 337708 191840 337736
rect 182140 337696 182146 337708
rect 191834 337696 191840 337708
rect 191892 337696 191898 337748
rect 201402 337696 201408 337748
rect 201460 337736 201466 337748
rect 211154 337736 211160 337748
rect 201460 337708 211160 337736
rect 201460 337696 201466 337708
rect 211154 337696 211160 337708
rect 211212 337696 211218 337748
rect 220722 337696 220728 337748
rect 220780 337736 220786 337748
rect 229097 337739 229155 337745
rect 229097 337736 229109 337739
rect 220780 337708 229109 337736
rect 220780 337696 220786 337708
rect 229097 337705 229109 337708
rect 229143 337705 229155 337739
rect 229097 337699 229155 337705
rect 238680 337708 238800 337736
rect 32398 337628 32404 337680
rect 32456 337668 32462 337680
rect 87049 337671 87107 337677
rect 87049 337668 87061 337671
rect 32456 337640 87061 337668
rect 32456 337628 32462 337640
rect 87049 337637 87061 337640
rect 87095 337637 87107 337671
rect 87049 337631 87107 337637
rect 87417 337671 87475 337677
rect 87417 337637 87429 337671
rect 87463 337668 87475 337671
rect 230569 337671 230627 337677
rect 230569 337668 230581 337671
rect 87463 337640 230581 337668
rect 87463 337637 87475 337640
rect 87417 337631 87475 337637
rect 230569 337637 230581 337640
rect 230615 337637 230627 337671
rect 230569 337631 230627 337637
rect 230658 337628 230664 337680
rect 230716 337668 230722 337680
rect 231118 337668 231124 337680
rect 230716 337640 231124 337668
rect 230716 337628 230722 337640
rect 231118 337628 231124 337640
rect 231176 337628 231182 337680
rect 238680 337677 238708 337708
rect 238772 337677 238800 337708
rect 254578 337696 254584 337748
rect 254636 337736 254642 337748
rect 262306 337736 262312 337748
rect 254636 337708 262312 337736
rect 254636 337696 254642 337708
rect 262306 337696 262312 337708
rect 262364 337696 262370 337748
rect 302237 337739 302295 337745
rect 302237 337705 302249 337739
rect 302283 337736 302295 337739
rect 307754 337736 307760 337748
rect 302283 337708 307760 337736
rect 302283 337705 302295 337708
rect 302237 337699 302295 337705
rect 307754 337696 307760 337708
rect 307812 337696 307818 337748
rect 317322 337696 317328 337748
rect 317380 337736 317386 337748
rect 327077 337739 327135 337745
rect 327077 337736 327089 337739
rect 317380 337708 327089 337736
rect 317380 337696 317386 337708
rect 327077 337705 327089 337708
rect 327123 337705 327135 337739
rect 327077 337699 327135 337705
rect 336645 337739 336703 337745
rect 336645 337705 336657 337739
rect 336691 337736 336703 337739
rect 346397 337739 346455 337745
rect 346397 337736 346409 337739
rect 336691 337708 346409 337736
rect 336691 337705 336703 337708
rect 336645 337699 336703 337705
rect 346397 337705 346409 337708
rect 346443 337705 346455 337739
rect 346397 337699 346455 337705
rect 356698 337696 356704 337748
rect 356756 337736 356762 337748
rect 360746 337736 360752 337748
rect 356756 337708 360752 337736
rect 356756 337696 356762 337708
rect 360746 337696 360752 337708
rect 360804 337696 360810 337748
rect 370424 337736 370452 337776
rect 377398 337764 377404 337776
rect 377456 337764 377462 337816
rect 404354 337764 404360 337816
rect 404412 337804 404418 337816
rect 413848 337804 413876 337844
rect 404412 337776 413876 337804
rect 404412 337764 404418 337776
rect 416130 337764 416136 337816
rect 416188 337804 416194 337816
rect 416682 337804 416688 337816
rect 416188 337776 416688 337804
rect 416188 337764 416194 337776
rect 416682 337764 416688 337776
rect 416740 337764 416746 337816
rect 416792 337804 416820 337844
rect 417602 337832 417608 337884
rect 417660 337872 417666 337884
rect 451384 337872 451412 337912
rect 455598 337900 455604 337912
rect 455656 337900 455662 337952
rect 458726 337900 458732 337952
rect 458784 337940 458790 337952
rect 459370 337940 459376 337952
rect 458784 337912 459376 337940
rect 458784 337900 458790 337912
rect 459370 337900 459376 337912
rect 459428 337900 459434 337952
rect 467098 337900 467104 337952
rect 467156 337940 467162 337952
rect 467742 337940 467748 337952
rect 467156 337912 467748 337940
rect 467156 337900 467162 337912
rect 467742 337900 467748 337912
rect 467800 337900 467806 337952
rect 468018 337900 468024 337952
rect 468076 337940 468082 337952
rect 469122 337940 469128 337952
rect 468076 337912 469128 337940
rect 468076 337900 468082 337912
rect 469122 337900 469128 337912
rect 469180 337900 469186 337952
rect 469217 337943 469275 337949
rect 469217 337909 469229 337943
rect 469263 337940 469275 337943
rect 527818 337940 527824 337952
rect 469263 337912 527824 337940
rect 469263 337909 469275 337912
rect 469217 337903 469275 337909
rect 527818 337900 527824 337912
rect 527876 337900 527882 337952
rect 417660 337844 451412 337872
rect 451461 337875 451519 337881
rect 417660 337832 417666 337844
rect 451461 337841 451473 337875
rect 451507 337872 451519 337875
rect 461397 337875 461455 337881
rect 461397 337872 461409 337875
rect 451507 337844 461409 337872
rect 451507 337841 451519 337844
rect 451461 337835 451519 337841
rect 461397 337841 461409 337844
rect 461443 337841 461455 337875
rect 523678 337872 523684 337884
rect 461397 337835 461455 337841
rect 461504 337844 523684 337872
rect 420270 337804 420276 337816
rect 416792 337776 420276 337804
rect 420270 337764 420276 337776
rect 420328 337764 420334 337816
rect 422018 337764 422024 337816
rect 422076 337804 422082 337816
rect 438118 337804 438124 337816
rect 422076 337776 438124 337804
rect 422076 337764 422082 337776
rect 438118 337764 438124 337776
rect 438176 337764 438182 337816
rect 438670 337764 438676 337816
rect 438728 337804 438734 337816
rect 438728 337776 440280 337804
rect 438728 337764 438734 337776
rect 375926 337736 375932 337748
rect 361592 337708 370452 337736
rect 370516 337708 375932 337736
rect 231213 337671 231271 337677
rect 231213 337637 231225 337671
rect 231259 337668 231271 337671
rect 234433 337671 234491 337677
rect 234433 337668 234445 337671
rect 231259 337640 234445 337668
rect 231259 337637 231271 337640
rect 231213 337631 231271 337637
rect 234433 337637 234445 337640
rect 234479 337637 234491 337671
rect 234433 337631 234491 337637
rect 238665 337671 238723 337677
rect 238665 337637 238677 337671
rect 238711 337637 238723 337671
rect 238665 337631 238723 337637
rect 238757 337671 238815 337677
rect 238757 337637 238769 337671
rect 238803 337637 238815 337671
rect 238757 337631 238815 337637
rect 255958 337628 255964 337680
rect 256016 337668 256022 337680
rect 259733 337671 259791 337677
rect 259733 337668 259745 337671
rect 256016 337640 259745 337668
rect 256016 337628 256022 337640
rect 259733 337637 259745 337640
rect 259779 337637 259791 337671
rect 259733 337631 259791 337637
rect 260098 337628 260104 337680
rect 260156 337668 260162 337680
rect 277026 337668 277032 337680
rect 260156 337640 277032 337668
rect 260156 337628 260162 337640
rect 277026 337628 277032 337640
rect 277084 337628 277090 337680
rect 285582 337628 285588 337680
rect 285640 337668 285646 337680
rect 336001 337671 336059 337677
rect 336001 337668 336013 337671
rect 285640 337640 336013 337668
rect 285640 337628 285646 337640
rect 336001 337637 336013 337640
rect 336047 337637 336059 337671
rect 336001 337631 336059 337637
rect 336090 337628 336096 337680
rect 336148 337668 336154 337680
rect 344554 337668 344560 337680
rect 336148 337640 344560 337668
rect 336148 337628 336154 337640
rect 344554 337628 344560 337640
rect 344612 337628 344618 337680
rect 344649 337671 344707 337677
rect 344649 337637 344661 337671
rect 344695 337668 344707 337671
rect 349982 337668 349988 337680
rect 344695 337640 349988 337668
rect 344695 337637 344707 337640
rect 344649 337631 344707 337637
rect 349982 337628 349988 337640
rect 350040 337628 350046 337680
rect 354858 337668 354864 337680
rect 350276 337640 354864 337668
rect 35158 337560 35164 337612
rect 35216 337600 35222 337612
rect 115661 337603 115719 337609
rect 115661 337600 115673 337603
rect 35216 337572 115673 337600
rect 35216 337560 35222 337572
rect 115661 337569 115673 337572
rect 115707 337569 115719 337603
rect 115661 337563 115719 337569
rect 115845 337603 115903 337609
rect 115845 337569 115857 337603
rect 115891 337600 115903 337603
rect 134981 337603 135039 337609
rect 134981 337600 134993 337603
rect 115891 337572 134993 337600
rect 115891 337569 115903 337572
rect 115845 337563 115903 337569
rect 134981 337569 134993 337572
rect 135027 337569 135039 337603
rect 134981 337563 135039 337569
rect 135165 337603 135223 337609
rect 135165 337569 135177 337603
rect 135211 337600 135223 337603
rect 154301 337603 154359 337609
rect 154301 337600 154313 337603
rect 135211 337572 154313 337600
rect 135211 337569 135223 337572
rect 135165 337563 135223 337569
rect 154301 337569 154313 337572
rect 154347 337569 154359 337603
rect 154301 337563 154359 337569
rect 154485 337603 154543 337609
rect 154485 337569 154497 337603
rect 154531 337600 154543 337603
rect 173621 337603 173679 337609
rect 173621 337600 173633 337603
rect 154531 337572 173633 337600
rect 154531 337569 154543 337572
rect 154485 337563 154543 337569
rect 173621 337569 173633 337572
rect 173667 337569 173679 337603
rect 173621 337563 173679 337569
rect 173805 337603 173863 337609
rect 173805 337569 173817 337603
rect 173851 337600 173863 337603
rect 192941 337603 192999 337609
rect 192941 337600 192953 337603
rect 173851 337572 192953 337600
rect 173851 337569 173863 337572
rect 173805 337563 173863 337569
rect 192941 337569 192953 337572
rect 192987 337569 192999 337603
rect 192941 337563 192999 337569
rect 193125 337603 193183 337609
rect 193125 337569 193137 337603
rect 193171 337600 193183 337603
rect 212261 337603 212319 337609
rect 212261 337600 212273 337603
rect 193171 337572 212273 337600
rect 193171 337569 193183 337572
rect 193125 337563 193183 337569
rect 212261 337569 212273 337572
rect 212307 337569 212319 337603
rect 212261 337563 212319 337569
rect 212445 337603 212503 337609
rect 212445 337569 212457 337603
rect 212491 337600 212503 337603
rect 220909 337603 220967 337609
rect 220909 337600 220921 337603
rect 212491 337572 220921 337600
rect 212491 337569 212503 337572
rect 212445 337563 212503 337569
rect 220909 337569 220921 337572
rect 220955 337569 220967 337603
rect 220909 337563 220967 337569
rect 221093 337603 221151 337609
rect 221093 337569 221105 337603
rect 221139 337600 221151 337603
rect 241698 337600 241704 337612
rect 221139 337572 241704 337600
rect 221139 337569 221151 337572
rect 221093 337563 221151 337569
rect 241698 337560 241704 337572
rect 241756 337560 241762 337612
rect 261386 337560 261392 337612
rect 261444 337600 261450 337612
rect 279970 337600 279976 337612
rect 261444 337572 279976 337600
rect 261444 337560 261450 337572
rect 279970 337560 279976 337572
rect 280028 337560 280034 337612
rect 281442 337560 281448 337612
rect 281500 337600 281506 337612
rect 318889 337603 318947 337609
rect 318889 337600 318901 337603
rect 281500 337572 318901 337600
rect 281500 337560 281506 337572
rect 318889 337569 318901 337572
rect 318935 337569 318947 337603
rect 318889 337563 318947 337569
rect 318981 337603 319039 337609
rect 318981 337569 318993 337603
rect 319027 337600 319039 337603
rect 345566 337600 345572 337612
rect 319027 337572 345572 337600
rect 319027 337569 319039 337572
rect 318981 337563 319039 337569
rect 345566 337560 345572 337572
rect 345624 337560 345630 337612
rect 345750 337560 345756 337612
rect 345808 337600 345814 337612
rect 350166 337600 350172 337612
rect 345808 337572 350172 337600
rect 345808 337560 345814 337572
rect 350166 337560 350172 337572
rect 350224 337560 350230 337612
rect 28258 337492 28264 337544
rect 28316 337532 28322 337544
rect 220814 337532 220820 337544
rect 28316 337504 220820 337532
rect 28316 337492 28322 337504
rect 220814 337492 220820 337504
rect 220872 337492 220878 337544
rect 220998 337492 221004 337544
rect 221056 337532 221062 337544
rect 230477 337535 230535 337541
rect 230477 337532 230489 337535
rect 221056 337504 230489 337532
rect 221056 337492 221062 337504
rect 230477 337501 230489 337504
rect 230523 337501 230535 337535
rect 230477 337495 230535 337501
rect 230569 337535 230627 337541
rect 230569 337501 230581 337535
rect 230615 337532 230627 337535
rect 237834 337532 237840 337544
rect 230615 337504 237840 337532
rect 230615 337501 230627 337504
rect 230569 337495 230627 337501
rect 237834 337492 237840 337504
rect 237892 337492 237898 337544
rect 253198 337492 253204 337544
rect 253256 337532 253262 337544
rect 259362 337532 259368 337544
rect 253256 337504 259368 337532
rect 253256 337492 253262 337504
rect 259362 337492 259368 337504
rect 259420 337492 259426 337544
rect 275554 337532 275560 337544
rect 259472 337504 275560 337532
rect 19978 337424 19984 337476
rect 20036 337464 20042 337476
rect 87049 337467 87107 337473
rect 87049 337464 87061 337467
rect 20036 337436 87061 337464
rect 20036 337424 20042 337436
rect 87049 337433 87061 337436
rect 87095 337433 87107 337467
rect 87049 337427 87107 337433
rect 87141 337467 87199 337473
rect 87141 337433 87153 337467
rect 87187 337464 87199 337467
rect 220909 337467 220967 337473
rect 220909 337464 220921 337467
rect 87187 337436 220921 337464
rect 87187 337433 87199 337436
rect 87141 337427 87199 337433
rect 220909 337433 220921 337436
rect 220955 337433 220967 337467
rect 220909 337427 220967 337433
rect 221093 337467 221151 337473
rect 221093 337433 221105 337467
rect 221139 337464 221151 337467
rect 234338 337464 234344 337476
rect 221139 337436 234344 337464
rect 221139 337433 221151 337436
rect 221093 337427 221151 337433
rect 234338 337424 234344 337436
rect 234396 337424 234402 337476
rect 234433 337467 234491 337473
rect 234433 337433 234445 337467
rect 234479 337464 234491 337467
rect 238294 337464 238300 337476
rect 234479 337436 238300 337464
rect 234479 337433 234491 337436
rect 234433 337427 234491 337433
rect 238294 337424 238300 337436
rect 238352 337424 238358 337476
rect 258810 337424 258816 337476
rect 258868 337464 258874 337476
rect 259472 337464 259500 337504
rect 275554 337492 275560 337504
rect 275612 337492 275618 337544
rect 275922 337492 275928 337544
rect 275980 337532 275986 337544
rect 335817 337535 335875 337541
rect 335817 337532 335829 337535
rect 275980 337504 335829 337532
rect 275980 337492 275986 337504
rect 335817 337501 335829 337504
rect 335863 337501 335875 337535
rect 341610 337532 341616 337544
rect 335817 337495 335875 337501
rect 336016 337504 341616 337532
rect 269666 337464 269672 337476
rect 258868 337436 259500 337464
rect 259656 337436 269672 337464
rect 258868 337424 258874 337436
rect 13078 337356 13084 337408
rect 13136 337396 13142 337408
rect 220814 337396 220820 337408
rect 13136 337368 220820 337396
rect 13136 337356 13142 337368
rect 220814 337356 220820 337368
rect 220872 337356 220878 337408
rect 220998 337356 221004 337408
rect 221056 337396 221062 337408
rect 233510 337396 233516 337408
rect 221056 337368 233516 337396
rect 221056 337356 221062 337368
rect 233510 337356 233516 337368
rect 233568 337356 233574 337408
rect 233878 337356 233884 337408
rect 233936 337396 233942 337408
rect 241238 337396 241244 337408
rect 233936 337368 241244 337396
rect 233936 337356 233942 337368
rect 241238 337356 241244 337368
rect 241296 337356 241302 337408
rect 250438 337356 250444 337408
rect 250496 337396 250502 337408
rect 253474 337396 253480 337408
rect 250496 337368 253480 337396
rect 250496 337356 250502 337368
rect 253474 337356 253480 337368
rect 253532 337356 253538 337408
rect 257338 337356 257344 337408
rect 257396 337396 257402 337408
rect 259656 337396 259684 337436
rect 269666 337424 269672 337436
rect 269724 337424 269730 337476
rect 271782 337424 271788 337476
rect 271840 337464 271846 337476
rect 318797 337467 318855 337473
rect 318797 337464 318809 337467
rect 271840 337436 318809 337464
rect 271840 337424 271846 337436
rect 318797 337433 318809 337436
rect 318843 337433 318855 337467
rect 318797 337427 318855 337433
rect 319073 337467 319131 337473
rect 319073 337433 319085 337467
rect 319119 337464 319131 337467
rect 336016 337464 336044 337504
rect 341610 337492 341616 337504
rect 341668 337492 341674 337544
rect 341705 337535 341763 337541
rect 341705 337501 341717 337535
rect 341751 337532 341763 337535
rect 342714 337532 342720 337544
rect 341751 337504 342720 337532
rect 341751 337501 341763 337504
rect 341705 337495 341763 337501
rect 342714 337492 342720 337504
rect 342772 337492 342778 337544
rect 342809 337535 342867 337541
rect 342809 337501 342821 337535
rect 342855 337532 342867 337535
rect 344189 337535 344247 337541
rect 344189 337532 344201 337535
rect 342855 337504 344201 337532
rect 342855 337501 342867 337504
rect 342809 337495 342867 337501
rect 344189 337501 344201 337504
rect 344235 337501 344247 337535
rect 344189 337495 344247 337501
rect 344278 337492 344284 337544
rect 344336 337532 344342 337544
rect 350276 337532 350304 337640
rect 354858 337628 354864 337640
rect 354916 337628 354922 337680
rect 358722 337628 358728 337680
rect 358780 337668 358786 337680
rect 361592 337668 361620 337708
rect 358780 337640 361620 337668
rect 364981 337671 365039 337677
rect 358780 337628 358786 337640
rect 364981 337637 364993 337671
rect 365027 337668 365039 337671
rect 370516 337668 370544 337708
rect 375926 337696 375932 337708
rect 375984 337696 375990 337748
rect 380158 337696 380164 337748
rect 380216 337736 380222 337748
rect 381354 337736 381360 337748
rect 380216 337708 381360 337736
rect 380216 337696 380222 337708
rect 381354 337696 381360 337708
rect 381412 337696 381418 337748
rect 381538 337696 381544 337748
rect 381596 337736 381602 337748
rect 382826 337736 382832 337748
rect 381596 337708 382832 337736
rect 381596 337696 381602 337708
rect 382826 337696 382832 337708
rect 382884 337696 382890 337748
rect 384942 337696 384948 337748
rect 385000 337736 385006 337748
rect 388162 337736 388168 337748
rect 385000 337708 388168 337736
rect 385000 337696 385006 337708
rect 388162 337696 388168 337708
rect 388220 337696 388226 337748
rect 399478 337696 399484 337748
rect 399536 337736 399542 337748
rect 400122 337736 400128 337748
rect 399536 337708 400128 337736
rect 399536 337696 399542 337708
rect 400122 337696 400128 337708
rect 400180 337696 400186 337748
rect 402422 337696 402428 337748
rect 402480 337736 402486 337748
rect 402882 337736 402888 337748
rect 402480 337708 402888 337736
rect 402480 337696 402486 337708
rect 402882 337696 402888 337708
rect 402940 337696 402946 337748
rect 403342 337696 403348 337748
rect 403400 337736 403406 337748
rect 403400 337708 410196 337736
rect 403400 337696 403406 337708
rect 365027 337640 370544 337668
rect 376757 337671 376815 337677
rect 365027 337637 365039 337640
rect 364981 337631 365039 337637
rect 376757 337637 376769 337671
rect 376803 337668 376815 337671
rect 380802 337668 380808 337680
rect 376803 337640 380808 337668
rect 376803 337637 376815 337640
rect 376757 337631 376815 337637
rect 380802 337628 380808 337640
rect 380860 337628 380866 337680
rect 384298 337628 384304 337680
rect 384356 337668 384362 337680
rect 387702 337668 387708 337680
rect 384356 337640 387708 337668
rect 384356 337628 384362 337640
rect 387702 337628 387708 337640
rect 387760 337628 387766 337680
rect 398926 337628 398932 337680
rect 398984 337668 398990 337680
rect 406378 337668 406384 337680
rect 398984 337640 406384 337668
rect 398984 337628 398990 337640
rect 406378 337628 406384 337640
rect 406436 337628 406442 337680
rect 410168 337668 410196 337708
rect 410242 337696 410248 337748
rect 410300 337736 410306 337748
rect 411070 337736 411076 337748
rect 410300 337708 411076 337736
rect 410300 337696 410306 337708
rect 411070 337696 411076 337708
rect 411128 337696 411134 337748
rect 414109 337739 414167 337745
rect 414109 337736 414121 337739
rect 411180 337708 414121 337736
rect 411180 337668 411208 337708
rect 414109 337705 414121 337708
rect 414155 337705 414167 337739
rect 414109 337699 414167 337705
rect 414198 337696 414204 337748
rect 414256 337736 414262 337748
rect 415302 337736 415308 337748
rect 414256 337708 415308 337736
rect 414256 337696 414262 337708
rect 415302 337696 415308 337708
rect 415360 337696 415366 337748
rect 415578 337696 415584 337748
rect 415636 337736 415642 337748
rect 416498 337736 416504 337748
rect 415636 337708 416504 337736
rect 415636 337696 415642 337708
rect 416498 337696 416504 337708
rect 416556 337696 416562 337748
rect 417050 337696 417056 337748
rect 417108 337736 417114 337748
rect 417970 337736 417976 337748
rect 417108 337708 417976 337736
rect 417108 337696 417114 337708
rect 417970 337696 417976 337708
rect 418028 337696 418034 337748
rect 425422 337696 425428 337748
rect 425480 337736 425486 337748
rect 428458 337736 428464 337748
rect 425480 337708 428464 337736
rect 425480 337696 425486 337708
rect 428458 337696 428464 337708
rect 428516 337696 428522 337748
rect 429378 337696 429384 337748
rect 429436 337736 429442 337748
rect 430482 337736 430488 337748
rect 429436 337708 430488 337736
rect 429436 337696 429442 337708
rect 430482 337696 430488 337708
rect 430540 337696 430546 337748
rect 432233 337739 432291 337745
rect 432233 337736 432245 337739
rect 430592 337708 432245 337736
rect 410168 337640 411208 337668
rect 411254 337628 411260 337680
rect 411312 337668 411318 337680
rect 412358 337668 412364 337680
rect 411312 337640 412364 337668
rect 411312 337628 411318 337640
rect 412358 337628 412364 337640
rect 412416 337628 412422 337680
rect 427078 337668 427084 337680
rect 412468 337640 427084 337668
rect 351178 337560 351184 337612
rect 351236 337600 351242 337612
rect 365165 337603 365223 337609
rect 365165 337600 365177 337603
rect 351236 337572 365177 337600
rect 351236 337560 351242 337572
rect 365165 337569 365177 337572
rect 365211 337569 365223 337603
rect 365165 337563 365223 337569
rect 367002 337560 367008 337612
rect 367060 337600 367066 337612
rect 374641 337603 374699 337609
rect 374641 337600 374653 337603
rect 367060 337572 374653 337600
rect 367060 337560 367066 337572
rect 374641 337569 374653 337572
rect 374687 337569 374699 337603
rect 383286 337600 383292 337612
rect 374641 337563 374699 337569
rect 374748 337572 383292 337600
rect 344336 337504 350304 337532
rect 344336 337492 344342 337504
rect 351822 337492 351828 337544
rect 351880 337532 351886 337544
rect 365073 337535 365131 337541
rect 365073 337532 365085 337535
rect 351880 337504 365085 337532
rect 351880 337492 351886 337504
rect 365073 337501 365085 337504
rect 365119 337501 365131 337535
rect 365073 337495 365131 337501
rect 365257 337535 365315 337541
rect 365257 337501 365269 337535
rect 365303 337532 365315 337535
rect 365303 337504 372200 337532
rect 365303 337501 365315 337504
rect 365257 337495 365315 337501
rect 344094 337464 344100 337476
rect 319119 337436 336044 337464
rect 336108 337436 344100 337464
rect 319119 337433 319131 337436
rect 319073 337427 319131 337433
rect 257396 337368 259684 337396
rect 259733 337399 259791 337405
rect 257396 337356 257402 337368
rect 259733 337365 259745 337399
rect 259779 337396 259791 337399
rect 266722 337396 266728 337408
rect 259779 337368 266728 337396
rect 259779 337365 259791 337368
rect 259733 337359 259791 337365
rect 266722 337356 266728 337368
rect 266780 337356 266786 337408
rect 269022 337356 269028 337408
rect 269080 337396 269086 337408
rect 334713 337399 334771 337405
rect 334713 337396 334725 337399
rect 269080 337368 334725 337396
rect 269080 337356 269086 337368
rect 334713 337365 334725 337368
rect 334759 337365 334771 337399
rect 334713 337359 334771 337365
rect 335909 337399 335967 337405
rect 335909 337365 335921 337399
rect 335955 337396 335967 337399
rect 336108 337396 336136 337436
rect 344094 337424 344100 337436
rect 344152 337424 344158 337476
rect 347498 337464 347504 337476
rect 344204 337436 347504 337464
rect 335955 337368 336136 337396
rect 336185 337399 336243 337405
rect 335955 337365 335967 337368
rect 335909 337359 335967 337365
rect 336185 337365 336197 337399
rect 336231 337396 336243 337399
rect 340785 337399 340843 337405
rect 340785 337396 340797 337399
rect 336231 337368 340797 337396
rect 336231 337365 336243 337368
rect 336185 337359 336243 337365
rect 340785 337365 340797 337368
rect 340831 337365 340843 337399
rect 340785 337359 340843 337365
rect 340877 337399 340935 337405
rect 340877 337365 340889 337399
rect 340923 337396 340935 337399
rect 344204 337396 344232 337436
rect 347498 337424 347504 337436
rect 347556 337424 347562 337476
rect 349062 337424 349068 337476
rect 349120 337464 349126 337476
rect 372172 337464 372200 337504
rect 373902 337492 373908 337544
rect 373960 337532 373966 337544
rect 374748 337532 374776 337572
rect 383286 337560 383292 337572
rect 383344 337560 383350 337612
rect 398006 337560 398012 337612
rect 398064 337600 398070 337612
rect 399478 337600 399484 337612
rect 398064 337572 399484 337600
rect 398064 337560 398070 337572
rect 399478 337560 399484 337572
rect 399536 337560 399542 337612
rect 407298 337560 407304 337612
rect 407356 337600 407362 337612
rect 412468 337600 412496 337640
rect 427078 337628 427084 337640
rect 427136 337628 427142 337680
rect 430592 337668 430620 337708
rect 432233 337705 432245 337708
rect 432279 337705 432291 337739
rect 432233 337699 432291 337705
rect 432322 337696 432328 337748
rect 432380 337736 432386 337748
rect 433242 337736 433248 337748
rect 432380 337708 433248 337736
rect 432380 337696 432386 337708
rect 433242 337696 433248 337708
rect 433300 337696 433306 337748
rect 433702 337696 433708 337748
rect 433760 337736 433766 337748
rect 434622 337736 434628 337748
rect 433760 337708 434628 337736
rect 433760 337696 433766 337708
rect 434622 337696 434628 337708
rect 434680 337696 434686 337748
rect 435174 337696 435180 337748
rect 435232 337736 435238 337748
rect 436002 337736 436008 337748
rect 435232 337708 436008 337736
rect 435232 337696 435238 337708
rect 436002 337696 436008 337708
rect 436060 337696 436066 337748
rect 436646 337696 436652 337748
rect 436704 337736 436710 337748
rect 437382 337736 437388 337748
rect 436704 337708 437388 337736
rect 436704 337696 436710 337708
rect 437382 337696 437388 337708
rect 437440 337696 437446 337748
rect 437658 337696 437664 337748
rect 437716 337736 437722 337748
rect 438762 337736 438768 337748
rect 437716 337708 438768 337736
rect 437716 337696 437722 337708
rect 438762 337696 438768 337708
rect 438820 337696 438826 337748
rect 439130 337696 439136 337748
rect 439188 337736 439194 337748
rect 440142 337736 440148 337748
rect 439188 337708 440148 337736
rect 439188 337696 439194 337708
rect 440142 337696 440148 337708
rect 440200 337696 440206 337748
rect 440252 337736 440280 337776
rect 440602 337764 440608 337816
rect 440660 337804 440666 337816
rect 441522 337804 441528 337816
rect 440660 337776 441528 337804
rect 440660 337764 440666 337776
rect 441522 337764 441528 337776
rect 441580 337764 441586 337816
rect 441614 337764 441620 337816
rect 441672 337804 441678 337816
rect 443638 337804 443644 337816
rect 441672 337776 443644 337804
rect 441672 337764 441678 337776
rect 443638 337764 443644 337776
rect 443696 337764 443702 337816
rect 444558 337764 444564 337816
rect 444616 337804 444622 337816
rect 445662 337804 445668 337816
rect 444616 337776 445668 337804
rect 444616 337764 444622 337776
rect 445662 337764 445668 337776
rect 445720 337764 445726 337816
rect 446401 337807 446459 337813
rect 446401 337773 446413 337807
rect 446447 337804 446459 337807
rect 448517 337807 448575 337813
rect 448517 337804 448529 337807
rect 446447 337776 448529 337804
rect 446447 337773 446459 337776
rect 446401 337767 446459 337773
rect 448517 337773 448529 337776
rect 448563 337773 448575 337807
rect 448517 337767 448575 337773
rect 448974 337764 448980 337816
rect 449032 337804 449038 337816
rect 449032 337776 451228 337804
rect 449032 337764 449038 337776
rect 449161 337739 449219 337745
rect 449161 337736 449173 337739
rect 440252 337708 449173 337736
rect 449161 337705 449173 337708
rect 449207 337705 449219 337739
rect 449161 337699 449219 337705
rect 428292 337640 430620 337668
rect 407356 337572 412496 337600
rect 412545 337603 412603 337609
rect 407356 337560 407362 337572
rect 412545 337569 412557 337603
rect 412591 337600 412603 337603
rect 424686 337600 424692 337612
rect 412591 337572 424692 337600
rect 412591 337569 412603 337572
rect 412545 337563 412603 337569
rect 424686 337560 424692 337572
rect 424744 337560 424750 337612
rect 426434 337560 426440 337612
rect 426492 337600 426498 337612
rect 428292 337600 428320 337640
rect 430850 337628 430856 337680
rect 430908 337668 430914 337680
rect 431862 337668 431868 337680
rect 430908 337640 431868 337668
rect 430908 337628 430914 337640
rect 431862 337628 431868 337640
rect 431920 337628 431926 337680
rect 434714 337628 434720 337680
rect 434772 337668 434778 337680
rect 435910 337668 435916 337680
rect 434772 337640 435916 337668
rect 434772 337628 434778 337640
rect 435910 337628 435916 337640
rect 435968 337628 435974 337680
rect 436186 337628 436192 337680
rect 436244 337668 436250 337680
rect 437290 337668 437296 337680
rect 436244 337640 437296 337668
rect 436244 337628 436250 337640
rect 437290 337628 437296 337640
rect 437348 337628 437354 337680
rect 437492 337640 441844 337668
rect 426492 337572 428320 337600
rect 426492 337560 426498 337572
rect 428366 337560 428372 337612
rect 428424 337600 428430 337612
rect 431218 337600 431224 337612
rect 428424 337572 431224 337600
rect 428424 337560 428430 337572
rect 431218 337560 431224 337572
rect 431276 337560 431282 337612
rect 431310 337560 431316 337612
rect 431368 337600 431374 337612
rect 437385 337603 437443 337609
rect 437385 337600 437397 337603
rect 431368 337572 437397 337600
rect 431368 337560 431374 337572
rect 437385 337569 437397 337572
rect 437431 337569 437443 337603
rect 437385 337563 437443 337569
rect 373960 337504 374776 337532
rect 373960 337492 373966 337504
rect 375282 337492 375288 337544
rect 375340 337532 375346 337544
rect 383746 337532 383752 337544
rect 375340 337504 383752 337532
rect 375340 337492 375346 337504
rect 383746 337492 383752 337504
rect 383804 337492 383810 337544
rect 405826 337492 405832 337544
rect 405884 337532 405890 337544
rect 405884 337504 422340 337532
rect 405884 337492 405890 337504
rect 374454 337464 374460 337476
rect 349120 337436 364564 337464
rect 372172 337436 374460 337464
rect 349120 337424 349126 337436
rect 340923 337368 344232 337396
rect 345569 337399 345627 337405
rect 340923 337365 340935 337368
rect 340877 337359 340935 337365
rect 345569 337365 345581 337399
rect 345615 337396 345627 337399
rect 354033 337399 354091 337405
rect 354033 337396 354045 337399
rect 345615 337368 354045 337396
rect 345615 337365 345627 337368
rect 345569 337359 345627 337365
rect 354033 337365 354045 337368
rect 354079 337365 354091 337399
rect 354033 337359 354091 337365
rect 79318 337288 79324 337340
rect 79376 337328 79382 337340
rect 220909 337331 220967 337337
rect 220909 337328 220921 337331
rect 79376 337300 220921 337328
rect 79376 337288 79382 337300
rect 220909 337297 220921 337300
rect 220955 337297 220967 337331
rect 220909 337291 220967 337297
rect 221093 337331 221151 337337
rect 221093 337297 221105 337331
rect 221139 337328 221151 337331
rect 260834 337328 260840 337340
rect 221139 337300 260840 337328
rect 221139 337297 221151 337300
rect 221093 337291 221151 337297
rect 260834 337288 260840 337300
rect 260892 337288 260898 337340
rect 272610 337328 272616 337340
rect 268120 337300 272616 337328
rect 103425 337263 103483 337269
rect 103425 337229 103437 337263
rect 103471 337260 103483 337263
rect 113177 337263 113235 337269
rect 113177 337260 113189 337263
rect 103471 337232 113189 337260
rect 103471 337229 103483 337232
rect 103425 337223 103483 337229
rect 113177 337229 113189 337232
rect 113223 337229 113235 337263
rect 113177 337223 113235 337229
rect 122745 337263 122803 337269
rect 122745 337229 122757 337263
rect 122791 337260 122803 337263
rect 132494 337260 132500 337272
rect 122791 337232 132500 337260
rect 122791 337229 122803 337232
rect 122745 337223 122803 337229
rect 132494 337220 132500 337232
rect 132552 337220 132558 337272
rect 142062 337220 142068 337272
rect 142120 337260 142126 337272
rect 151814 337260 151820 337272
rect 142120 337232 151820 337260
rect 142120 337220 142126 337232
rect 151814 337220 151820 337232
rect 151872 337220 151878 337272
rect 161382 337220 161388 337272
rect 161440 337260 161446 337272
rect 171134 337260 171140 337272
rect 161440 337232 171140 337260
rect 161440 337220 161446 337232
rect 171134 337220 171140 337232
rect 171192 337220 171198 337272
rect 180702 337220 180708 337272
rect 180760 337260 180766 337272
rect 190454 337260 190460 337272
rect 180760 337232 190460 337260
rect 180760 337220 180766 337232
rect 190454 337220 190460 337232
rect 190512 337220 190518 337272
rect 200022 337220 200028 337272
rect 200080 337260 200086 337272
rect 209774 337260 209780 337272
rect 200080 337232 209780 337260
rect 200080 337220 200086 337232
rect 209774 337220 209780 337232
rect 209832 337220 209838 337272
rect 219342 337220 219348 337272
rect 219400 337260 219406 337272
rect 220817 337263 220875 337269
rect 220817 337260 220829 337263
rect 219400 337232 220829 337260
rect 219400 337220 219406 337232
rect 220817 337229 220829 337232
rect 220863 337229 220875 337263
rect 220998 337260 221004 337272
rect 220959 337232 221004 337260
rect 220817 337223 220875 337229
rect 220998 337220 221004 337232
rect 221056 337220 221062 337272
rect 234614 337220 234620 337272
rect 234672 337260 234678 337272
rect 257890 337260 257896 337272
rect 234672 337232 257896 337260
rect 234672 337220 234678 337232
rect 257890 337220 257896 337232
rect 257948 337220 257954 337272
rect 258718 337220 258724 337272
rect 258776 337260 258782 337272
rect 268120 337260 268148 337300
rect 272610 337288 272616 337300
rect 272668 337288 272674 337340
rect 272794 337288 272800 337340
rect 272852 337328 272858 337340
rect 272852 337300 306236 337328
rect 272852 337288 272858 337300
rect 258776 337232 268148 337260
rect 258776 337220 258782 337232
rect 271322 337220 271328 337272
rect 271380 337260 271386 337272
rect 271380 337232 306144 337260
rect 271380 337220 271386 337232
rect 84838 337152 84844 337204
rect 84896 337192 84902 337204
rect 263778 337192 263784 337204
rect 84896 337164 263784 337192
rect 84896 337152 84902 337164
rect 263778 337152 263784 337164
rect 263836 337152 263842 337204
rect 297910 337152 297916 337204
rect 297968 337192 297974 337204
rect 303985 337195 304043 337201
rect 303985 337192 303997 337195
rect 297968 337164 303997 337192
rect 297968 337152 297974 337164
rect 303985 337161 303997 337164
rect 304031 337161 304043 337195
rect 303985 337155 304043 337161
rect 86957 337127 87015 337133
rect 86957 337093 86969 337127
rect 87003 337124 87015 337127
rect 87003 337096 93900 337124
rect 87003 337093 87015 337096
rect 86957 337087 87015 337093
rect 77938 336948 77944 337000
rect 77996 336988 78002 337000
rect 86957 336991 87015 336997
rect 86957 336988 86969 336991
rect 77996 336960 86969 336988
rect 77996 336948 78002 336960
rect 86957 336957 86969 336960
rect 87003 336957 87015 336991
rect 93872 336988 93900 337096
rect 100662 337084 100668 337136
rect 100720 337124 100726 337136
rect 271138 337124 271144 337136
rect 100720 337096 271144 337124
rect 100720 337084 100726 337096
rect 271138 337084 271144 337096
rect 271196 337084 271202 337136
rect 306116 337124 306144 337232
rect 306208 337192 306236 337300
rect 309778 337288 309784 337340
rect 309836 337328 309842 337340
rect 315485 337331 315543 337337
rect 315485 337328 315497 337331
rect 309836 337300 315497 337328
rect 309836 337288 309842 337300
rect 315485 337297 315497 337300
rect 315531 337297 315543 337331
rect 315485 337291 315543 337297
rect 316034 337288 316040 337340
rect 316092 337328 316098 337340
rect 316862 337328 316868 337340
rect 316092 337300 316868 337328
rect 316092 337288 316098 337300
rect 316862 337288 316868 337300
rect 316920 337288 316926 337340
rect 317414 337288 317420 337340
rect 317472 337328 317478 337340
rect 318334 337328 318340 337340
rect 317472 337300 318340 337328
rect 317472 337288 317478 337300
rect 318334 337288 318340 337300
rect 318392 337288 318398 337340
rect 318886 337288 318892 337340
rect 318944 337328 318950 337340
rect 319254 337328 319260 337340
rect 318944 337300 319260 337328
rect 318944 337288 318950 337300
rect 319254 337288 319260 337300
rect 319312 337288 319318 337340
rect 320174 337288 320180 337340
rect 320232 337328 320238 337340
rect 320726 337328 320732 337340
rect 320232 337300 320732 337328
rect 320232 337288 320238 337300
rect 320726 337288 320732 337300
rect 320784 337288 320790 337340
rect 326341 337331 326399 337337
rect 326341 337297 326353 337331
rect 326387 337328 326399 337331
rect 361758 337328 361764 337340
rect 326387 337300 361764 337328
rect 326387 337297 326399 337300
rect 326341 337291 326399 337297
rect 361758 337288 361764 337300
rect 361816 337288 361822 337340
rect 312538 337220 312544 337272
rect 312596 337260 312602 337272
rect 341705 337263 341763 337269
rect 341705 337260 341717 337263
rect 312596 337232 341717 337260
rect 312596 337220 312602 337232
rect 341705 337229 341717 337232
rect 341751 337229 341763 337263
rect 341705 337223 341763 337229
rect 341794 337220 341800 337272
rect 341852 337260 341858 337272
rect 348970 337260 348976 337272
rect 341852 337232 348976 337260
rect 341852 337220 341858 337232
rect 348970 337220 348976 337232
rect 349028 337220 349034 337272
rect 359458 337220 359464 337272
rect 359516 337260 359522 337272
rect 363690 337260 363696 337272
rect 359516 337232 363696 337260
rect 359516 337220 359522 337232
rect 363690 337220 363696 337232
rect 363748 337220 363754 337272
rect 364536 337260 364564 337436
rect 374454 337424 374460 337436
rect 374512 337424 374518 337476
rect 374641 337467 374699 337473
rect 374641 337433 374653 337467
rect 374687 337464 374699 337467
rect 381814 337464 381820 337476
rect 374687 337436 381820 337464
rect 374687 337433 374699 337436
rect 374641 337427 374699 337433
rect 381814 337424 381820 337436
rect 381872 337424 381878 337476
rect 387058 337424 387064 337476
rect 387116 337464 387122 337476
rect 388714 337464 388720 337476
rect 387116 337436 388720 337464
rect 387116 337424 387122 337436
rect 388714 337424 388720 337436
rect 388772 337424 388778 337476
rect 396994 337424 397000 337476
rect 397052 337464 397058 337476
rect 405918 337464 405924 337476
rect 397052 337436 405924 337464
rect 397052 337424 397058 337436
rect 405918 337424 405924 337436
rect 405976 337424 405982 337476
rect 414109 337467 414167 337473
rect 414109 337433 414121 337467
rect 414155 337464 414167 337467
rect 421190 337464 421196 337476
rect 414155 337436 421196 337464
rect 414155 337433 414167 337436
rect 414109 337427 414167 337433
rect 421190 337424 421196 337436
rect 421248 337424 421254 337476
rect 369762 337356 369768 337408
rect 369820 337396 369826 337408
rect 369857 337399 369915 337405
rect 369857 337396 369869 337399
rect 369820 337368 369869 337396
rect 369820 337356 369826 337368
rect 369857 337365 369869 337368
rect 369903 337365 369915 337399
rect 369857 337359 369915 337365
rect 382182 337356 382188 337408
rect 382240 337396 382246 337408
rect 386690 337396 386696 337408
rect 382240 337368 386696 337396
rect 382240 337356 382246 337368
rect 386690 337356 386696 337368
rect 386748 337356 386754 337408
rect 400950 337356 400956 337408
rect 401008 337396 401014 337408
rect 402238 337396 402244 337408
rect 401008 337368 402244 337396
rect 401008 337356 401014 337368
rect 402238 337356 402244 337368
rect 402296 337356 402302 337408
rect 407758 337356 407764 337408
rect 407816 337396 407822 337408
rect 409138 337396 409144 337408
rect 407816 337368 409144 337396
rect 407816 337356 407822 337368
rect 409138 337356 409144 337368
rect 409196 337356 409202 337408
rect 422312 337396 422340 337504
rect 427906 337492 427912 337544
rect 427964 337532 427970 337544
rect 437492 337532 437520 337640
rect 437569 337603 437627 337609
rect 437569 337569 437581 337603
rect 437615 337600 437627 337603
rect 441816 337600 441844 337640
rect 442074 337628 442080 337680
rect 442132 337668 442138 337680
rect 442902 337668 442908 337680
rect 442132 337640 442908 337668
rect 442132 337628 442138 337640
rect 442902 337628 442908 337640
rect 442960 337628 442966 337680
rect 443546 337628 443552 337680
rect 443604 337668 443610 337680
rect 444282 337668 444288 337680
rect 443604 337640 444288 337668
rect 443604 337628 443610 337640
rect 444282 337628 444288 337640
rect 444340 337628 444346 337680
rect 445018 337628 445024 337680
rect 445076 337668 445082 337680
rect 445570 337668 445576 337680
rect 445076 337640 445576 337668
rect 445076 337628 445082 337640
rect 445570 337628 445576 337640
rect 445628 337628 445634 337680
rect 446490 337628 446496 337680
rect 446548 337668 446554 337680
rect 447042 337668 447048 337680
rect 446548 337640 447048 337668
rect 446548 337628 446554 337640
rect 447042 337628 447048 337640
rect 447100 337628 447106 337680
rect 448238 337628 448244 337680
rect 448296 337668 448302 337680
rect 448422 337668 448428 337680
rect 448296 337640 448428 337668
rect 448296 337628 448302 337640
rect 448422 337628 448428 337640
rect 448480 337628 448486 337680
rect 449894 337628 449900 337680
rect 449952 337668 449958 337680
rect 450998 337668 451004 337680
rect 449952 337640 451004 337668
rect 449952 337628 449958 337640
rect 450998 337628 451004 337640
rect 451056 337628 451062 337680
rect 451200 337668 451228 337776
rect 452838 337764 452844 337816
rect 452896 337804 452902 337816
rect 453758 337804 453764 337816
rect 452896 337776 453764 337804
rect 452896 337764 452902 337776
rect 453758 337764 453764 337776
rect 453816 337764 453822 337816
rect 454310 337764 454316 337816
rect 454368 337804 454374 337816
rect 455230 337804 455236 337816
rect 454368 337776 455236 337804
rect 454368 337764 454374 337776
rect 455230 337764 455236 337776
rect 455288 337764 455294 337816
rect 455782 337764 455788 337816
rect 455840 337804 455846 337816
rect 456610 337804 456616 337816
rect 455840 337776 456616 337804
rect 455840 337764 455846 337776
rect 456610 337764 456616 337776
rect 456668 337764 456674 337816
rect 457714 337764 457720 337816
rect 457772 337804 457778 337816
rect 461504 337804 461532 337844
rect 523678 337832 523684 337844
rect 523736 337832 523742 337884
rect 457772 337776 461532 337804
rect 461581 337807 461639 337813
rect 457772 337764 457778 337776
rect 461581 337773 461593 337807
rect 461627 337804 461639 337807
rect 521010 337804 521016 337816
rect 461627 337776 521016 337804
rect 461627 337773 461639 337776
rect 461581 337767 461639 337773
rect 521010 337764 521016 337776
rect 521068 337764 521074 337816
rect 451369 337739 451427 337745
rect 451369 337705 451381 337739
rect 451415 337736 451427 337739
rect 506474 337736 506480 337748
rect 451415 337708 506480 337736
rect 451415 337705 451427 337708
rect 451369 337699 451427 337705
rect 506474 337696 506480 337708
rect 506532 337696 506538 337748
rect 518158 337668 518164 337680
rect 451200 337640 518164 337668
rect 518158 337628 518164 337640
rect 518216 337628 518222 337680
rect 442258 337600 442264 337612
rect 437615 337572 441752 337600
rect 441816 337572 442264 337600
rect 437615 337569 437627 337572
rect 437569 337563 437627 337569
rect 427964 337504 437520 337532
rect 427964 337492 427970 337504
rect 440234 337492 440240 337544
rect 440292 337532 440298 337544
rect 441724 337532 441752 337572
rect 442258 337560 442264 337572
rect 442316 337560 442322 337612
rect 449158 337600 449164 337612
rect 442368 337572 449164 337600
rect 442368 337532 442396 337572
rect 449158 337560 449164 337572
rect 449216 337560 449222 337612
rect 450446 337560 450452 337612
rect 450504 337600 450510 337612
rect 451182 337600 451188 337612
rect 450504 337572 451188 337600
rect 450504 337560 450510 337572
rect 451182 337560 451188 337572
rect 451240 337560 451246 337612
rect 451366 337560 451372 337612
rect 451424 337600 451430 337612
rect 452470 337600 452476 337612
rect 451424 337572 452476 337600
rect 451424 337560 451430 337572
rect 452470 337560 452476 337572
rect 452528 337560 452534 337612
rect 453298 337560 453304 337612
rect 453356 337600 453362 337612
rect 453942 337600 453948 337612
rect 453356 337572 453948 337600
rect 453356 337560 453362 337572
rect 453942 337560 453948 337572
rect 454000 337560 454006 337612
rect 456981 337603 457039 337609
rect 456981 337569 456993 337603
rect 457027 337600 457039 337603
rect 459097 337603 459155 337609
rect 457027 337572 458220 337600
rect 457027 337569 457039 337572
rect 456981 337563 457039 337569
rect 446401 337535 446459 337541
rect 446401 337532 446413 337535
rect 440292 337504 441660 337532
rect 441724 337504 442396 337532
rect 442460 337504 446413 337532
rect 440292 337492 440298 337504
rect 422941 337467 422999 337473
rect 422941 337433 422953 337467
rect 422987 337464 422999 337467
rect 433978 337464 433984 337476
rect 422987 337436 433984 337464
rect 422987 337433 422999 337436
rect 422941 337427 422999 337433
rect 433978 337424 433984 337436
rect 434036 337424 434042 337476
rect 434254 337424 434260 337476
rect 434312 337464 434318 337476
rect 439590 337464 439596 337476
rect 434312 337436 439596 337464
rect 434312 337424 434318 337436
rect 439590 337424 439596 337436
rect 439648 337424 439654 337476
rect 441632 337464 441660 337504
rect 442460 337464 442488 337504
rect 446401 337501 446413 337504
rect 446447 337501 446459 337535
rect 446401 337495 446459 337501
rect 447502 337492 447508 337544
rect 447560 337532 447566 337544
rect 448422 337532 448428 337544
rect 447560 337504 448428 337532
rect 447560 337492 447566 337504
rect 448422 337492 448428 337504
rect 448480 337492 448486 337544
rect 448517 337535 448575 337541
rect 448517 337501 448529 337535
rect 448563 337532 448575 337535
rect 456061 337535 456119 337541
rect 456061 337532 456073 337535
rect 448563 337504 456073 337532
rect 448563 337501 448575 337504
rect 448517 337495 448575 337501
rect 456061 337501 456073 337504
rect 456107 337501 456119 337535
rect 456061 337495 456119 337501
rect 456794 337492 456800 337544
rect 456852 337532 456858 337544
rect 458082 337532 458088 337544
rect 456852 337504 458088 337532
rect 456852 337492 456858 337504
rect 458082 337492 458088 337504
rect 458140 337492 458146 337544
rect 458192 337532 458220 337572
rect 459097 337569 459109 337603
rect 459143 337600 459155 337603
rect 520918 337600 520924 337612
rect 459143 337572 520924 337600
rect 459143 337569 459155 337572
rect 459097 337563 459155 337569
rect 520918 337560 520924 337572
rect 520976 337560 520982 337612
rect 460385 337535 460443 337541
rect 460385 337532 460397 337535
rect 458192 337504 460397 337532
rect 460385 337501 460397 337504
rect 460431 337501 460443 337535
rect 460385 337495 460443 337501
rect 461397 337535 461455 337541
rect 461397 337501 461409 337535
rect 461443 337532 461455 337535
rect 516778 337532 516784 337544
rect 461443 337504 516784 337532
rect 461443 337501 461455 337504
rect 461397 337495 461455 337501
rect 516778 337492 516784 337504
rect 516836 337492 516842 337544
rect 441632 337436 442488 337464
rect 443086 337424 443092 337476
rect 443144 337464 443150 337476
rect 514018 337464 514024 337476
rect 443144 337436 514024 337464
rect 443144 337424 443150 337436
rect 514018 337424 514024 337436
rect 514076 337424 514082 337476
rect 426434 337396 426440 337408
rect 422312 337368 426440 337396
rect 426434 337356 426440 337368
rect 426492 337356 426498 337408
rect 429838 337356 429844 337408
rect 429896 337396 429902 337408
rect 436741 337399 436799 337405
rect 436741 337396 436753 337399
rect 429896 337368 436753 337396
rect 429896 337356 429902 337368
rect 436741 337365 436753 337368
rect 436787 337365 436799 337399
rect 436741 337359 436799 337365
rect 449161 337399 449219 337405
rect 449161 337365 449173 337399
rect 449207 337396 449219 337399
rect 451369 337399 451427 337405
rect 451369 337396 451381 337399
rect 449207 337368 451381 337396
rect 449207 337365 449219 337368
rect 449161 337359 449219 337365
rect 451369 337365 451381 337368
rect 451415 337365 451427 337399
rect 451369 337359 451427 337365
rect 456061 337399 456119 337405
rect 456061 337365 456073 337399
rect 456107 337396 456119 337399
rect 470781 337399 470839 337405
rect 470781 337396 470793 337399
rect 456107 337368 470793 337396
rect 456107 337365 456119 337368
rect 456061 337359 456119 337365
rect 470781 337365 470793 337368
rect 470827 337365 470839 337399
rect 470781 337359 470839 337365
rect 480901 337399 480959 337405
rect 480901 337365 480913 337399
rect 480947 337396 480959 337399
rect 489917 337399 489975 337405
rect 489917 337396 489929 337399
rect 480947 337368 489929 337396
rect 480947 337365 480959 337368
rect 480901 337359 480959 337365
rect 489917 337365 489929 337368
rect 489963 337365 489975 337399
rect 489917 337359 489975 337365
rect 500221 337399 500279 337405
rect 500221 337365 500233 337399
rect 500267 337396 500279 337399
rect 509234 337396 509240 337408
rect 500267 337368 509240 337396
rect 500267 337365 500279 337368
rect 500221 337359 500279 337365
rect 509234 337356 509240 337368
rect 509292 337356 509298 337408
rect 366910 337288 366916 337340
rect 366968 337328 366974 337340
rect 380342 337328 380348 337340
rect 366968 337300 380348 337328
rect 366968 337288 366974 337300
rect 380342 337288 380348 337300
rect 380400 337288 380406 337340
rect 398466 337288 398472 337340
rect 398524 337328 398530 337340
rect 408770 337328 408776 337340
rect 398524 337300 408776 337328
rect 398524 337288 398530 337300
rect 408770 337288 408776 337300
rect 408828 337288 408834 337340
rect 409230 337288 409236 337340
rect 409288 337328 409294 337340
rect 409288 337300 417464 337328
rect 409288 337288 409294 337300
rect 372982 337260 372988 337272
rect 364536 337232 372988 337260
rect 372982 337220 372988 337232
rect 373040 337220 373046 337272
rect 417436 337260 417464 337300
rect 421006 337288 421012 337340
rect 421064 337328 421070 337340
rect 456981 337331 457039 337337
rect 456981 337328 456993 337331
rect 421064 337300 456993 337328
rect 421064 337288 421070 337300
rect 456981 337297 456993 337300
rect 457027 337297 457039 337331
rect 461581 337331 461639 337337
rect 461581 337328 461593 337331
rect 456981 337291 457039 337297
rect 457088 337300 461593 337328
rect 422941 337263 422999 337269
rect 422941 337260 422953 337263
rect 417436 337232 422953 337260
rect 422941 337229 422953 337232
rect 422987 337229 422999 337263
rect 422941 337223 422999 337229
rect 423490 337220 423496 337272
rect 423548 337260 423554 337272
rect 457088 337260 457116 337300
rect 461581 337297 461593 337300
rect 461627 337297 461639 337331
rect 463878 337328 463884 337340
rect 461581 337291 461639 337297
rect 461688 337300 463884 337328
rect 423548 337232 457116 337260
rect 457165 337263 457223 337269
rect 423548 337220 423554 337232
rect 457165 337229 457177 337263
rect 457211 337260 457223 337263
rect 460290 337260 460296 337272
rect 457211 337232 460296 337260
rect 457211 337229 457223 337232
rect 457165 337223 457223 337229
rect 460290 337220 460296 337232
rect 460348 337220 460354 337272
rect 460385 337263 460443 337269
rect 460385 337229 460397 337263
rect 460431 337260 460443 337263
rect 461688 337260 461716 337300
rect 463878 337288 463884 337300
rect 463936 337288 463942 337340
rect 465074 337288 465080 337340
rect 465132 337328 465138 337340
rect 466362 337328 466368 337340
rect 465132 337300 466368 337328
rect 465132 337288 465138 337300
rect 466362 337288 466368 337300
rect 466420 337288 466426 337340
rect 466457 337331 466515 337337
rect 466457 337297 466469 337331
rect 466503 337328 466515 337331
rect 470594 337328 470600 337340
rect 466503 337300 470600 337328
rect 466503 337297 466515 337300
rect 466457 337291 466515 337297
rect 470594 337288 470600 337300
rect 470652 337288 470658 337340
rect 470686 337288 470692 337340
rect 470744 337328 470750 337340
rect 529198 337328 529204 337340
rect 470744 337300 529204 337328
rect 470744 337288 470750 337300
rect 529198 337288 529204 337300
rect 529256 337288 529262 337340
rect 460431 337232 461716 337260
rect 460431 337229 460443 337232
rect 460385 337223 460443 337229
rect 463602 337220 463608 337272
rect 463660 337260 463666 337272
rect 469217 337263 469275 337269
rect 469217 337260 469229 337263
rect 463660 337232 469229 337260
rect 463660 337220 463666 337232
rect 469217 337229 469229 337232
rect 469263 337229 469275 337263
rect 469217 337223 469275 337229
rect 469490 337220 469496 337272
rect 469548 337260 469554 337272
rect 530578 337260 530584 337272
rect 469548 337232 530584 337260
rect 469548 337220 469554 337232
rect 530578 337220 530584 337232
rect 530636 337220 530642 337272
rect 314194 337192 314200 337204
rect 306208 337164 314200 337192
rect 314194 337152 314200 337164
rect 314252 337152 314258 337204
rect 321462 337152 321468 337204
rect 321520 337192 321526 337204
rect 326341 337195 326399 337201
rect 326341 337192 326353 337195
rect 321520 337164 326353 337192
rect 321520 337152 321526 337164
rect 326341 337161 326353 337164
rect 326387 337161 326399 337195
rect 342809 337195 342867 337201
rect 342809 337192 342821 337195
rect 326341 337155 326399 337161
rect 326448 337164 342821 337192
rect 312722 337124 312728 337136
rect 306116 337096 312728 337124
rect 312722 337084 312728 337096
rect 312780 337084 312786 337136
rect 316678 337084 316684 337136
rect 316736 337124 316742 337136
rect 326448 337124 326476 337164
rect 342809 337161 342821 337164
rect 342855 337161 342867 337195
rect 342809 337155 342867 337161
rect 342898 337152 342904 337204
rect 342956 337192 342962 337204
rect 345845 337195 345903 337201
rect 345845 337192 345857 337195
rect 342956 337164 345857 337192
rect 342956 337152 342962 337164
rect 345845 337161 345857 337164
rect 345891 337161 345903 337195
rect 345845 337155 345903 337161
rect 355962 337152 355968 337204
rect 356020 337192 356026 337204
rect 364981 337195 365039 337201
rect 364981 337192 364993 337195
rect 356020 337164 364993 337192
rect 356020 337152 356026 337164
rect 364981 337161 364993 337164
rect 365027 337161 365039 337195
rect 364981 337155 365039 337161
rect 369857 337195 369915 337201
rect 369857 337161 369869 337195
rect 369903 337192 369915 337195
rect 374641 337195 374699 337201
rect 374641 337192 374653 337195
rect 369903 337164 374653 337192
rect 369903 337161 369915 337164
rect 369857 337155 369915 337161
rect 374641 337161 374653 337164
rect 374687 337161 374699 337195
rect 374641 337155 374699 337161
rect 401870 337152 401876 337204
rect 401928 337192 401934 337204
rect 416958 337192 416964 337204
rect 401928 337164 416964 337192
rect 401928 337152 401934 337164
rect 416958 337152 416964 337164
rect 417016 337152 417022 337204
rect 423950 337152 423956 337204
rect 424008 337192 424014 337204
rect 427909 337195 427967 337201
rect 427909 337192 427921 337195
rect 424008 337164 427921 337192
rect 424008 337152 424014 337164
rect 427909 337161 427921 337164
rect 427955 337161 427967 337195
rect 427909 337155 427967 337161
rect 432782 337152 432788 337204
rect 432840 337192 432846 337204
rect 492674 337192 492680 337204
rect 432840 337164 492680 337192
rect 432840 337152 432846 337164
rect 492674 337152 492680 337164
rect 492732 337152 492738 337204
rect 509234 337152 509240 337204
rect 509292 337192 509298 337204
rect 510614 337192 510620 337204
rect 509292 337164 510620 337192
rect 509292 337152 509298 337164
rect 510614 337152 510620 337164
rect 510672 337152 510678 337204
rect 316736 337096 326476 337124
rect 316736 337084 316742 337096
rect 335262 337084 335268 337136
rect 335320 337124 335326 337136
rect 340785 337127 340843 337133
rect 335320 337096 340736 337124
rect 335320 337084 335326 337096
rect 95878 337016 95884 337068
rect 95936 337056 95942 337068
rect 265250 337056 265256 337068
rect 95936 337028 265256 337056
rect 95936 337016 95942 337028
rect 265250 337016 265256 337028
rect 265308 337016 265314 337068
rect 335817 337059 335875 337065
rect 335817 337025 335829 337059
rect 335863 337056 335875 337059
rect 340601 337059 340659 337065
rect 340601 337056 340613 337059
rect 335863 337028 340613 337056
rect 335863 337025 335875 337028
rect 335817 337019 335875 337025
rect 340601 337025 340613 337028
rect 340647 337025 340659 337059
rect 340708 337056 340736 337096
rect 340785 337093 340797 337127
rect 340831 337124 340843 337127
rect 366634 337124 366640 337136
rect 340831 337096 366640 337124
rect 340831 337093 340843 337096
rect 340785 337087 340843 337093
rect 366634 337084 366640 337096
rect 366692 337084 366698 337136
rect 369118 337084 369124 337136
rect 369176 337124 369182 337136
rect 371050 337124 371056 337136
rect 369176 337096 371056 337124
rect 369176 337084 369182 337096
rect 371050 337084 371056 337096
rect 371108 337084 371114 337136
rect 415118 337084 415124 337136
rect 415176 337124 415182 337136
rect 421558 337124 421564 337136
rect 415176 337096 421564 337124
rect 415176 337084 415182 337096
rect 421558 337084 421564 337096
rect 421616 337084 421622 337136
rect 433518 337124 433524 337136
rect 422956 337096 433524 337124
rect 367646 337056 367652 337068
rect 340708 337028 367652 337056
rect 340601 337019 340659 337025
rect 367646 337016 367652 337028
rect 367704 337016 367710 337068
rect 393590 337016 393596 337068
rect 393648 337056 393654 337068
rect 397454 337056 397460 337068
rect 393648 337028 397460 337056
rect 393648 337016 393654 337028
rect 397454 337016 397460 337028
rect 397512 337016 397518 337068
rect 103425 336991 103483 336997
rect 103425 336988 103437 336991
rect 93872 336960 103437 336988
rect 86957 336951 87015 336957
rect 103425 336957 103437 336960
rect 103471 336957 103483 336991
rect 103425 336951 103483 336957
rect 107562 336948 107568 337000
rect 107620 336988 107626 337000
rect 274082 336988 274088 337000
rect 107620 336960 274088 336988
rect 107620 336948 107626 336960
rect 274082 336948 274088 336960
rect 274140 336948 274146 337000
rect 319438 336948 319444 337000
rect 319496 336988 319502 337000
rect 345845 336991 345903 336997
rect 319496 336960 345704 336988
rect 319496 336948 319502 336960
rect 102778 336880 102784 336932
rect 102836 336920 102842 336932
rect 268194 336920 268200 336932
rect 102836 336892 268200 336920
rect 102836 336880 102842 336892
rect 268194 336880 268200 336892
rect 268252 336880 268258 336932
rect 333238 336880 333244 336932
rect 333296 336920 333302 336932
rect 336185 336923 336243 336929
rect 336185 336920 336197 336923
rect 333296 336892 336197 336920
rect 333296 336880 333302 336892
rect 336185 336889 336197 336892
rect 336231 336889 336243 336923
rect 336185 336883 336243 336889
rect 338758 336880 338764 336932
rect 338816 336920 338822 336932
rect 338816 336892 340736 336920
rect 338816 336880 338822 336892
rect 118602 336812 118608 336864
rect 118660 336852 118666 336864
rect 278498 336852 278504 336864
rect 118660 336824 278504 336852
rect 118660 336812 118666 336824
rect 278498 336812 278504 336824
rect 278556 336812 278562 336864
rect 327718 336812 327724 336864
rect 327776 336852 327782 336864
rect 340708 336852 340736 336892
rect 340782 336880 340788 336932
rect 340840 336920 340846 336932
rect 345569 336923 345627 336929
rect 345569 336920 345581 336923
rect 340840 336892 345581 336920
rect 340840 336880 340846 336892
rect 345569 336889 345581 336892
rect 345615 336889 345627 336923
rect 345569 336883 345627 336889
rect 340877 336855 340935 336861
rect 340877 336852 340889 336855
rect 327776 336824 340552 336852
rect 340708 336824 340889 336852
rect 327776 336812 327782 336824
rect 113177 336787 113235 336793
rect 113177 336753 113189 336787
rect 113223 336784 113235 336787
rect 122745 336787 122803 336793
rect 122745 336784 122757 336787
rect 113223 336756 122757 336784
rect 113223 336753 113235 336756
rect 113177 336747 113235 336753
rect 122745 336753 122757 336756
rect 122791 336753 122803 336787
rect 122745 336747 122803 336753
rect 125502 336744 125508 336796
rect 125560 336784 125566 336796
rect 281166 336784 281172 336796
rect 125560 336756 281172 336784
rect 125560 336744 125566 336756
rect 281166 336744 281172 336756
rect 281224 336744 281230 336796
rect 334713 336787 334771 336793
rect 334713 336753 334725 336787
rect 334759 336784 334771 336787
rect 340230 336784 340236 336796
rect 334759 336756 340236 336784
rect 334759 336753 334771 336756
rect 334713 336747 334771 336753
rect 340230 336744 340236 336756
rect 340288 336744 340294 336796
rect 249058 336676 249064 336728
rect 249116 336716 249122 336728
rect 250530 336716 250536 336728
rect 249116 336688 250536 336716
rect 249116 336676 249122 336688
rect 250530 336676 250536 336688
rect 250588 336676 250594 336728
rect 251818 336676 251824 336728
rect 251876 336716 251882 336728
rect 256418 336716 256424 336728
rect 251876 336688 256424 336716
rect 251876 336676 251882 336688
rect 256418 336676 256424 336688
rect 256476 336676 256482 336728
rect 262858 336676 262864 336728
rect 262916 336716 262922 336728
rect 263042 336716 263048 336728
rect 262916 336688 263048 336716
rect 262916 336676 262922 336688
rect 263042 336676 263048 336688
rect 263100 336676 263106 336728
rect 284386 336716 284392 336728
rect 284347 336688 284392 336716
rect 284386 336676 284392 336688
rect 284444 336676 284450 336728
rect 288805 336719 288863 336725
rect 288805 336685 288817 336719
rect 288851 336716 288863 336719
rect 288986 336716 288992 336728
rect 288851 336688 288992 336716
rect 288851 336685 288863 336688
rect 288805 336679 288863 336685
rect 288986 336676 288992 336688
rect 289044 336676 289050 336728
rect 327261 336719 327319 336725
rect 327261 336685 327273 336719
rect 327307 336716 327319 336719
rect 327626 336716 327632 336728
rect 327307 336688 327632 336716
rect 327307 336685 327319 336688
rect 327261 336679 327319 336685
rect 327626 336676 327632 336688
rect 327684 336676 327690 336728
rect 337378 336716 337384 336728
rect 337339 336688 337384 336716
rect 337378 336676 337384 336688
rect 337436 336676 337442 336728
rect 339773 336719 339831 336725
rect 339773 336685 339785 336719
rect 339819 336716 339831 336719
rect 340322 336716 340328 336728
rect 339819 336688 340328 336716
rect 339819 336685 339831 336688
rect 339773 336679 339831 336685
rect 340322 336676 340328 336688
rect 340380 336676 340386 336728
rect 340524 336580 340552 336824
rect 340877 336821 340889 336824
rect 340923 336821 340935 336855
rect 340877 336815 340935 336821
rect 341076 336824 343220 336852
rect 340785 336787 340843 336793
rect 340785 336753 340797 336787
rect 340831 336784 340843 336787
rect 340969 336787 341027 336793
rect 340969 336784 340981 336787
rect 340831 336756 340981 336784
rect 340831 336753 340843 336756
rect 340785 336747 340843 336753
rect 340969 336753 340981 336756
rect 341015 336753 341027 336787
rect 340969 336747 341027 336753
rect 341076 336580 341104 336824
rect 341153 336787 341211 336793
rect 341153 336753 341165 336787
rect 341199 336784 341211 336787
rect 343082 336784 343088 336796
rect 341199 336756 343088 336784
rect 341199 336753 341211 336756
rect 341153 336747 341211 336753
rect 343082 336744 343088 336756
rect 343140 336744 343146 336796
rect 343192 336784 343220 336824
rect 344370 336812 344376 336864
rect 344428 336852 344434 336864
rect 345477 336855 345535 336861
rect 345477 336852 345489 336855
rect 344428 336824 345489 336852
rect 344428 336812 344434 336824
rect 345477 336821 345489 336824
rect 345523 336821 345535 336855
rect 345477 336815 345535 336821
rect 345566 336784 345572 336796
rect 343192 336756 345572 336784
rect 345566 336744 345572 336756
rect 345624 336744 345630 336796
rect 345676 336784 345704 336960
rect 345845 336957 345857 336991
rect 345891 336988 345903 336991
rect 353386 336988 353392 337000
rect 345891 336960 353392 336988
rect 345891 336957 345903 336960
rect 345845 336951 345903 336957
rect 353386 336948 353392 336960
rect 353444 336948 353450 337000
rect 354033 336991 354091 336997
rect 354033 336957 354045 336991
rect 354079 336988 354091 336991
rect 369578 336988 369584 337000
rect 354079 336960 369584 336988
rect 354079 336957 354091 336960
rect 354033 336951 354091 336957
rect 369578 336948 369584 336960
rect 369636 336948 369642 337000
rect 378042 336948 378048 337000
rect 378100 336988 378106 337000
rect 385218 336988 385224 337000
rect 378100 336960 385224 336988
rect 378100 336948 378106 336960
rect 385218 336948 385224 336960
rect 385276 336948 385282 337000
rect 412726 336948 412732 337000
rect 412784 336988 412790 337000
rect 413830 336988 413836 337000
rect 412784 336960 413836 336988
rect 412784 336948 412790 336960
rect 413830 336948 413836 336960
rect 413888 336948 413894 337000
rect 345934 336880 345940 336932
rect 345992 336920 345998 336932
rect 360286 336920 360292 336932
rect 345992 336892 360292 336920
rect 345992 336880 345998 336892
rect 360286 336880 360292 336892
rect 360344 336880 360350 336932
rect 380802 336880 380808 336932
rect 380860 336920 380866 336932
rect 386230 336920 386236 336932
rect 380860 336892 386236 336920
rect 380860 336880 380866 336892
rect 386230 336880 386236 336892
rect 386288 336880 386294 336932
rect 392118 336880 392124 336932
rect 392176 336920 392182 336932
rect 393590 336920 393596 336932
rect 392176 336892 393596 336920
rect 392176 336880 392182 336892
rect 393590 336880 393596 336892
rect 393648 336880 393654 336932
rect 401410 336880 401416 336932
rect 401468 336920 401474 336932
rect 404998 336920 405004 336932
rect 401468 336892 405004 336920
rect 401468 336880 401474 336892
rect 404998 336880 405004 336892
rect 405056 336880 405062 336932
rect 409046 336880 409052 336932
rect 409104 336920 409110 336932
rect 422956 336920 422984 337096
rect 433518 337084 433524 337096
rect 433576 337084 433582 337136
rect 436741 337127 436799 337133
rect 436741 337093 436753 337127
rect 436787 337124 436799 337127
rect 485774 337124 485780 337136
rect 436787 337096 485780 337124
rect 436787 337093 436799 337096
rect 436741 337087 436799 337093
rect 485774 337084 485780 337096
rect 485832 337084 485838 337136
rect 489917 337127 489975 337133
rect 489917 337093 489929 337127
rect 489963 337124 489975 337127
rect 500221 337127 500279 337133
rect 500221 337124 500233 337127
rect 489963 337096 500233 337124
rect 489963 337093 489975 337096
rect 489917 337087 489975 337093
rect 500221 337093 500233 337096
rect 500267 337093 500279 337127
rect 500221 337087 500279 337093
rect 426894 337016 426900 337068
rect 426952 337056 426958 337068
rect 477586 337056 477592 337068
rect 426952 337028 477592 337056
rect 426952 337016 426958 337028
rect 477586 337016 477592 337028
rect 477644 337016 477650 337068
rect 432233 336991 432291 336997
rect 432233 336957 432245 336991
rect 432279 336988 432291 336991
rect 475378 336988 475384 337000
rect 432279 336960 475384 336988
rect 432279 336957 432291 336960
rect 432233 336951 432291 336957
rect 475378 336948 475384 336960
rect 475436 336948 475442 337000
rect 409104 336892 422984 336920
rect 427909 336923 427967 336929
rect 409104 336880 409110 336892
rect 427909 336889 427921 336923
rect 427955 336920 427967 336923
rect 466457 336923 466515 336929
rect 466457 336920 466469 336923
rect 427955 336892 466469 336920
rect 427955 336889 427967 336892
rect 427909 336883 427967 336889
rect 466457 336889 466469 336892
rect 466503 336889 466515 336923
rect 466457 336883 466515 336889
rect 466546 336880 466552 336932
rect 466604 336920 466610 336932
rect 470502 336920 470508 336932
rect 466604 336892 470508 336920
rect 466604 336880 466610 336892
rect 470502 336880 470508 336892
rect 470560 336880 470566 336932
rect 470781 336923 470839 336929
rect 470781 336889 470793 336923
rect 470827 336920 470839 336923
rect 480901 336923 480959 336929
rect 480901 336920 480913 336923
rect 470827 336892 480913 336920
rect 470827 336889 470839 336892
rect 470781 336883 470839 336889
rect 480901 336889 480913 336892
rect 480947 336889 480959 336923
rect 480901 336883 480959 336889
rect 345753 336855 345811 336861
rect 345753 336821 345765 336855
rect 345799 336852 345811 336855
rect 357342 336852 357348 336864
rect 345799 336824 357348 336852
rect 345799 336821 345811 336824
rect 345753 336815 345811 336821
rect 357342 336812 357348 336824
rect 357400 336812 357406 336864
rect 362218 336812 362224 336864
rect 362276 336852 362282 336864
rect 365162 336852 365168 336864
rect 362276 336824 365168 336852
rect 362276 336812 362282 336824
rect 365162 336812 365168 336824
rect 365220 336812 365226 336864
rect 381630 336812 381636 336864
rect 381688 336852 381694 336864
rect 384758 336852 384764 336864
rect 381688 336824 384764 336852
rect 381688 336812 381694 336824
rect 384758 336812 384764 336824
rect 384816 336812 384822 336864
rect 396074 336812 396080 336864
rect 396132 336852 396138 336864
rect 398098 336852 398104 336864
rect 396132 336824 398104 336852
rect 396132 336812 396138 336824
rect 398098 336812 398104 336824
rect 398156 336812 398162 336864
rect 419994 336812 420000 336864
rect 420052 336852 420058 336864
rect 420730 336852 420736 336864
rect 420052 336824 420736 336852
rect 420052 336812 420058 336824
rect 420730 336812 420736 336824
rect 420788 336812 420794 336864
rect 424962 336812 424968 336864
rect 425020 336852 425026 336864
rect 439498 336852 439504 336864
rect 425020 336824 439504 336852
rect 425020 336812 425026 336824
rect 439498 336812 439504 336824
rect 439556 336812 439562 336864
rect 441617 336855 441675 336861
rect 441617 336821 441629 336855
rect 441663 336852 441675 336855
rect 451093 336855 451151 336861
rect 451093 336852 451105 336855
rect 441663 336824 451105 336852
rect 441663 336821 441675 336824
rect 441617 336815 441675 336821
rect 451093 336821 451105 336824
rect 451139 336821 451151 336855
rect 451093 336815 451151 336821
rect 451826 336812 451832 336864
rect 451884 336852 451890 336864
rect 459097 336855 459155 336861
rect 459097 336852 459109 336855
rect 451884 336824 459109 336852
rect 451884 336812 451890 336824
rect 459097 336821 459109 336824
rect 459143 336821 459155 336855
rect 459097 336815 459155 336821
rect 459186 336812 459192 336864
rect 459244 336852 459250 336864
rect 460198 336852 460204 336864
rect 459244 336824 460204 336852
rect 459244 336812 459250 336824
rect 460198 336812 460204 336824
rect 460256 336812 460262 336864
rect 460382 336812 460388 336864
rect 460440 336852 460446 336864
rect 460750 336852 460756 336864
rect 460440 336824 460756 336852
rect 460440 336812 460446 336824
rect 460750 336812 460756 336824
rect 460808 336812 460814 336864
rect 461581 336855 461639 336861
rect 461581 336821 461593 336855
rect 461627 336852 461639 336855
rect 469214 336852 469220 336864
rect 461627 336824 469220 336852
rect 461627 336821 461639 336824
rect 461581 336815 461639 336821
rect 469214 336812 469220 336824
rect 469272 336812 469278 336864
rect 509878 336852 509884 336864
rect 469324 336824 509884 336852
rect 351454 336784 351460 336796
rect 345676 336756 351460 336784
rect 351454 336744 351460 336756
rect 351512 336744 351518 336796
rect 352558 336744 352564 336796
rect 352616 336784 352622 336796
rect 357802 336784 357808 336796
rect 352616 336756 357808 336784
rect 352616 336744 352622 336756
rect 357802 336744 357808 336756
rect 357860 336744 357866 336796
rect 363598 336744 363604 336796
rect 363656 336784 363662 336796
rect 364702 336784 364708 336796
rect 363656 336756 364708 336784
rect 363656 336744 363662 336756
rect 364702 336744 364708 336756
rect 364760 336744 364766 336796
rect 370498 336744 370504 336796
rect 370556 336784 370562 336796
rect 372522 336784 372528 336796
rect 370556 336756 372528 336784
rect 370556 336744 370562 336756
rect 372522 336744 372528 336756
rect 372580 336744 372586 336796
rect 376018 336744 376024 336796
rect 376076 336784 376082 336796
rect 376938 336784 376944 336796
rect 376076 336756 376944 336784
rect 376076 336744 376082 336756
rect 376938 336744 376944 336756
rect 376996 336744 377002 336796
rect 377674 336744 377680 336796
rect 377732 336784 377738 336796
rect 378410 336784 378416 336796
rect 377732 336756 378416 336784
rect 377732 336744 377738 336756
rect 378410 336744 378416 336756
rect 378468 336744 378474 336796
rect 395062 336744 395068 336796
rect 395120 336784 395126 336796
rect 395982 336784 395988 336796
rect 395120 336756 395988 336784
rect 395120 336744 395126 336756
rect 395982 336744 395988 336756
rect 396040 336744 396046 336796
rect 396534 336744 396540 336796
rect 396592 336784 396598 336796
rect 398190 336784 398196 336796
rect 396592 336756 398196 336784
rect 396592 336744 396598 336756
rect 398190 336744 398196 336756
rect 398248 336744 398254 336796
rect 418522 336744 418528 336796
rect 418580 336784 418586 336796
rect 419442 336784 419448 336796
rect 418580 336756 419448 336784
rect 418580 336744 418586 336756
rect 419442 336744 419448 336756
rect 419500 336744 419506 336796
rect 419534 336744 419540 336796
rect 419592 336784 419598 336796
rect 420822 336784 420828 336796
rect 419592 336756 420828 336784
rect 419592 336744 419598 336756
rect 420822 336744 420828 336756
rect 420880 336744 420886 336796
rect 421466 336744 421472 336796
rect 421524 336784 421530 336796
rect 422202 336784 422208 336796
rect 421524 336756 422208 336784
rect 421524 336744 421530 336756
rect 422202 336744 422208 336756
rect 422260 336744 422266 336796
rect 422478 336744 422484 336796
rect 422536 336784 422542 336796
rect 424318 336784 424324 336796
rect 422536 336756 424324 336784
rect 422536 336744 422542 336756
rect 424318 336744 424324 336756
rect 424376 336744 424382 336796
rect 424410 336744 424416 336796
rect 424468 336784 424474 336796
rect 451277 336787 451335 336793
rect 424468 336756 425008 336784
rect 424468 336744 424474 336756
rect 424980 336728 425008 336756
rect 451277 336753 451289 336787
rect 451323 336784 451335 336787
rect 457165 336787 457223 336793
rect 457165 336784 457177 336787
rect 451323 336756 457177 336784
rect 451323 336753 451335 336756
rect 451277 336747 451335 336753
rect 457165 336753 457177 336756
rect 457211 336753 457223 336787
rect 457165 336747 457223 336753
rect 457254 336744 457260 336796
rect 457312 336784 457318 336796
rect 457990 336784 457996 336796
rect 457312 336756 457996 336784
rect 457312 336744 457318 336756
rect 457990 336744 457996 336756
rect 458048 336744 458054 336796
rect 458266 336744 458272 336796
rect 458324 336784 458330 336796
rect 459462 336784 459468 336796
rect 458324 336756 459468 336784
rect 458324 336744 458330 336756
rect 459462 336744 459468 336756
rect 459520 336744 459526 336796
rect 459738 336744 459744 336796
rect 459796 336784 459802 336796
rect 460842 336784 460848 336796
rect 459796 336756 460848 336784
rect 459796 336744 459802 336756
rect 460842 336744 460848 336756
rect 460900 336744 460906 336796
rect 461210 336744 461216 336796
rect 461268 336784 461274 336796
rect 462130 336784 462136 336796
rect 461268 336756 462136 336784
rect 461268 336744 461274 336756
rect 462130 336744 462136 336756
rect 462188 336744 462194 336796
rect 462682 336744 462688 336796
rect 462740 336784 462746 336796
rect 463510 336784 463516 336796
rect 462740 336756 463516 336784
rect 462740 336744 462746 336756
rect 463510 336744 463516 336756
rect 463568 336744 463574 336796
rect 464154 336744 464160 336796
rect 464212 336784 464218 336796
rect 464982 336784 464988 336796
rect 464212 336756 464988 336784
rect 464212 336744 464218 336756
rect 464982 336744 464988 336756
rect 465040 336744 465046 336796
rect 465074 336744 465080 336796
rect 465132 336784 465138 336796
rect 469324 336784 469352 336824
rect 509878 336812 509884 336824
rect 509936 336812 509942 336864
rect 505738 336784 505744 336796
rect 465132 336756 469352 336784
rect 469416 336756 505744 336784
rect 465132 336744 465138 336756
rect 424962 336676 424968 336728
rect 425020 336676 425026 336728
rect 466273 336719 466331 336725
rect 466273 336685 466285 336719
rect 466319 336716 466331 336719
rect 469416 336716 469444 336756
rect 505738 336744 505744 336756
rect 505796 336744 505802 336796
rect 466319 336688 469444 336716
rect 466319 336685 466331 336688
rect 466273 336679 466331 336685
rect 340524 336552 341104 336580
rect 247218 336404 247224 336456
rect 247276 336444 247282 336456
rect 248138 336444 248144 336456
rect 247276 336416 248144 336444
rect 247276 336404 247282 336416
rect 248138 336404 248144 336416
rect 248196 336404 248202 336456
rect 251450 335792 251456 335844
rect 251508 335832 251514 335844
rect 252462 335832 252468 335844
rect 251508 335804 252468 335832
rect 251508 335792 251514 335804
rect 252462 335792 252468 335804
rect 252520 335792 252526 335844
rect 236178 335656 236184 335708
rect 236236 335696 236242 335708
rect 237006 335696 237012 335708
rect 236236 335668 237012 335696
rect 236236 335656 236242 335668
rect 237006 335656 237012 335668
rect 237064 335656 237070 335708
rect 302234 335656 302240 335708
rect 302292 335696 302298 335708
rect 302694 335696 302700 335708
rect 302292 335668 302700 335696
rect 302292 335656 302298 335668
rect 302694 335656 302700 335668
rect 302752 335656 302758 335708
rect 332686 335656 332692 335708
rect 332744 335696 332750 335708
rect 333422 335696 333428 335708
rect 332744 335668 333428 335696
rect 332744 335656 332750 335668
rect 333422 335656 333428 335668
rect 333480 335656 333486 335708
rect 334066 335656 334072 335708
rect 334124 335696 334130 335708
rect 334894 335696 334900 335708
rect 334124 335668 334900 335696
rect 334124 335656 334130 335668
rect 334894 335656 334900 335668
rect 334952 335656 334958 335708
rect 390646 335656 390652 335708
rect 390704 335656 390710 335708
rect 236086 335588 236092 335640
rect 236144 335628 236150 335640
rect 236546 335628 236552 335640
rect 236144 335600 236552 335628
rect 236144 335588 236150 335600
rect 236546 335588 236552 335600
rect 236604 335588 236610 335640
rect 241606 335588 241612 335640
rect 241664 335628 241670 335640
rect 242342 335628 242348 335640
rect 241664 335600 242348 335628
rect 241664 335588 241670 335600
rect 242342 335588 242348 335600
rect 242400 335588 242406 335640
rect 260926 335588 260932 335640
rect 260984 335628 260990 335640
rect 261478 335628 261484 335640
rect 260984 335600 261484 335628
rect 260984 335588 260990 335600
rect 261478 335588 261484 335600
rect 261536 335588 261542 335640
rect 263686 335588 263692 335640
rect 263744 335628 263750 335640
rect 264422 335628 264428 335640
rect 263744 335600 264428 335628
rect 263744 335588 263750 335600
rect 264422 335588 264428 335600
rect 264480 335588 264486 335640
rect 265066 335588 265072 335640
rect 265124 335628 265130 335640
rect 265894 335628 265900 335640
rect 265124 335600 265900 335628
rect 265124 335588 265130 335600
rect 265894 335588 265900 335600
rect 265952 335588 265958 335640
rect 266446 335588 266452 335640
rect 266504 335628 266510 335640
rect 267366 335628 267372 335640
rect 266504 335600 267372 335628
rect 266504 335588 266510 335600
rect 267366 335588 267372 335600
rect 267424 335588 267430 335640
rect 280246 335588 280252 335640
rect 280304 335628 280310 335640
rect 280614 335628 280620 335640
rect 280304 335600 280620 335628
rect 280304 335588 280310 335600
rect 280614 335588 280620 335600
rect 280672 335588 280678 335640
rect 281534 335588 281540 335640
rect 281592 335628 281598 335640
rect 282086 335628 282092 335640
rect 281592 335600 282092 335628
rect 281592 335588 281598 335600
rect 282086 335588 282092 335600
rect 282144 335588 282150 335640
rect 283006 335588 283012 335640
rect 283064 335628 283070 335640
rect 283558 335628 283564 335640
rect 283064 335600 283564 335628
rect 283064 335588 283070 335600
rect 283558 335588 283564 335600
rect 283616 335588 283622 335640
rect 285674 335588 285680 335640
rect 285732 335628 285738 335640
rect 285950 335628 285956 335640
rect 285732 335600 285956 335628
rect 285732 335588 285738 335600
rect 285950 335588 285956 335600
rect 286008 335588 286014 335640
rect 286042 335588 286048 335640
rect 286100 335628 286106 335640
rect 286594 335628 286600 335640
rect 286100 335600 286600 335628
rect 286100 335588 286106 335600
rect 286594 335588 286600 335600
rect 286652 335588 286658 335640
rect 287054 335588 287060 335640
rect 287112 335628 287118 335640
rect 287974 335628 287980 335640
rect 287112 335600 287980 335628
rect 287112 335588 287118 335600
rect 287974 335588 287980 335600
rect 288032 335588 288038 335640
rect 288434 335588 288440 335640
rect 288492 335628 288498 335640
rect 289446 335628 289452 335640
rect 288492 335600 289452 335628
rect 288492 335588 288498 335600
rect 289446 335588 289452 335600
rect 289504 335588 289510 335640
rect 292758 335588 292764 335640
rect 292816 335628 292822 335640
rect 293310 335628 293316 335640
rect 292816 335600 293316 335628
rect 292816 335588 292822 335600
rect 293310 335588 293316 335600
rect 293368 335588 293374 335640
rect 298278 335588 298284 335640
rect 298336 335628 298342 335640
rect 298646 335628 298652 335640
rect 298336 335600 298652 335628
rect 298336 335588 298342 335600
rect 298646 335588 298652 335600
rect 298704 335588 298710 335640
rect 300854 335588 300860 335640
rect 300912 335628 300918 335640
rect 301222 335628 301228 335640
rect 300912 335600 301228 335628
rect 300912 335588 300918 335600
rect 301222 335588 301228 335600
rect 301280 335588 301286 335640
rect 303614 335588 303620 335640
rect 303672 335628 303678 335640
rect 304166 335628 304172 335640
rect 303672 335600 304172 335628
rect 303672 335588 303678 335600
rect 304166 335588 304172 335600
rect 304224 335588 304230 335640
rect 304994 335588 305000 335640
rect 305052 335628 305058 335640
rect 305638 335628 305644 335640
rect 305052 335600 305644 335628
rect 305052 335588 305058 335600
rect 305638 335588 305644 335600
rect 305696 335588 305702 335640
rect 307754 335588 307760 335640
rect 307812 335628 307818 335640
rect 308582 335628 308588 335640
rect 307812 335600 308588 335628
rect 307812 335588 307818 335600
rect 308582 335588 308588 335600
rect 308640 335588 308646 335640
rect 309134 335588 309140 335640
rect 309192 335628 309198 335640
rect 310054 335628 310060 335640
rect 309192 335600 310060 335628
rect 309192 335588 309198 335600
rect 310054 335588 310060 335600
rect 310112 335588 310118 335640
rect 321646 335588 321652 335640
rect 321704 335628 321710 335640
rect 322198 335628 322204 335640
rect 321704 335600 322204 335628
rect 321704 335588 321710 335600
rect 322198 335588 322204 335600
rect 322256 335588 322262 335640
rect 329834 335588 329840 335640
rect 329892 335628 329898 335640
rect 330110 335628 330116 335640
rect 329892 335600 330116 335628
rect 329892 335588 329898 335600
rect 330110 335588 330116 335600
rect 330168 335588 330174 335640
rect 332594 335588 332600 335640
rect 332652 335628 332658 335640
rect 333054 335628 333060 335640
rect 332652 335600 333060 335628
rect 332652 335588 332658 335600
rect 333054 335588 333060 335600
rect 333112 335588 333118 335640
rect 333974 335588 333980 335640
rect 334032 335628 334038 335640
rect 334526 335628 334532 335640
rect 334032 335600 334532 335628
rect 334032 335588 334038 335600
rect 334526 335588 334532 335600
rect 334584 335588 334590 335640
rect 335354 335588 335360 335640
rect 335412 335628 335418 335640
rect 335998 335628 336004 335640
rect 335412 335600 336004 335628
rect 335412 335588 335418 335600
rect 335998 335588 336004 335600
rect 336056 335588 336062 335640
rect 338114 335588 338120 335640
rect 338172 335628 338178 335640
rect 338942 335628 338948 335640
rect 338172 335600 338948 335628
rect 338172 335588 338178 335600
rect 338942 335588 338948 335600
rect 339000 335588 339006 335640
rect 361666 335588 361672 335640
rect 361724 335628 361730 335640
rect 362310 335628 362316 335640
rect 361724 335600 362316 335628
rect 361724 335588 361730 335600
rect 362310 335588 362316 335600
rect 362368 335588 362374 335640
rect 363046 335588 363052 335640
rect 363104 335628 363110 335640
rect 363782 335628 363788 335640
rect 363104 335600 363788 335628
rect 363104 335588 363110 335600
rect 363782 335588 363788 335600
rect 363840 335588 363846 335640
rect 367278 335588 367284 335640
rect 367336 335628 367342 335640
rect 367922 335628 367928 335640
rect 367336 335600 367928 335628
rect 367336 335588 367342 335600
rect 367922 335588 367928 335600
rect 367980 335588 367986 335640
rect 372614 335588 372620 335640
rect 372672 335628 372678 335640
rect 373258 335628 373264 335640
rect 372672 335600 373264 335628
rect 372672 335588 372678 335600
rect 373258 335588 373264 335600
rect 373316 335588 373322 335640
rect 390664 335504 390692 335656
rect 390646 335452 390652 335504
rect 390704 335452 390710 335504
rect 265250 335288 265256 335300
rect 265211 335260 265256 335288
rect 265250 335248 265256 335260
rect 265308 335248 265314 335300
rect 284389 335223 284447 335229
rect 284389 335189 284401 335223
rect 284435 335220 284447 335223
rect 284478 335220 284484 335232
rect 284435 335192 284484 335220
rect 284435 335189 284447 335192
rect 284389 335183 284447 335189
rect 284478 335180 284484 335192
rect 284536 335180 284542 335232
rect 248506 334908 248512 334960
rect 248564 334948 248570 334960
rect 249518 334948 249524 334960
rect 248564 334920 249524 334948
rect 248564 334908 248570 334920
rect 249518 334908 249524 334920
rect 249576 334908 249582 334960
rect 278774 334772 278780 334824
rect 278832 334812 278838 334824
rect 278958 334812 278964 334824
rect 278832 334784 278964 334812
rect 278832 334772 278838 334784
rect 278958 334772 278964 334784
rect 279016 334772 279022 334824
rect 302602 334704 302608 334756
rect 302660 334744 302666 334756
rect 303062 334744 303068 334756
rect 302660 334716 303068 334744
rect 302660 334704 302666 334716
rect 303062 334704 303068 334716
rect 303120 334704 303126 334756
rect 258166 334568 258172 334620
rect 258224 334608 258230 334620
rect 258534 334608 258540 334620
rect 258224 334580 258540 334608
rect 258224 334568 258230 334580
rect 258534 334568 258540 334580
rect 258592 334568 258598 334620
rect 234982 334500 234988 334552
rect 235040 334540 235046 334552
rect 235626 334540 235632 334552
rect 235040 334512 235632 334540
rect 235040 334500 235046 334512
rect 235626 334500 235632 334512
rect 235684 334500 235690 334552
rect 336734 334500 336740 334552
rect 336792 334540 336798 334552
rect 336918 334540 336924 334552
rect 336792 334512 336924 334540
rect 336792 334500 336798 334512
rect 336918 334500 336924 334512
rect 336976 334500 336982 334552
rect 250165 334475 250223 334481
rect 250165 334441 250177 334475
rect 250211 334472 250223 334475
rect 250622 334472 250628 334484
rect 250211 334444 250628 334472
rect 250211 334441 250223 334444
rect 250165 334435 250223 334441
rect 250622 334432 250628 334444
rect 250680 334432 250686 334484
rect 270773 334339 270831 334345
rect 270773 334305 270785 334339
rect 270819 334336 270831 334339
rect 271230 334336 271236 334348
rect 270819 334308 271236 334336
rect 270819 334305 270831 334308
rect 270773 334299 270831 334305
rect 271230 334296 271236 334308
rect 271288 334296 271294 334348
rect 272245 334339 272303 334345
rect 272245 334305 272257 334339
rect 272291 334336 272303 334339
rect 272702 334336 272708 334348
rect 272291 334308 272708 334336
rect 272291 334305 272303 334308
rect 272245 334299 272303 334305
rect 272702 334296 272708 334308
rect 272760 334296 272766 334348
rect 247862 333956 247868 334008
rect 247920 333996 247926 334008
rect 248598 333996 248604 334008
rect 247920 333968 248604 333996
rect 247920 333956 247926 333968
rect 248598 333956 248604 333968
rect 248656 333956 248662 334008
rect 325970 333276 325976 333328
rect 326028 333316 326034 333328
rect 326522 333316 326528 333328
rect 326028 333288 326528 333316
rect 326028 333276 326034 333288
rect 326522 333276 326528 333288
rect 326580 333276 326586 333328
rect 374086 333140 374092 333192
rect 374144 333180 374150 333192
rect 374730 333180 374736 333192
rect 374144 333152 374736 333180
rect 374144 333140 374150 333152
rect 374730 333140 374736 333152
rect 374788 333140 374794 333192
rect 356146 332800 356152 332852
rect 356204 332840 356210 332852
rect 356606 332840 356612 332852
rect 356204 332812 356612 332840
rect 356204 332800 356210 332812
rect 356606 332800 356612 332812
rect 356664 332800 356670 332852
rect 284662 332528 284668 332580
rect 284720 332568 284726 332580
rect 285122 332568 285128 332580
rect 284720 332540 285128 332568
rect 284720 332528 284726 332540
rect 285122 332528 285128 332540
rect 285180 332528 285186 332580
rect 331214 332120 331220 332172
rect 331272 332160 331278 332172
rect 331490 332160 331496 332172
rect 331272 332132 331496 332160
rect 331272 332120 331278 332132
rect 331490 332120 331496 332132
rect 331548 332120 331554 332172
rect 242986 332052 242992 332104
rect 243044 332092 243050 332104
rect 243446 332092 243452 332104
rect 243044 332064 243452 332092
rect 243044 332052 243050 332064
rect 243446 332052 243452 332064
rect 243504 332052 243510 332104
rect 310514 332052 310520 332104
rect 310572 332092 310578 332104
rect 311526 332092 311532 332104
rect 310572 332064 311532 332092
rect 310572 332052 310578 332064
rect 311526 332052 311532 332064
rect 311584 332052 311590 332104
rect 331306 331712 331312 331764
rect 331364 331752 331370 331764
rect 331950 331752 331956 331764
rect 331364 331724 331956 331752
rect 331364 331712 331370 331724
rect 331950 331712 331956 331724
rect 332008 331712 332014 331764
rect 299566 331304 299572 331356
rect 299624 331304 299630 331356
rect 328546 331304 328552 331356
rect 328604 331344 328610 331356
rect 329006 331344 329012 331356
rect 328604 331316 329012 331344
rect 328604 331304 328610 331316
rect 329006 331304 329012 331316
rect 329064 331304 329070 331356
rect 259638 331168 259644 331220
rect 259696 331208 259702 331220
rect 259822 331208 259828 331220
rect 259696 331180 259828 331208
rect 259696 331168 259702 331180
rect 259822 331168 259828 331180
rect 259880 331168 259886 331220
rect 299584 331084 299612 331304
rect 336826 331236 336832 331288
rect 336884 331236 336890 331288
rect 336844 331152 336872 331236
rect 341150 331168 341156 331220
rect 341208 331208 341214 331220
rect 341334 331208 341340 331220
rect 341208 331180 341340 331208
rect 341208 331168 341214 331180
rect 341334 331168 341340 331180
rect 341392 331168 341398 331220
rect 360286 331168 360292 331220
rect 360344 331208 360350 331220
rect 360470 331208 360476 331220
rect 360344 331180 360476 331208
rect 360344 331168 360350 331180
rect 360470 331168 360476 331180
rect 360528 331168 360534 331220
rect 389266 331168 389272 331220
rect 389324 331208 389330 331220
rect 389450 331208 389456 331220
rect 389324 331180 389456 331208
rect 389324 331168 389330 331180
rect 389450 331168 389456 331180
rect 389508 331168 389514 331220
rect 336826 331100 336832 331152
rect 336884 331100 336890 331152
rect 299566 331032 299572 331084
rect 299624 331032 299630 331084
rect 306466 331032 306472 331084
rect 306524 331072 306530 331084
rect 306650 331072 306656 331084
rect 306524 331044 306656 331072
rect 306524 331032 306530 331044
rect 306650 331032 306656 331044
rect 306708 331032 306714 331084
rect 299474 330964 299480 331016
rect 299532 331004 299538 331016
rect 299658 331004 299664 331016
rect 299532 330976 299664 331004
rect 299532 330964 299538 330976
rect 299658 330964 299664 330976
rect 299716 330964 299722 331016
rect 301130 330488 301136 330540
rect 301188 330528 301194 330540
rect 301682 330528 301688 330540
rect 301188 330500 301688 330528
rect 301188 330488 301194 330500
rect 301682 330488 301688 330500
rect 301740 330488 301746 330540
rect 284294 329536 284300 329588
rect 284352 329576 284358 329588
rect 284570 329576 284576 329588
rect 284352 329548 284576 329576
rect 284352 329536 284358 329548
rect 284570 329536 284576 329548
rect 284628 329536 284634 329588
rect 270770 328488 270776 328500
rect 270731 328460 270776 328488
rect 270770 328448 270776 328460
rect 270828 328448 270834 328500
rect 272242 328488 272248 328500
rect 272203 328460 272248 328488
rect 272242 328448 272248 328460
rect 272300 328448 272306 328500
rect 278866 328448 278872 328500
rect 278924 328488 278930 328500
rect 279050 328488 279056 328500
rect 278924 328460 279056 328488
rect 278924 328448 278930 328460
rect 279050 328448 279056 328460
rect 279108 328448 279114 328500
rect 303890 328448 303896 328500
rect 303948 328488 303954 328500
rect 304626 328488 304632 328500
rect 303948 328460 304632 328488
rect 303948 328448 303954 328460
rect 304626 328448 304632 328460
rect 304684 328448 304690 328500
rect 323302 328448 323308 328500
rect 323360 328488 323366 328500
rect 323670 328488 323676 328500
rect 323360 328460 323676 328488
rect 323360 328448 323366 328460
rect 323670 328448 323676 328460
rect 323728 328448 323734 328500
rect 324682 328448 324688 328500
rect 324740 328488 324746 328500
rect 325142 328488 325148 328500
rect 324740 328460 325148 328488
rect 324740 328448 324746 328460
rect 325142 328448 325148 328460
rect 325200 328448 325206 328500
rect 330202 328448 330208 328500
rect 330260 328488 330266 328500
rect 330478 328488 330484 328500
rect 330260 328460 330484 328488
rect 330260 328448 330266 328460
rect 330478 328448 330484 328460
rect 330536 328448 330542 328500
rect 259822 328420 259828 328432
rect 259783 328392 259828 328420
rect 259822 328380 259828 328392
rect 259880 328380 259886 328432
rect 295518 328380 295524 328432
rect 295576 328420 295582 328432
rect 295702 328420 295708 328432
rect 295576 328392 295708 328420
rect 295576 328380 295582 328392
rect 295702 328380 295708 328392
rect 295760 328380 295766 328432
rect 296806 328380 296812 328432
rect 296864 328420 296870 328432
rect 296990 328420 296996 328432
rect 296864 328392 296996 328420
rect 296864 328380 296870 328392
rect 296990 328380 296996 328392
rect 297048 328380 297054 328432
rect 302602 328420 302608 328432
rect 302563 328392 302608 328420
rect 302602 328380 302608 328392
rect 302660 328380 302666 328432
rect 337378 328420 337384 328432
rect 337339 328392 337384 328420
rect 337378 328380 337384 328392
rect 337436 328380 337442 328432
rect 341334 328420 341340 328432
rect 341295 328392 341340 328420
rect 341334 328380 341340 328392
rect 341392 328380 341398 328432
rect 389450 328420 389456 328432
rect 389411 328392 389456 328420
rect 389450 328380 389456 328392
rect 389508 328380 389514 328432
rect 470594 328420 470600 328432
rect 470555 328392 470600 328420
rect 470594 328380 470600 328392
rect 470652 328380 470658 328432
rect 250162 327128 250168 327140
rect 250123 327100 250168 327128
rect 250162 327088 250168 327100
rect 250220 327088 250226 327140
rect 327258 327128 327264 327140
rect 327219 327100 327264 327128
rect 327258 327088 327264 327100
rect 327316 327088 327322 327140
rect 273533 327063 273591 327069
rect 273533 327029 273545 327063
rect 273579 327060 273591 327063
rect 273622 327060 273628 327072
rect 273579 327032 273628 327060
rect 273579 327029 273591 327032
rect 273533 327023 273591 327029
rect 273622 327020 273628 327032
rect 273680 327020 273686 327072
rect 284662 327020 284668 327072
rect 284720 327060 284726 327072
rect 284754 327060 284760 327072
rect 284720 327032 284760 327060
rect 284720 327020 284726 327032
rect 284754 327020 284760 327032
rect 284812 327020 284818 327072
rect 285953 327063 286011 327069
rect 285953 327029 285965 327063
rect 285999 327060 286011 327063
rect 286042 327060 286048 327072
rect 285999 327032 286048 327060
rect 285999 327029 286011 327032
rect 285953 327023 286011 327029
rect 286042 327020 286048 327032
rect 286100 327020 286106 327072
rect 330110 327060 330116 327072
rect 330071 327032 330116 327060
rect 330110 327020 330116 327032
rect 330168 327020 330174 327072
rect 357618 326476 357624 326528
rect 357676 326516 357682 326528
rect 357894 326516 357900 326528
rect 357676 326488 357900 326516
rect 357676 326476 357682 326488
rect 357894 326476 357900 326488
rect 357952 326476 357958 326528
rect 358630 325728 358636 325780
rect 358688 325768 358694 325780
rect 358722 325768 358728 325780
rect 358688 325740 358728 325768
rect 358688 325728 358694 325740
rect 358722 325728 358728 325740
rect 358780 325728 358786 325780
rect 262674 325660 262680 325712
rect 262732 325700 262738 325712
rect 262858 325700 262864 325712
rect 262732 325672 262864 325700
rect 262732 325660 262738 325672
rect 262858 325660 262864 325672
rect 262916 325660 262922 325712
rect 265250 325660 265256 325712
rect 265308 325700 265314 325712
rect 265308 325672 265353 325700
rect 265308 325660 265314 325672
rect 463694 325660 463700 325712
rect 463752 325700 463758 325712
rect 463878 325700 463884 325712
rect 463752 325672 463884 325700
rect 463752 325660 463758 325672
rect 463878 325660 463884 325672
rect 463936 325660 463942 325712
rect 358538 325592 358544 325644
rect 358596 325632 358602 325644
rect 358630 325632 358636 325644
rect 358596 325604 358636 325632
rect 358596 325592 358602 325604
rect 358630 325592 358636 325604
rect 358688 325592 358694 325644
rect 3326 324232 3332 324284
rect 3384 324272 3390 324284
rect 14458 324272 14464 324284
rect 3384 324244 14464 324272
rect 3384 324232 3390 324244
rect 14458 324232 14464 324244
rect 14516 324232 14522 324284
rect 470042 322872 470048 322924
rect 470100 322912 470106 322924
rect 579982 322912 579988 322924
rect 470100 322884 579988 322912
rect 470100 322872 470106 322884
rect 579982 322872 579988 322884
rect 580040 322872 580046 322924
rect 236454 321688 236460 321700
rect 236415 321660 236460 321688
rect 236454 321648 236460 321660
rect 236512 321648 236518 321700
rect 244458 321620 244464 321632
rect 244384 321592 244464 321620
rect 244384 321564 244412 321592
rect 244458 321580 244464 321592
rect 244516 321580 244522 321632
rect 310790 321580 310796 321632
rect 310848 321580 310854 321632
rect 337378 321620 337384 321632
rect 337339 321592 337384 321620
rect 337378 321580 337384 321592
rect 337436 321580 337442 321632
rect 375834 321580 375840 321632
rect 375892 321580 375898 321632
rect 377122 321580 377128 321632
rect 377180 321580 377186 321632
rect 244366 321512 244372 321564
rect 244424 321512 244430 321564
rect 273530 321552 273536 321564
rect 273491 321524 273536 321552
rect 273530 321512 273536 321524
rect 273588 321512 273594 321564
rect 310808 321484 310836 321580
rect 310882 321484 310888 321496
rect 310808 321456 310888 321484
rect 310882 321444 310888 321456
rect 310940 321444 310946 321496
rect 375852 321416 375880 321580
rect 375926 321416 375932 321428
rect 375852 321388 375932 321416
rect 375926 321376 375932 321388
rect 375984 321376 375990 321428
rect 377140 321416 377168 321580
rect 377214 321416 377220 321428
rect 377140 321388 377220 321416
rect 377214 321376 377220 321388
rect 377272 321376 377278 321428
rect 359182 318900 359188 318912
rect 359108 318872 359188 318900
rect 359108 318844 359136 318872
rect 359182 318860 359188 318872
rect 359240 318860 359246 318912
rect 362310 318900 362316 318912
rect 362236 318872 362316 318900
rect 362236 318844 362264 318872
rect 362310 318860 362316 318872
rect 362368 318860 362374 318912
rect 236454 318832 236460 318844
rect 236415 318804 236460 318832
rect 236454 318792 236460 318804
rect 236512 318792 236518 318844
rect 259825 318835 259883 318841
rect 259825 318801 259837 318835
rect 259871 318832 259883 318835
rect 259914 318832 259920 318844
rect 259871 318804 259920 318832
rect 259871 318801 259883 318804
rect 259825 318795 259883 318801
rect 259914 318792 259920 318804
rect 259972 318792 259978 318844
rect 299842 318792 299848 318844
rect 299900 318832 299906 318844
rect 300210 318832 300216 318844
rect 299900 318804 300216 318832
rect 299900 318792 299906 318804
rect 300210 318792 300216 318804
rect 300268 318792 300274 318844
rect 302602 318832 302608 318844
rect 302563 318804 302608 318832
rect 302602 318792 302608 318804
rect 302660 318792 302666 318844
rect 330113 318835 330171 318841
rect 330113 318801 330125 318835
rect 330159 318832 330171 318835
rect 330202 318832 330208 318844
rect 330159 318804 330208 318832
rect 330159 318801 330171 318804
rect 330113 318795 330171 318801
rect 330202 318792 330208 318804
rect 330260 318792 330266 318844
rect 337378 318832 337384 318844
rect 337339 318804 337384 318832
rect 337378 318792 337384 318804
rect 337436 318792 337442 318844
rect 339770 318832 339776 318844
rect 339731 318804 339776 318832
rect 339770 318792 339776 318804
rect 339828 318792 339834 318844
rect 341337 318835 341395 318841
rect 341337 318801 341349 318835
rect 341383 318832 341395 318835
rect 341426 318832 341432 318844
rect 341383 318804 341432 318832
rect 341383 318801 341395 318804
rect 341337 318795 341395 318801
rect 341426 318792 341432 318804
rect 341484 318792 341490 318844
rect 359090 318792 359096 318844
rect 359148 318792 359154 318844
rect 362218 318792 362224 318844
rect 362276 318792 362282 318844
rect 389453 318835 389511 318841
rect 389453 318801 389465 318835
rect 389499 318832 389511 318835
rect 389542 318832 389548 318844
rect 389499 318804 389548 318832
rect 389499 318801 389511 318804
rect 389453 318795 389511 318801
rect 389542 318792 389548 318804
rect 389600 318792 389606 318844
rect 424594 318792 424600 318844
rect 424652 318832 424658 318844
rect 424686 318832 424692 318844
rect 424652 318804 424692 318832
rect 424652 318792 424658 318804
rect 424686 318792 424692 318804
rect 424744 318792 424750 318844
rect 470594 318832 470600 318844
rect 470555 318804 470600 318832
rect 470594 318792 470600 318804
rect 470652 318792 470658 318844
rect 372706 318764 372712 318776
rect 372667 318736 372712 318764
rect 372706 318724 372712 318736
rect 372764 318724 372770 318776
rect 288805 318631 288863 318637
rect 288805 318597 288817 318631
rect 288851 318628 288863 318631
rect 288986 318628 288992 318640
rect 288851 318600 288992 318628
rect 288851 318597 288863 318600
rect 288805 318591 288863 318597
rect 288986 318588 288992 318600
rect 289044 318588 289050 318640
rect 285950 317540 285956 317552
rect 285911 317512 285956 317540
rect 285950 317500 285956 317512
rect 286008 317500 286014 317552
rect 306742 317472 306748 317484
rect 306703 317444 306748 317472
rect 306742 317432 306748 317444
rect 306800 317432 306806 317484
rect 236270 317364 236276 317416
rect 236328 317404 236334 317416
rect 236454 317404 236460 317416
rect 236328 317376 236460 317404
rect 236328 317364 236334 317376
rect 236454 317364 236460 317376
rect 236512 317364 236518 317416
rect 250162 317404 250168 317416
rect 250123 317376 250168 317404
rect 250162 317364 250168 317376
rect 250220 317364 250226 317416
rect 251542 317404 251548 317416
rect 251503 317376 251548 317404
rect 251542 317364 251548 317376
rect 251600 317364 251606 317416
rect 266630 317364 266636 317416
rect 266688 317404 266694 317416
rect 266722 317404 266728 317416
rect 266688 317376 266728 317404
rect 266688 317364 266694 317376
rect 266722 317364 266728 317376
rect 266780 317364 266786 317416
rect 267734 317364 267740 317416
rect 267792 317404 267798 317416
rect 267826 317404 267832 317416
rect 267792 317376 267832 317404
rect 267792 317364 267798 317376
rect 267826 317364 267832 317376
rect 267884 317364 267890 317416
rect 273254 317364 273260 317416
rect 273312 317404 273318 317416
rect 273530 317404 273536 317416
rect 273312 317376 273536 317404
rect 273312 317364 273318 317376
rect 273530 317364 273536 317376
rect 273588 317364 273594 317416
rect 299753 317407 299811 317413
rect 299753 317373 299765 317407
rect 299799 317404 299811 317407
rect 299842 317404 299848 317416
rect 299799 317376 299848 317404
rect 299799 317373 299811 317376
rect 299753 317367 299811 317373
rect 299842 317364 299848 317376
rect 299900 317364 299906 317416
rect 325881 317407 325939 317413
rect 325881 317373 325893 317407
rect 325927 317404 325939 317407
rect 325970 317404 325976 317416
rect 325927 317376 325976 317404
rect 325927 317373 325939 317376
rect 325881 317367 325939 317373
rect 325970 317364 325976 317376
rect 326028 317364 326034 317416
rect 421190 317404 421196 317416
rect 421151 317376 421196 317404
rect 421190 317364 421196 317376
rect 421248 317364 421254 317416
rect 245838 316004 245844 316056
rect 245896 316044 245902 316056
rect 246114 316044 246120 316056
rect 245896 316016 246120 316044
rect 245896 316004 245902 316016
rect 246114 316004 246120 316016
rect 246172 316004 246178 316056
rect 265158 316004 265164 316056
rect 265216 316044 265222 316056
rect 265342 316044 265348 316056
rect 265216 316016 265348 316044
rect 265216 316004 265222 316016
rect 265342 316004 265348 316016
rect 265400 316004 265406 316056
rect 301130 316004 301136 316056
rect 301188 316044 301194 316056
rect 301314 316044 301320 316056
rect 301188 316016 301320 316044
rect 301188 316004 301194 316016
rect 301314 316004 301320 316016
rect 301372 316004 301378 316056
rect 306742 316044 306748 316056
rect 306703 316016 306748 316044
rect 306742 316004 306748 316016
rect 306800 316004 306806 316056
rect 357434 316004 357440 316056
rect 357492 316044 357498 316056
rect 357618 316044 357624 316056
rect 357492 316016 357624 316044
rect 357492 316004 357498 316016
rect 357618 316004 357624 316016
rect 357676 316004 357682 316056
rect 244366 315936 244372 315988
rect 244424 315936 244430 315988
rect 244384 315840 244412 315936
rect 244550 315840 244556 315852
rect 244384 315812 244556 315840
rect 244550 315800 244556 315812
rect 244608 315800 244614 315852
rect 290090 313256 290096 313268
rect 290051 313228 290096 313256
rect 290090 313216 290096 313228
rect 290148 313216 290154 313268
rect 302602 311964 302608 311976
rect 302528 311936 302608 311964
rect 239030 311856 239036 311908
rect 239088 311896 239094 311908
rect 239214 311896 239220 311908
rect 239088 311868 239220 311896
rect 239088 311856 239094 311868
rect 239214 311856 239220 311868
rect 239272 311856 239278 311908
rect 284573 311899 284631 311905
rect 284573 311865 284585 311899
rect 284619 311896 284631 311899
rect 284662 311896 284668 311908
rect 284619 311868 284668 311896
rect 284619 311865 284631 311868
rect 284573 311859 284631 311865
rect 284662 311856 284668 311868
rect 284720 311856 284726 311908
rect 285950 311896 285956 311908
rect 285911 311868 285956 311896
rect 285950 311856 285956 311868
rect 286008 311856 286014 311908
rect 302528 311840 302556 311936
rect 302602 311924 302608 311936
rect 302660 311924 302666 311976
rect 310882 311964 310888 311976
rect 310843 311936 310888 311964
rect 310882 311924 310888 311936
rect 310940 311924 310946 311976
rect 323302 311964 323308 311976
rect 323228 311936 323308 311964
rect 323228 311908 323256 311936
rect 323302 311924 323308 311936
rect 323360 311924 323366 311976
rect 323210 311856 323216 311908
rect 323268 311856 323274 311908
rect 337194 311856 337200 311908
rect 337252 311896 337258 311908
rect 337378 311896 337384 311908
rect 337252 311868 337384 311896
rect 337252 311856 337258 311868
rect 337378 311856 337384 311868
rect 337436 311856 337442 311908
rect 341242 311856 341248 311908
rect 341300 311896 341306 311908
rect 341426 311896 341432 311908
rect 341300 311868 341432 311896
rect 341300 311856 341306 311868
rect 341426 311856 341432 311868
rect 341484 311856 341490 311908
rect 360194 311856 360200 311908
rect 360252 311896 360258 311908
rect 360562 311896 360568 311908
rect 360252 311868 360568 311896
rect 360252 311856 360258 311868
rect 360562 311856 360568 311868
rect 360620 311856 360626 311908
rect 424134 311856 424140 311908
rect 424192 311896 424198 311908
rect 424594 311896 424600 311908
rect 424192 311868 424600 311896
rect 424192 311856 424198 311868
rect 424594 311856 424600 311868
rect 424652 311856 424658 311908
rect 302510 311788 302516 311840
rect 302568 311788 302574 311840
rect 339678 311788 339684 311840
rect 339736 311828 339742 311840
rect 339862 311828 339868 311840
rect 339736 311800 339868 311828
rect 339736 311788 339742 311800
rect 339862 311788 339868 311800
rect 339920 311788 339926 311840
rect 291470 309136 291476 309188
rect 291528 309176 291534 309188
rect 291562 309176 291568 309188
rect 291528 309148 291568 309176
rect 291528 309136 291534 309148
rect 291562 309136 291568 309148
rect 291620 309136 291626 309188
rect 372706 309176 372712 309188
rect 372667 309148 372712 309176
rect 372706 309136 372712 309148
rect 372764 309136 372770 309188
rect 389358 309136 389364 309188
rect 389416 309176 389422 309188
rect 389542 309176 389548 309188
rect 389416 309148 389548 309176
rect 389416 309136 389422 309148
rect 389542 309136 389548 309148
rect 389600 309136 389606 309188
rect 239122 309108 239128 309120
rect 239083 309080 239128 309108
rect 239122 309068 239128 309080
rect 239180 309068 239186 309120
rect 327166 309068 327172 309120
rect 327224 309108 327230 309120
rect 327258 309108 327264 309120
rect 327224 309080 327264 309108
rect 327224 309068 327230 309080
rect 327258 309068 327264 309080
rect 327316 309068 327322 309120
rect 339862 309108 339868 309120
rect 339823 309080 339868 309108
rect 339862 309068 339868 309080
rect 339920 309068 339926 309120
rect 341153 309111 341211 309117
rect 341153 309077 341165 309111
rect 341199 309108 341211 309111
rect 341242 309108 341248 309120
rect 341199 309080 341248 309108
rect 341199 309077 341211 309080
rect 341153 309071 341211 309077
rect 341242 309068 341248 309080
rect 341300 309068 341306 309120
rect 360194 309068 360200 309120
rect 360252 309108 360258 309120
rect 360286 309108 360292 309120
rect 360252 309080 360292 309108
rect 360252 309068 360258 309080
rect 360286 309068 360292 309080
rect 360344 309068 360350 309120
rect 367002 309108 367008 309120
rect 366963 309080 367008 309108
rect 367002 309068 367008 309080
rect 367060 309068 367066 309120
rect 470594 309108 470600 309120
rect 470555 309080 470600 309108
rect 470594 309068 470600 309080
rect 470652 309068 470658 309120
rect 389269 309043 389327 309049
rect 389269 309009 389281 309043
rect 389315 309040 389327 309043
rect 389358 309040 389364 309052
rect 389315 309012 389364 309040
rect 389315 309009 389327 309012
rect 389269 309003 389327 309009
rect 389358 309000 389364 309012
rect 389416 309000 389422 309052
rect 2774 308796 2780 308848
rect 2832 308836 2838 308848
rect 5350 308836 5356 308848
rect 2832 308808 5356 308836
rect 2832 308796 2838 308808
rect 5350 308796 5356 308808
rect 5408 308796 5414 308848
rect 288713 308431 288771 308437
rect 288713 308397 288725 308431
rect 288759 308428 288771 308431
rect 288986 308428 288992 308440
rect 288759 308400 288992 308428
rect 288759 308397 288771 308400
rect 288713 308391 288771 308397
rect 288986 308388 288992 308400
rect 289044 308388 289050 308440
rect 310698 307844 310704 307896
rect 310756 307884 310762 307896
rect 310885 307887 310943 307893
rect 310885 307884 310897 307887
rect 310756 307856 310897 307884
rect 310756 307844 310762 307856
rect 310885 307853 310897 307856
rect 310931 307853 310943 307887
rect 310885 307847 310943 307853
rect 250162 307816 250168 307828
rect 250123 307788 250168 307816
rect 250162 307776 250168 307788
rect 250220 307776 250226 307828
rect 251542 307816 251548 307828
rect 251503 307788 251548 307816
rect 251542 307776 251548 307788
rect 251600 307776 251606 307828
rect 259730 307776 259736 307828
rect 259788 307816 259794 307828
rect 259914 307816 259920 307828
rect 259788 307788 259920 307816
rect 259788 307776 259794 307788
rect 259914 307776 259920 307788
rect 259972 307776 259978 307828
rect 301130 307776 301136 307828
rect 301188 307776 301194 307828
rect 306742 307776 306748 307828
rect 306800 307776 306806 307828
rect 325878 307816 325884 307828
rect 325839 307788 325884 307816
rect 325878 307776 325884 307788
rect 325936 307776 325942 307828
rect 421190 307816 421196 307828
rect 421151 307788 421196 307816
rect 421190 307776 421196 307788
rect 421248 307776 421254 307828
rect 232314 307748 232320 307760
rect 232275 307720 232320 307748
rect 232314 307708 232320 307720
rect 232372 307708 232378 307760
rect 301148 307680 301176 307776
rect 301222 307680 301228 307692
rect 301148 307652 301228 307680
rect 301222 307640 301228 307652
rect 301280 307640 301286 307692
rect 306760 307680 306788 307776
rect 310698 307748 310704 307760
rect 310659 307720 310704 307748
rect 310698 307708 310704 307720
rect 310756 307708 310762 307760
rect 337013 307751 337071 307757
rect 337013 307717 337025 307751
rect 337059 307748 337071 307751
rect 337194 307748 337200 307760
rect 337059 307720 337200 307748
rect 337059 307717 337071 307720
rect 337013 307711 337071 307717
rect 337194 307708 337200 307720
rect 337252 307708 337258 307760
rect 306926 307680 306932 307692
rect 306760 307652 306932 307680
rect 306926 307640 306932 307652
rect 306984 307640 306990 307692
rect 285766 306416 285772 306468
rect 285824 306456 285830 306468
rect 285953 306459 286011 306465
rect 285953 306456 285965 306459
rect 285824 306428 285965 306456
rect 285824 306416 285830 306428
rect 285953 306425 285965 306428
rect 285999 306425 286011 306459
rect 285953 306419 286011 306425
rect 267826 306348 267832 306400
rect 267884 306388 267890 306400
rect 268010 306388 268016 306400
rect 267884 306360 268016 306388
rect 267884 306348 267890 306360
rect 268010 306348 268016 306360
rect 268068 306348 268074 306400
rect 273070 306348 273076 306400
rect 273128 306388 273134 306400
rect 273254 306388 273260 306400
rect 273128 306360 273260 306388
rect 273128 306348 273134 306360
rect 273254 306348 273260 306360
rect 273312 306348 273318 306400
rect 284570 306388 284576 306400
rect 284531 306360 284576 306388
rect 284570 306348 284576 306360
rect 284628 306348 284634 306400
rect 317506 306348 317512 306400
rect 317564 306388 317570 306400
rect 317690 306388 317696 306400
rect 317564 306360 317696 306388
rect 317564 306348 317570 306360
rect 317690 306348 317696 306360
rect 317748 306348 317754 306400
rect 330202 306348 330208 306400
rect 330260 306388 330266 306400
rect 330386 306388 330392 306400
rect 330260 306360 330392 306388
rect 330260 306348 330266 306360
rect 330386 306348 330392 306360
rect 330444 306348 330450 306400
rect 358538 306348 358544 306400
rect 358596 306388 358602 306400
rect 358722 306388 358728 306400
rect 358596 306360 358728 306388
rect 358596 306348 358602 306360
rect 358722 306348 358728 306360
rect 358780 306348 358786 306400
rect 463694 306348 463700 306400
rect 463752 306388 463758 306400
rect 463878 306388 463884 306400
rect 463752 306360 463884 306388
rect 463752 306348 463758 306360
rect 463878 306348 463884 306360
rect 463936 306348 463942 306400
rect 290093 306323 290151 306329
rect 290093 306289 290105 306323
rect 290139 306320 290151 306323
rect 290182 306320 290188 306332
rect 290139 306292 290188 306320
rect 290139 306289 290151 306292
rect 290093 306283 290151 306289
rect 290182 306280 290188 306292
rect 290240 306280 290246 306332
rect 294322 304920 294328 304972
rect 294380 304920 294386 304972
rect 294230 304852 294236 304904
rect 294288 304892 294294 304904
rect 294340 304892 294368 304920
rect 294288 304864 294368 304892
rect 294288 304852 294294 304864
rect 245930 302444 245936 302456
rect 245891 302416 245936 302444
rect 245930 302404 245936 302416
rect 245988 302404 245994 302456
rect 270678 302268 270684 302320
rect 270736 302268 270742 302320
rect 272150 302268 272156 302320
rect 272208 302268 272214 302320
rect 330202 302308 330208 302320
rect 330128 302280 330208 302308
rect 270696 302104 270724 302268
rect 270770 302104 270776 302116
rect 270696 302076 270776 302104
rect 270770 302064 270776 302076
rect 270828 302064 270834 302116
rect 272168 302104 272196 302268
rect 330128 302184 330156 302280
rect 330202 302268 330208 302280
rect 330260 302268 330266 302320
rect 424134 302200 424140 302252
rect 424192 302240 424198 302252
rect 424502 302240 424508 302252
rect 424192 302212 424508 302240
rect 424192 302200 424198 302212
rect 424502 302200 424508 302212
rect 424560 302200 424566 302252
rect 330110 302132 330116 302184
rect 330168 302132 330174 302184
rect 272242 302104 272248 302116
rect 272168 302076 272248 302104
rect 272242 302064 272248 302076
rect 272300 302064 272306 302116
rect 339862 299928 339868 299940
rect 339823 299900 339868 299928
rect 339862 299888 339868 299900
rect 339920 299888 339926 299940
rect 239125 299523 239183 299529
rect 239125 299489 239137 299523
rect 239171 299520 239183 299523
rect 239214 299520 239220 299532
rect 239171 299492 239220 299520
rect 239171 299489 239183 299492
rect 239125 299483 239183 299489
rect 239214 299480 239220 299492
rect 239272 299480 239278 299532
rect 299753 299523 299811 299529
rect 299753 299489 299765 299523
rect 299799 299520 299811 299523
rect 299842 299520 299848 299532
rect 299799 299492 299848 299520
rect 299799 299489 299811 299492
rect 299753 299483 299811 299489
rect 299842 299480 299848 299492
rect 299900 299480 299906 299532
rect 302510 299480 302516 299532
rect 302568 299520 302574 299532
rect 302602 299520 302608 299532
rect 302568 299492 302608 299520
rect 302568 299480 302574 299492
rect 302602 299480 302608 299492
rect 302660 299480 302666 299532
rect 306834 299520 306840 299532
rect 306795 299492 306840 299520
rect 306834 299480 306840 299492
rect 306892 299480 306898 299532
rect 341150 299520 341156 299532
rect 341111 299492 341156 299520
rect 341150 299480 341156 299492
rect 341208 299480 341214 299532
rect 367002 299520 367008 299532
rect 366963 299492 367008 299520
rect 367002 299480 367008 299492
rect 367060 299480 367066 299532
rect 389266 299520 389272 299532
rect 389227 299492 389272 299520
rect 389266 299480 389272 299492
rect 389324 299480 389330 299532
rect 470594 299520 470600 299532
rect 470555 299492 470600 299520
rect 470594 299480 470600 299492
rect 470652 299480 470658 299532
rect 323302 299452 323308 299464
rect 323263 299424 323308 299452
rect 323302 299412 323308 299424
rect 323360 299412 323366 299464
rect 324682 299452 324688 299464
rect 324643 299424 324688 299452
rect 324682 299412 324688 299424
rect 324740 299412 324746 299464
rect 325878 299412 325884 299464
rect 325936 299412 325942 299464
rect 372706 299452 372712 299464
rect 372667 299424 372712 299452
rect 372706 299412 372712 299424
rect 372764 299412 372770 299464
rect 469950 299412 469956 299464
rect 470008 299452 470014 299464
rect 579798 299452 579804 299464
rect 470008 299424 579804 299452
rect 470008 299412 470014 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 325896 299384 325924 299412
rect 325970 299384 325976 299396
rect 325896 299356 325976 299384
rect 325970 299344 325976 299356
rect 326028 299344 326034 299396
rect 295610 298228 295616 298240
rect 295536 298200 295616 298228
rect 232314 298160 232320 298172
rect 232275 298132 232320 298160
rect 232314 298120 232320 298132
rect 232372 298120 232378 298172
rect 262490 298120 262496 298172
rect 262548 298160 262554 298172
rect 262674 298160 262680 298172
rect 262548 298132 262680 298160
rect 262548 298120 262554 298132
rect 262674 298120 262680 298132
rect 262732 298120 262738 298172
rect 236270 298092 236276 298104
rect 236231 298064 236276 298092
rect 236270 298052 236276 298064
rect 236328 298052 236334 298104
rect 250162 298092 250168 298104
rect 250123 298064 250168 298092
rect 250162 298052 250168 298064
rect 250220 298052 250226 298104
rect 251361 298095 251419 298101
rect 251361 298061 251373 298095
rect 251407 298092 251419 298095
rect 251542 298092 251548 298104
rect 251407 298064 251548 298092
rect 251407 298061 251419 298064
rect 251361 298055 251419 298061
rect 251542 298052 251548 298064
rect 251600 298052 251606 298104
rect 295536 298036 295564 298200
rect 295610 298188 295616 298200
rect 295668 298188 295674 298240
rect 337010 298228 337016 298240
rect 336971 298200 337016 298228
rect 337010 298188 337016 298200
rect 337068 298188 337074 298240
rect 358722 298228 358728 298240
rect 358648 298200 358728 298228
rect 358648 298172 358676 298200
rect 358722 298188 358728 298200
rect 358780 298188 358786 298240
rect 310701 298163 310759 298169
rect 310701 298129 310713 298163
rect 310747 298160 310759 298163
rect 310882 298160 310888 298172
rect 310747 298132 310888 298160
rect 310747 298129 310759 298132
rect 310701 298123 310759 298129
rect 310882 298120 310888 298132
rect 310940 298120 310946 298172
rect 358630 298120 358636 298172
rect 358688 298120 358694 298172
rect 325970 298092 325976 298104
rect 325931 298064 325976 298092
rect 325970 298052 325976 298064
rect 326028 298052 326034 298104
rect 327169 298095 327227 298101
rect 327169 298061 327181 298095
rect 327215 298092 327227 298095
rect 327258 298092 327264 298104
rect 327215 298064 327264 298092
rect 327215 298061 327227 298064
rect 327169 298055 327227 298061
rect 327258 298052 327264 298064
rect 327316 298052 327322 298104
rect 337010 298052 337016 298104
rect 337068 298092 337074 298104
rect 337197 298095 337255 298101
rect 337197 298092 337209 298095
rect 337068 298064 337209 298092
rect 337068 298052 337074 298064
rect 337197 298061 337209 298064
rect 337243 298061 337255 298095
rect 337197 298055 337255 298061
rect 359090 298052 359096 298104
rect 359148 298092 359154 298104
rect 359182 298092 359188 298104
rect 359148 298064 359188 298092
rect 359148 298052 359154 298064
rect 359182 298052 359188 298064
rect 359240 298052 359246 298104
rect 421190 298092 421196 298104
rect 421151 298064 421196 298092
rect 421190 298052 421196 298064
rect 421248 298052 421254 298104
rect 232225 298027 232283 298033
rect 232225 297993 232237 298027
rect 232271 298024 232283 298027
rect 232314 298024 232320 298036
rect 232271 297996 232320 298024
rect 232271 297993 232283 297996
rect 232225 297987 232283 297993
rect 232314 297984 232320 297996
rect 232372 297984 232378 298036
rect 245933 298027 245991 298033
rect 245933 297993 245945 298027
rect 245979 298024 245991 298027
rect 246022 298024 246028 298036
rect 245979 297996 246028 298024
rect 245979 297993 245991 297996
rect 245933 297987 245991 297993
rect 246022 297984 246028 297996
rect 246080 297984 246086 298036
rect 295518 297984 295524 298036
rect 295576 297984 295582 298036
rect 273254 296692 273260 296744
rect 273312 296732 273318 296744
rect 273530 296732 273536 296744
rect 273312 296704 273536 296732
rect 273312 296692 273318 296704
rect 273530 296692 273536 296704
rect 273588 296692 273594 296744
rect 285766 296692 285772 296744
rect 285824 296732 285830 296744
rect 286042 296732 286048 296744
rect 285824 296704 286048 296732
rect 285824 296692 285830 296704
rect 286042 296692 286048 296704
rect 286100 296692 286106 296744
rect 296806 296692 296812 296744
rect 296864 296732 296870 296744
rect 296898 296732 296904 296744
rect 296864 296704 296904 296732
rect 296864 296692 296870 296704
rect 296898 296692 296904 296704
rect 296956 296692 296962 296744
rect 301038 296692 301044 296744
rect 301096 296732 301102 296744
rect 301406 296732 301412 296744
rect 301096 296704 301412 296732
rect 301096 296692 301102 296704
rect 301406 296692 301412 296704
rect 301464 296692 301470 296744
rect 306834 296732 306840 296744
rect 306795 296704 306840 296732
rect 306834 296692 306840 296704
rect 306892 296692 306898 296744
rect 362218 296692 362224 296744
rect 362276 296732 362282 296744
rect 362402 296732 362408 296744
rect 362276 296704 362408 296732
rect 362276 296692 362282 296704
rect 362402 296692 362408 296704
rect 362460 296692 362466 296744
rect 273622 296664 273628 296676
rect 273583 296636 273628 296664
rect 273622 296624 273628 296636
rect 273680 296624 273686 296676
rect 299842 296624 299848 296676
rect 299900 296664 299906 296676
rect 299934 296664 299940 296676
rect 299900 296636 299940 296664
rect 299900 296624 299906 296636
rect 299934 296624 299940 296636
rect 299992 296624 299998 296676
rect 302602 296624 302608 296676
rect 302660 296664 302666 296676
rect 302694 296664 302700 296676
rect 302660 296636 302700 296664
rect 302660 296624 302666 296636
rect 302694 296624 302700 296636
rect 302752 296624 302758 296676
rect 310882 293060 310888 293072
rect 310843 293032 310888 293060
rect 310882 293020 310888 293032
rect 310940 293020 310946 293072
rect 306834 292652 306840 292664
rect 306760 292624 306840 292652
rect 239030 292544 239036 292596
rect 239088 292584 239094 292596
rect 239214 292584 239220 292596
rect 239088 292556 239220 292584
rect 239088 292544 239094 292556
rect 239214 292544 239220 292556
rect 239272 292544 239278 292596
rect 306760 292528 306788 292624
rect 306834 292612 306840 292624
rect 306892 292612 306898 292664
rect 306742 292476 306748 292528
rect 306800 292476 306806 292528
rect 337194 292448 337200 292460
rect 337155 292420 337200 292448
rect 337194 292408 337200 292420
rect 337252 292408 337258 292460
rect 285766 291864 285772 291916
rect 285824 291904 285830 291916
rect 286042 291904 286048 291916
rect 285824 291876 286048 291904
rect 285824 291864 285830 291876
rect 286042 291864 286048 291876
rect 286100 291864 286106 291916
rect 288710 290000 288716 290012
rect 288671 289972 288716 290000
rect 288710 289960 288716 289972
rect 288768 289960 288774 290012
rect 262490 289824 262496 289876
rect 262548 289864 262554 289876
rect 262674 289864 262680 289876
rect 262548 289836 262680 289864
rect 262548 289824 262554 289836
rect 262674 289824 262680 289836
rect 262732 289824 262738 289876
rect 267826 289824 267832 289876
rect 267884 289864 267890 289876
rect 267918 289864 267924 289876
rect 267884 289836 267924 289864
rect 267884 289824 267890 289836
rect 267918 289824 267924 289836
rect 267976 289824 267982 289876
rect 324682 289864 324688 289876
rect 324643 289836 324688 289864
rect 324682 289824 324688 289836
rect 324740 289824 324746 289876
rect 372706 289864 372712 289876
rect 372667 289836 372712 289864
rect 372706 289824 372712 289836
rect 372764 289824 372770 289876
rect 375834 289824 375840 289876
rect 375892 289864 375898 289876
rect 375926 289864 375932 289876
rect 375892 289836 375932 289864
rect 375892 289824 375898 289836
rect 375926 289824 375932 289836
rect 375984 289824 375990 289876
rect 377122 289824 377128 289876
rect 377180 289864 377186 289876
rect 377214 289864 377220 289876
rect 377180 289836 377220 289864
rect 377180 289824 377186 289836
rect 377214 289824 377220 289836
rect 377272 289824 377278 289876
rect 250162 289796 250168 289808
rect 250123 289768 250168 289796
rect 250162 289756 250168 289768
rect 250220 289756 250226 289808
rect 270678 289756 270684 289808
rect 270736 289796 270742 289808
rect 270770 289796 270776 289808
rect 270736 289768 270776 289796
rect 270736 289756 270742 289768
rect 270770 289756 270776 289768
rect 270828 289756 270834 289808
rect 272153 289799 272211 289805
rect 272153 289765 272165 289799
rect 272199 289796 272211 289799
rect 272242 289796 272248 289808
rect 272199 289768 272248 289796
rect 272199 289765 272211 289768
rect 272153 289759 272211 289765
rect 272242 289756 272248 289768
rect 272300 289756 272306 289808
rect 284570 289756 284576 289808
rect 284628 289756 284634 289808
rect 288710 289756 288716 289808
rect 288768 289796 288774 289808
rect 288802 289796 288808 289808
rect 288768 289768 288808 289796
rect 288768 289756 288774 289768
rect 288802 289756 288808 289768
rect 288860 289756 288866 289808
rect 341153 289799 341211 289805
rect 341153 289765 341165 289799
rect 341199 289796 341211 289799
rect 341242 289796 341248 289808
rect 341199 289768 341248 289796
rect 341199 289765 341211 289768
rect 341153 289759 341211 289765
rect 341242 289756 341248 289768
rect 341300 289756 341306 289808
rect 367002 289796 367008 289808
rect 366963 289768 367008 289796
rect 367002 289756 367008 289768
rect 367060 289756 367066 289808
rect 389361 289799 389419 289805
rect 389361 289765 389373 289799
rect 389407 289796 389419 289799
rect 389450 289796 389456 289808
rect 389407 289768 389456 289796
rect 389407 289765 389419 289768
rect 389361 289759 389419 289765
rect 389450 289756 389456 289768
rect 389508 289756 389514 289808
rect 470594 289796 470600 289808
rect 470555 289768 470600 289796
rect 470594 289756 470600 289768
rect 470652 289756 470658 289808
rect 284588 289728 284616 289756
rect 284754 289728 284760 289740
rect 284588 289700 284760 289728
rect 284754 289688 284760 289700
rect 284812 289688 284818 289740
rect 232222 288436 232228 288448
rect 232183 288408 232228 288436
rect 232222 288396 232228 288408
rect 232280 288396 232286 288448
rect 236270 288436 236276 288448
rect 236231 288408 236276 288436
rect 236270 288396 236276 288408
rect 236328 288396 236334 288448
rect 251358 288436 251364 288448
rect 251319 288408 251364 288436
rect 251358 288396 251364 288408
rect 251416 288396 251422 288448
rect 323305 288439 323363 288445
rect 323305 288405 323317 288439
rect 323351 288436 323363 288439
rect 323486 288436 323492 288448
rect 323351 288408 323492 288436
rect 323351 288405 323363 288408
rect 323305 288399 323363 288405
rect 323486 288396 323492 288408
rect 323544 288396 323550 288448
rect 325970 288436 325976 288448
rect 325931 288408 325976 288436
rect 325970 288396 325976 288408
rect 326028 288396 326034 288448
rect 327166 288436 327172 288448
rect 327127 288408 327172 288436
rect 327166 288396 327172 288408
rect 327224 288396 327230 288448
rect 330294 288436 330300 288448
rect 330255 288408 330300 288436
rect 330294 288396 330300 288408
rect 330352 288396 330358 288448
rect 357434 288396 357440 288448
rect 357492 288436 357498 288448
rect 357618 288436 357624 288448
rect 357492 288408 357624 288436
rect 357492 288396 357498 288408
rect 357618 288396 357624 288408
rect 357676 288396 357682 288448
rect 358630 288396 358636 288448
rect 358688 288436 358694 288448
rect 358722 288436 358728 288448
rect 358688 288408 358728 288436
rect 358688 288396 358694 288408
rect 358722 288396 358728 288408
rect 358780 288396 358786 288448
rect 421190 288436 421196 288448
rect 421151 288408 421196 288436
rect 421190 288396 421196 288408
rect 421248 288396 421254 288448
rect 273622 287076 273628 287088
rect 273583 287048 273628 287076
rect 273622 287036 273628 287048
rect 273680 287036 273686 287088
rect 330294 287076 330300 287088
rect 330255 287048 330300 287076
rect 330294 287036 330300 287048
rect 330352 287036 330358 287088
rect 463694 287036 463700 287088
rect 463752 287076 463758 287088
rect 463878 287076 463884 287088
rect 463752 287048 463884 287076
rect 463752 287036 463758 287048
rect 463878 287036 463884 287048
rect 463936 287036 463942 287088
rect 259546 285608 259552 285660
rect 259604 285648 259610 285660
rect 259914 285648 259920 285660
rect 259604 285620 259920 285648
rect 259604 285608 259610 285620
rect 259914 285608 259920 285620
rect 259972 285608 259978 285660
rect 272153 283611 272211 283617
rect 272153 283577 272165 283611
rect 272199 283608 272211 283611
rect 272334 283608 272340 283620
rect 272199 283580 272340 283608
rect 272199 283577 272211 283580
rect 272153 283571 272211 283577
rect 272334 283568 272340 283580
rect 272392 283568 272398 283620
rect 236270 282888 236276 282940
rect 236328 282888 236334 282940
rect 239122 282888 239128 282940
rect 239180 282888 239186 282940
rect 337102 282928 337108 282940
rect 337063 282900 337108 282928
rect 337102 282888 337108 282900
rect 337160 282888 337166 282940
rect 339678 282888 339684 282940
rect 339736 282928 339742 282940
rect 339862 282928 339868 282940
rect 339736 282900 339868 282928
rect 339736 282888 339742 282900
rect 339862 282888 339868 282900
rect 339920 282888 339926 282940
rect 424502 282888 424508 282940
rect 424560 282928 424566 282940
rect 424686 282928 424692 282940
rect 424560 282900 424692 282928
rect 424560 282888 424566 282900
rect 424686 282888 424692 282900
rect 424744 282888 424750 282940
rect 236288 282792 236316 282888
rect 236454 282792 236460 282804
rect 236288 282764 236460 282792
rect 236454 282752 236460 282764
rect 236512 282752 236518 282804
rect 239140 282792 239168 282888
rect 239214 282792 239220 282804
rect 239140 282764 239220 282792
rect 239214 282752 239220 282764
rect 239272 282752 239278 282804
rect 310882 282792 310888 282804
rect 310843 282764 310888 282792
rect 310882 282752 310888 282764
rect 310940 282752 310946 282804
rect 232222 280168 232228 280220
rect 232280 280208 232286 280220
rect 232314 280208 232320 280220
rect 232280 280180 232320 280208
rect 232280 280168 232286 280180
rect 232314 280168 232320 280180
rect 232372 280168 232378 280220
rect 341150 280208 341156 280220
rect 341111 280180 341156 280208
rect 341150 280168 341156 280180
rect 341208 280168 341214 280220
rect 367002 280208 367008 280220
rect 366963 280180 367008 280208
rect 367002 280168 367008 280180
rect 367060 280168 367066 280220
rect 389358 280208 389364 280220
rect 389319 280180 389364 280208
rect 389358 280168 389364 280180
rect 389416 280168 389422 280220
rect 470594 280208 470600 280220
rect 470555 280180 470600 280208
rect 470594 280168 470600 280180
rect 470652 280168 470658 280220
rect 250070 280100 250076 280152
rect 250128 280140 250134 280152
rect 250162 280140 250168 280152
rect 250128 280112 250168 280140
rect 250128 280100 250134 280112
rect 250162 280100 250168 280112
rect 250220 280100 250226 280152
rect 270678 280140 270684 280152
rect 270639 280112 270684 280140
rect 270678 280100 270684 280112
rect 270736 280100 270742 280152
rect 273530 280140 273536 280152
rect 273491 280112 273536 280140
rect 273530 280100 273536 280112
rect 273588 280100 273594 280152
rect 284570 280100 284576 280152
rect 284628 280140 284634 280152
rect 284754 280140 284760 280152
rect 284628 280112 284760 280140
rect 284628 280100 284634 280112
rect 284754 280100 284760 280112
rect 284812 280100 284818 280152
rect 288802 280100 288808 280152
rect 288860 280140 288866 280152
rect 288894 280140 288900 280152
rect 288860 280112 288900 280140
rect 288860 280100 288866 280112
rect 288894 280100 288900 280112
rect 288952 280100 288958 280152
rect 323302 280100 323308 280152
rect 323360 280140 323366 280152
rect 323394 280140 323400 280152
rect 323360 280112 323400 280140
rect 323360 280100 323366 280112
rect 323394 280100 323400 280112
rect 323452 280100 323458 280152
rect 372706 280140 372712 280152
rect 372667 280112 372712 280140
rect 372706 280100 372712 280112
rect 372764 280100 372770 280152
rect 375834 280140 375840 280152
rect 375795 280112 375840 280140
rect 375834 280100 375840 280112
rect 375892 280100 375898 280152
rect 377122 280140 377128 280152
rect 377083 280112 377128 280140
rect 377122 280100 377128 280112
rect 377180 280100 377186 280152
rect 424594 280140 424600 280152
rect 424555 280112 424600 280140
rect 424594 280100 424600 280112
rect 424652 280100 424658 280152
rect 265158 278740 265164 278792
rect 265216 278780 265222 278792
rect 265250 278780 265256 278792
rect 265216 278752 265256 278780
rect 265216 278740 265222 278752
rect 265250 278740 265256 278752
rect 265308 278740 265314 278792
rect 267734 278740 267740 278792
rect 267792 278780 267798 278792
rect 267826 278780 267832 278792
rect 267792 278752 267832 278780
rect 267792 278740 267798 278752
rect 267826 278740 267832 278752
rect 267884 278740 267890 278792
rect 285766 278740 285772 278792
rect 285824 278780 285830 278792
rect 286042 278780 286048 278792
rect 285824 278752 286048 278780
rect 285824 278740 285830 278752
rect 286042 278740 286048 278752
rect 286100 278740 286106 278792
rect 295242 278740 295248 278792
rect 295300 278780 295306 278792
rect 295518 278780 295524 278792
rect 295300 278752 295524 278780
rect 295300 278740 295306 278752
rect 295518 278740 295524 278752
rect 295576 278740 295582 278792
rect 301038 278740 301044 278792
rect 301096 278780 301102 278792
rect 301222 278780 301228 278792
rect 301096 278752 301228 278780
rect 301096 278740 301102 278752
rect 301222 278740 301228 278752
rect 301280 278740 301286 278792
rect 327350 278740 327356 278792
rect 327408 278780 327414 278792
rect 327534 278780 327540 278792
rect 327408 278752 327540 278780
rect 327408 278740 327414 278752
rect 327534 278740 327540 278752
rect 327592 278740 327598 278792
rect 337102 278780 337108 278792
rect 337063 278752 337108 278780
rect 337102 278740 337108 278752
rect 337160 278740 337166 278792
rect 310882 278712 310888 278724
rect 310843 278684 310888 278712
rect 310882 278672 310888 278684
rect 310940 278672 310946 278724
rect 324498 278712 324504 278724
rect 324459 278684 324504 278712
rect 324498 278672 324504 278684
rect 324556 278672 324562 278724
rect 295518 277856 295524 277908
rect 295576 277896 295582 277908
rect 295794 277896 295800 277908
rect 295576 277868 295800 277896
rect 295576 277856 295582 277868
rect 295794 277856 295800 277868
rect 295852 277856 295858 277908
rect 307018 277488 307024 277500
rect 306852 277460 307024 277488
rect 306852 277432 306880 277460
rect 307018 277448 307024 277460
rect 307076 277448 307082 277500
rect 289998 277380 290004 277432
rect 290056 277420 290062 277432
rect 290090 277420 290096 277432
rect 290056 277392 290096 277420
rect 290056 277380 290062 277392
rect 290090 277380 290096 277392
rect 290148 277380 290154 277432
rect 296806 277380 296812 277432
rect 296864 277420 296870 277432
rect 297082 277420 297088 277432
rect 296864 277392 297088 277420
rect 296864 277380 296870 277392
rect 297082 277380 297088 277392
rect 297140 277380 297146 277432
rect 306834 277380 306840 277432
rect 306892 277380 306898 277432
rect 330110 277380 330116 277432
rect 330168 277420 330174 277432
rect 330294 277420 330300 277432
rect 330168 277392 330300 277420
rect 330168 277380 330174 277392
rect 330294 277380 330300 277392
rect 330352 277380 330358 277432
rect 357710 277380 357716 277432
rect 357768 277420 357774 277432
rect 357802 277420 357808 277432
rect 357768 277392 357808 277420
rect 357768 277380 357774 277392
rect 357802 277380 357808 277392
rect 357860 277380 357866 277432
rect 362218 277352 362224 277364
rect 362179 277324 362224 277352
rect 362218 277312 362224 277324
rect 362276 277312 362282 277364
rect 330110 277284 330116 277296
rect 330071 277256 330116 277284
rect 330110 277244 330116 277256
rect 330168 277244 330174 277296
rect 270678 275312 270684 275324
rect 270639 275284 270684 275312
rect 270678 275272 270684 275284
rect 270736 275272 270742 275324
rect 236270 273232 236276 273284
rect 236328 273272 236334 273284
rect 236454 273272 236460 273284
rect 236328 273244 236460 273272
rect 236328 273232 236334 273244
rect 236454 273232 236460 273244
rect 236512 273232 236518 273284
rect 239030 273232 239036 273284
rect 239088 273272 239094 273284
rect 239214 273272 239220 273284
rect 239088 273244 239220 273272
rect 239088 273232 239094 273244
rect 239214 273232 239220 273244
rect 239272 273232 239278 273284
rect 301038 273232 301044 273284
rect 301096 273232 301102 273284
rect 337102 273232 337108 273284
rect 337160 273232 337166 273284
rect 301056 273204 301084 273232
rect 301130 273204 301136 273216
rect 301056 273176 301136 273204
rect 301130 273164 301136 273176
rect 301188 273164 301194 273216
rect 337120 273136 337148 273232
rect 358998 273164 359004 273216
rect 359056 273204 359062 273216
rect 359182 273204 359188 273216
rect 359056 273176 359188 273204
rect 359056 273164 359062 273176
rect 359182 273164 359188 273176
rect 359240 273164 359246 273216
rect 337194 273136 337200 273148
rect 337120 273108 337200 273136
rect 337194 273096 337200 273108
rect 337252 273096 337258 273148
rect 357434 272552 357440 272604
rect 357492 272592 357498 272604
rect 357894 272592 357900 272604
rect 357492 272564 357900 272592
rect 357492 272552 357498 272564
rect 357894 272552 357900 272564
rect 357952 272552 357958 272604
rect 294230 270580 294236 270632
rect 294288 270580 294294 270632
rect 232222 270552 232228 270564
rect 232183 270524 232228 270552
rect 232222 270512 232228 270524
rect 232280 270512 232286 270564
rect 251174 270512 251180 270564
rect 251232 270552 251238 270564
rect 251450 270552 251456 270564
rect 251232 270524 251456 270552
rect 251232 270512 251238 270524
rect 251450 270512 251456 270524
rect 251508 270512 251514 270564
rect 273533 270555 273591 270561
rect 273533 270521 273545 270555
rect 273579 270552 273591 270555
rect 273622 270552 273628 270564
rect 273579 270524 273628 270552
rect 273579 270521 273591 270524
rect 273533 270515 273591 270521
rect 273622 270512 273628 270524
rect 273680 270512 273686 270564
rect 294138 270444 294144 270496
rect 294196 270484 294202 270496
rect 294248 270484 294276 270580
rect 372706 270552 372712 270564
rect 372667 270524 372712 270552
rect 372706 270512 372712 270524
rect 372764 270512 372770 270564
rect 375834 270552 375840 270564
rect 375795 270524 375840 270552
rect 375834 270512 375840 270524
rect 375892 270512 375898 270564
rect 377122 270552 377128 270564
rect 377083 270524 377128 270552
rect 377122 270512 377128 270524
rect 377180 270512 377186 270564
rect 424597 270555 424655 270561
rect 424597 270521 424609 270555
rect 424643 270552 424655 270555
rect 424778 270552 424784 270564
rect 424643 270524 424784 270552
rect 424643 270521 424655 270524
rect 424597 270515 424655 270521
rect 424778 270512 424784 270524
rect 424836 270512 424842 270564
rect 294196 270456 294276 270484
rect 294196 270444 294202 270456
rect 301130 270444 301136 270496
rect 301188 270484 301194 270496
rect 301222 270484 301228 270496
rect 301188 270456 301228 270484
rect 301188 270444 301194 270456
rect 301222 270444 301228 270456
rect 301280 270444 301286 270496
rect 327258 270444 327264 270496
rect 327316 270484 327322 270496
rect 327350 270484 327356 270496
rect 327316 270456 327356 270484
rect 327316 270444 327322 270456
rect 327350 270444 327356 270456
rect 327408 270444 327414 270496
rect 341153 270487 341211 270493
rect 341153 270453 341165 270487
rect 341199 270484 341211 270487
rect 341242 270484 341248 270496
rect 341199 270456 341248 270484
rect 341199 270453 341211 270456
rect 341153 270447 341211 270453
rect 341242 270444 341248 270456
rect 341300 270444 341306 270496
rect 367002 270484 367008 270496
rect 366963 270456 367008 270484
rect 367002 270444 367008 270456
rect 367060 270444 367066 270496
rect 389361 270487 389419 270493
rect 389361 270453 389373 270487
rect 389407 270484 389419 270487
rect 389450 270484 389456 270496
rect 389407 270456 389456 270484
rect 389407 270453 389419 270456
rect 389361 270447 389419 270453
rect 389450 270444 389456 270456
rect 389508 270444 389514 270496
rect 470594 270484 470600 270496
rect 470555 270456 470600 270484
rect 470594 270444 470600 270456
rect 470652 270444 470658 270496
rect 232222 269124 232228 269136
rect 232183 269096 232228 269124
rect 232222 269084 232228 269096
rect 232280 269084 232286 269136
rect 250070 269084 250076 269136
rect 250128 269124 250134 269136
rect 250254 269124 250260 269136
rect 250128 269096 250260 269124
rect 250128 269084 250134 269096
rect 250254 269084 250260 269096
rect 250312 269084 250318 269136
rect 262582 269084 262588 269136
rect 262640 269124 262646 269136
rect 262674 269124 262680 269136
rect 262640 269096 262680 269124
rect 262640 269084 262646 269096
rect 262674 269084 262680 269096
rect 262732 269084 262738 269136
rect 284570 269084 284576 269136
rect 284628 269124 284634 269136
rect 284754 269124 284760 269136
rect 284628 269096 284760 269124
rect 284628 269084 284634 269096
rect 284754 269084 284760 269096
rect 284812 269084 284818 269136
rect 288802 269084 288808 269136
rect 288860 269124 288866 269136
rect 288894 269124 288900 269136
rect 288860 269096 288900 269124
rect 288860 269084 288866 269096
rect 288894 269084 288900 269096
rect 288952 269084 288958 269136
rect 324501 269127 324559 269133
rect 324501 269093 324513 269127
rect 324547 269124 324559 269127
rect 324590 269124 324596 269136
rect 324547 269096 324596 269124
rect 324547 269093 324559 269096
rect 324501 269087 324559 269093
rect 324590 269084 324596 269096
rect 324648 269084 324654 269136
rect 421190 269084 421196 269136
rect 421248 269124 421254 269136
rect 421374 269124 421380 269136
rect 421248 269096 421380 269124
rect 421248 269084 421254 269096
rect 421374 269084 421380 269096
rect 421432 269084 421438 269136
rect 267826 267724 267832 267776
rect 267884 267764 267890 267776
rect 268010 267764 268016 267776
rect 267884 267736 268016 267764
rect 267884 267724 267890 267736
rect 268010 267724 268016 267736
rect 268068 267724 268074 267776
rect 299658 267724 299664 267776
rect 299716 267764 299722 267776
rect 299842 267764 299848 267776
rect 299716 267736 299848 267764
rect 299716 267724 299722 267736
rect 299842 267724 299848 267736
rect 299900 267724 299906 267776
rect 463694 267724 463700 267776
rect 463752 267764 463758 267776
rect 463878 267764 463884 267776
rect 463752 267736 463884 267764
rect 463752 267724 463758 267736
rect 463878 267724 463884 267736
rect 463936 267724 463942 267776
rect 325970 263684 325976 263696
rect 325896 263656 325976 263684
rect 236270 263576 236276 263628
rect 236328 263576 236334 263628
rect 239122 263576 239128 263628
rect 239180 263576 239186 263628
rect 270678 263576 270684 263628
rect 270736 263576 270742 263628
rect 236288 263480 236316 263576
rect 236454 263480 236460 263492
rect 236288 263452 236460 263480
rect 236454 263440 236460 263452
rect 236512 263440 236518 263492
rect 239140 263480 239168 263576
rect 270696 263492 270724 263576
rect 325896 263560 325924 263656
rect 325970 263644 325976 263656
rect 326028 263644 326034 263696
rect 337102 263616 337108 263628
rect 337063 263588 337108 263616
rect 337102 263576 337108 263588
rect 337160 263576 337166 263628
rect 339678 263576 339684 263628
rect 339736 263616 339742 263628
rect 339862 263616 339868 263628
rect 339736 263588 339868 263616
rect 339736 263576 339742 263588
rect 339862 263576 339868 263588
rect 339920 263576 339926 263628
rect 360286 263576 360292 263628
rect 360344 263616 360350 263628
rect 360470 263616 360476 263628
rect 360344 263588 360476 263616
rect 360344 263576 360350 263588
rect 360470 263576 360476 263588
rect 360528 263576 360534 263628
rect 325878 263508 325884 263560
rect 325936 263508 325942 263560
rect 239214 263480 239220 263492
rect 239140 263452 239220 263480
rect 239214 263440 239220 263452
rect 239272 263440 239278 263492
rect 270678 263440 270684 263492
rect 270736 263440 270742 263492
rect 310882 263480 310888 263492
rect 310843 263452 310888 263480
rect 310882 263440 310888 263452
rect 310940 263440 310946 263492
rect 362218 263480 362224 263492
rect 362179 263452 362224 263480
rect 362218 263440 362224 263452
rect 362276 263440 362282 263492
rect 330110 263208 330116 263220
rect 330071 263180 330116 263208
rect 330110 263168 330116 263180
rect 330168 263168 330174 263220
rect 264974 262896 264980 262948
rect 265032 262936 265038 262948
rect 265158 262936 265164 262948
rect 265032 262908 265164 262936
rect 265032 262896 265038 262908
rect 265158 262896 265164 262908
rect 265216 262896 265222 262948
rect 306834 262936 306840 262948
rect 306795 262908 306840 262936
rect 306834 262896 306840 262908
rect 306892 262896 306898 262948
rect 272334 260964 272340 260976
rect 272168 260936 272340 260964
rect 232222 260856 232228 260908
rect 232280 260896 232286 260908
rect 232314 260896 232320 260908
rect 232280 260868 232320 260896
rect 232280 260856 232286 260868
rect 232314 260856 232320 260868
rect 232372 260856 232378 260908
rect 250070 260856 250076 260908
rect 250128 260896 250134 260908
rect 250162 260896 250168 260908
rect 250128 260868 250168 260896
rect 250128 260856 250134 260868
rect 250162 260856 250168 260868
rect 250220 260856 250226 260908
rect 266722 260856 266728 260908
rect 266780 260856 266786 260908
rect 266740 260772 266768 260856
rect 270678 260828 270684 260840
rect 270639 260800 270684 260828
rect 270678 260788 270684 260800
rect 270736 260788 270742 260840
rect 272168 260772 272196 260936
rect 272334 260924 272340 260936
rect 272392 260924 272398 260976
rect 284570 260856 284576 260908
rect 284628 260896 284634 260908
rect 284754 260896 284760 260908
rect 284628 260868 284760 260896
rect 284628 260856 284634 260868
rect 284754 260856 284760 260868
rect 284812 260856 284818 260908
rect 341150 260896 341156 260908
rect 341111 260868 341156 260896
rect 341150 260856 341156 260868
rect 341208 260856 341214 260908
rect 359090 260856 359096 260908
rect 359148 260896 359154 260908
rect 359182 260896 359188 260908
rect 359148 260868 359188 260896
rect 359148 260856 359154 260868
rect 359182 260856 359188 260868
rect 359240 260856 359246 260908
rect 367002 260896 367008 260908
rect 366963 260868 367008 260896
rect 367002 260856 367008 260868
rect 367060 260856 367066 260908
rect 389358 260896 389364 260908
rect 389319 260868 389364 260896
rect 389358 260856 389364 260868
rect 389416 260856 389422 260908
rect 470594 260896 470600 260908
rect 470555 260868 470600 260896
rect 470594 260856 470600 260868
rect 470652 260856 470658 260908
rect 273530 260828 273536 260840
rect 273491 260800 273536 260828
rect 273530 260788 273536 260800
rect 273588 260788 273594 260840
rect 324590 260788 324596 260840
rect 324648 260788 324654 260840
rect 372706 260828 372712 260840
rect 372667 260800 372712 260828
rect 372706 260788 372712 260800
rect 372764 260788 372770 260840
rect 375834 260828 375840 260840
rect 375795 260800 375840 260828
rect 375834 260788 375840 260800
rect 375892 260788 375898 260840
rect 377122 260828 377128 260840
rect 377083 260800 377128 260828
rect 377122 260788 377128 260800
rect 377180 260788 377186 260840
rect 424505 260831 424563 260837
rect 424505 260797 424517 260831
rect 424551 260828 424563 260831
rect 424594 260828 424600 260840
rect 424551 260800 424600 260828
rect 424551 260797 424563 260800
rect 424505 260791 424563 260797
rect 424594 260788 424600 260800
rect 424652 260788 424658 260840
rect 463697 260831 463755 260837
rect 463697 260797 463709 260831
rect 463743 260828 463755 260831
rect 463786 260828 463792 260840
rect 463743 260800 463792 260828
rect 463743 260797 463755 260800
rect 463697 260791 463755 260797
rect 463786 260788 463792 260800
rect 463844 260788 463850 260840
rect 266722 260720 266728 260772
rect 266780 260720 266786 260772
rect 272150 260720 272156 260772
rect 272208 260720 272214 260772
rect 324608 260760 324636 260788
rect 324682 260760 324688 260772
rect 324608 260732 324688 260760
rect 324682 260720 324688 260732
rect 324740 260720 324746 260772
rect 267734 259428 267740 259480
rect 267792 259468 267798 259480
rect 267826 259468 267832 259480
rect 267792 259440 267832 259468
rect 267792 259428 267798 259440
rect 267826 259428 267832 259440
rect 267884 259428 267890 259480
rect 296990 259428 296996 259480
rect 297048 259468 297054 259480
rect 297082 259468 297088 259480
rect 297048 259440 297088 259468
rect 297048 259428 297054 259440
rect 297082 259428 297088 259440
rect 297140 259428 297146 259480
rect 337102 259468 337108 259480
rect 337063 259440 337108 259468
rect 337102 259428 337108 259440
rect 337160 259428 337166 259480
rect 299842 259360 299848 259412
rect 299900 259400 299906 259412
rect 300026 259400 300032 259412
rect 299900 259372 300032 259400
rect 299900 259360 299906 259372
rect 300026 259360 300032 259372
rect 300084 259360 300090 259412
rect 330110 259360 330116 259412
rect 330168 259400 330174 259412
rect 330202 259400 330208 259412
rect 330168 259372 330208 259400
rect 330168 259360 330174 259372
rect 330202 259360 330208 259372
rect 330260 259360 330266 259412
rect 251174 259020 251180 259072
rect 251232 259060 251238 259072
rect 251358 259060 251364 259072
rect 251232 259032 251364 259060
rect 251232 259020 251238 259032
rect 251358 259020 251364 259032
rect 251416 259020 251422 259072
rect 288802 258000 288808 258052
rect 288860 258040 288866 258052
rect 288986 258040 288992 258052
rect 288860 258012 288992 258040
rect 288860 258000 288866 258012
rect 288986 258000 288992 258012
rect 289044 258000 289050 258052
rect 290001 258043 290059 258049
rect 290001 258009 290013 258043
rect 290047 258040 290059 258043
rect 290090 258040 290096 258052
rect 290047 258012 290096 258040
rect 290047 258009 290059 258012
rect 290001 258003 290059 258009
rect 290090 258000 290096 258012
rect 290148 258000 290154 258052
rect 294230 258040 294236 258052
rect 294191 258012 294236 258040
rect 294230 258000 294236 258012
rect 294288 258000 294294 258052
rect 296990 258000 296996 258052
rect 297048 258040 297054 258052
rect 297174 258040 297180 258052
rect 297048 258012 297180 258040
rect 297048 258000 297054 258012
rect 297174 258000 297180 258012
rect 297232 258000 297238 258052
rect 330202 258000 330208 258052
rect 330260 258040 330266 258052
rect 330386 258040 330392 258052
rect 330260 258012 330392 258040
rect 330260 258000 330266 258012
rect 330386 258000 330392 258012
rect 330444 258000 330450 258052
rect 245838 257932 245844 257984
rect 245896 257972 245902 257984
rect 245930 257972 245936 257984
rect 245896 257944 245936 257972
rect 245896 257932 245902 257944
rect 245930 257932 245936 257944
rect 245988 257932 245994 257984
rect 310882 256068 310888 256080
rect 310843 256040 310888 256068
rect 310882 256028 310888 256040
rect 310940 256028 310946 256080
rect 270678 256000 270684 256012
rect 270639 255972 270684 256000
rect 270678 255960 270684 255972
rect 270736 255960 270742 256012
rect 336734 254600 336740 254652
rect 336792 254640 336798 254652
rect 337102 254640 337108 254652
rect 336792 254612 337108 254640
rect 336792 254600 336798 254612
rect 337102 254600 337108 254612
rect 337160 254600 337166 254652
rect 236270 253920 236276 253972
rect 236328 253960 236334 253972
rect 236454 253960 236460 253972
rect 236328 253932 236460 253960
rect 236328 253920 236334 253932
rect 236454 253920 236460 253932
rect 236512 253920 236518 253972
rect 239030 253920 239036 253972
rect 239088 253960 239094 253972
rect 239214 253960 239220 253972
rect 239088 253932 239220 253960
rect 239088 253920 239094 253932
rect 239214 253920 239220 253932
rect 239272 253920 239278 253972
rect 250070 253960 250076 253972
rect 250031 253932 250076 253960
rect 250070 253920 250076 253932
rect 250128 253920 250134 253972
rect 362310 253960 362316 253972
rect 362236 253932 362316 253960
rect 362236 253904 362264 253932
rect 362310 253920 362316 253932
rect 362368 253920 362374 253972
rect 357526 253852 357532 253904
rect 357584 253892 357590 253904
rect 357710 253892 357716 253904
rect 357584 253864 357716 253892
rect 357584 253852 357590 253864
rect 357710 253852 357716 253864
rect 357768 253852 357774 253904
rect 358998 253852 359004 253904
rect 359056 253892 359062 253904
rect 359182 253892 359188 253904
rect 359056 253864 359188 253892
rect 359056 253852 359062 253864
rect 359182 253852 359188 253864
rect 359240 253852 359246 253904
rect 362218 253852 362224 253904
rect 362276 253852 362282 253904
rect 323394 252736 323400 252748
rect 323355 252708 323400 252736
rect 323394 252696 323400 252708
rect 323452 252696 323458 252748
rect 2774 252492 2780 252544
rect 2832 252532 2838 252544
rect 5258 252532 5264 252544
rect 2832 252504 5264 252532
rect 2832 252492 2838 252504
rect 5258 252492 5264 252504
rect 5316 252492 5322 252544
rect 469858 252492 469864 252544
rect 469916 252532 469922 252544
rect 580166 252532 580172 252544
rect 469916 252504 580172 252532
rect 469916 252492 469922 252504
rect 580166 252492 580172 252504
rect 580224 252492 580230 252544
rect 232314 251308 232320 251320
rect 232240 251280 232320 251308
rect 232240 251116 232268 251280
rect 232314 251268 232320 251280
rect 232372 251268 232378 251320
rect 310698 251268 310704 251320
rect 310756 251308 310762 251320
rect 310885 251311 310943 251317
rect 310885 251308 310897 251311
rect 310756 251280 310897 251308
rect 310756 251268 310762 251280
rect 310885 251277 310897 251280
rect 310931 251277 310943 251311
rect 310885 251271 310943 251277
rect 265158 251200 265164 251252
rect 265216 251240 265222 251252
rect 265250 251240 265256 251252
rect 265216 251212 265256 251240
rect 265216 251200 265222 251212
rect 265250 251200 265256 251212
rect 265308 251200 265314 251252
rect 267734 251200 267740 251252
rect 267792 251240 267798 251252
rect 267826 251240 267832 251252
rect 267792 251212 267832 251240
rect 267792 251200 267798 251212
rect 267826 251200 267832 251212
rect 267884 251200 267890 251252
rect 273533 251243 273591 251249
rect 273533 251209 273545 251243
rect 273579 251240 273591 251243
rect 273622 251240 273628 251252
rect 273579 251212 273628 251240
rect 273579 251209 273591 251212
rect 273533 251203 273591 251209
rect 273622 251200 273628 251212
rect 273680 251200 273686 251252
rect 291470 251200 291476 251252
rect 291528 251240 291534 251252
rect 291562 251240 291568 251252
rect 291528 251212 291568 251240
rect 291528 251200 291534 251212
rect 291562 251200 291568 251212
rect 291620 251200 291626 251252
rect 372706 251240 372712 251252
rect 372667 251212 372712 251240
rect 372706 251200 372712 251212
rect 372764 251200 372770 251252
rect 375834 251240 375840 251252
rect 375795 251212 375840 251240
rect 375834 251200 375840 251212
rect 375892 251200 375898 251252
rect 377122 251240 377128 251252
rect 377083 251212 377128 251240
rect 377122 251200 377128 251212
rect 377180 251200 377186 251252
rect 389174 251200 389180 251252
rect 389232 251240 389238 251252
rect 389358 251240 389364 251252
rect 389232 251212 389364 251240
rect 389232 251200 389238 251212
rect 389358 251200 389364 251212
rect 389416 251200 389422 251252
rect 424502 251240 424508 251252
rect 424463 251212 424508 251240
rect 424502 251200 424508 251212
rect 424560 251200 424566 251252
rect 463694 251200 463700 251252
rect 463752 251240 463758 251252
rect 463752 251212 463797 251240
rect 463752 251200 463758 251212
rect 239122 251132 239128 251184
rect 239180 251172 239186 251184
rect 239214 251172 239220 251184
rect 239180 251144 239220 251172
rect 239180 251132 239186 251144
rect 239214 251132 239220 251144
rect 239272 251132 239278 251184
rect 259641 251175 259699 251181
rect 259641 251141 259653 251175
rect 259687 251172 259699 251175
rect 259730 251172 259736 251184
rect 259687 251144 259736 251172
rect 259687 251141 259699 251144
rect 259641 251135 259699 251141
rect 259730 251132 259736 251144
rect 259788 251132 259794 251184
rect 262674 251132 262680 251184
rect 262732 251172 262738 251184
rect 262766 251172 262772 251184
rect 262732 251144 262772 251172
rect 262732 251132 262738 251144
rect 262766 251132 262772 251144
rect 262824 251132 262830 251184
rect 266722 251132 266728 251184
rect 266780 251132 266786 251184
rect 295518 251132 295524 251184
rect 295576 251172 295582 251184
rect 295702 251172 295708 251184
rect 295576 251144 295708 251172
rect 295576 251132 295582 251144
rect 295702 251132 295708 251144
rect 295760 251132 295766 251184
rect 310698 251172 310704 251184
rect 310659 251144 310704 251172
rect 310698 251132 310704 251144
rect 310756 251132 310762 251184
rect 325878 251172 325884 251184
rect 325839 251144 325884 251172
rect 325878 251132 325884 251144
rect 325936 251132 325942 251184
rect 357618 251132 357624 251184
rect 357676 251172 357682 251184
rect 357710 251172 357716 251184
rect 357676 251144 357716 251172
rect 357676 251132 357682 251144
rect 357710 251132 357716 251144
rect 357768 251132 357774 251184
rect 367002 251172 367008 251184
rect 366963 251144 367008 251172
rect 367002 251132 367008 251144
rect 367060 251132 367066 251184
rect 470594 251172 470600 251184
rect 470555 251144 470600 251172
rect 470594 251132 470600 251144
rect 470652 251132 470658 251184
rect 232222 251064 232228 251116
rect 232280 251064 232286 251116
rect 266740 251048 266768 251132
rect 266722 250996 266728 251048
rect 266780 250996 266786 251048
rect 327350 249948 327356 249960
rect 327184 249920 327356 249948
rect 327184 249892 327212 249920
rect 327350 249908 327356 249920
rect 327408 249908 327414 249960
rect 284662 249840 284668 249892
rect 284720 249880 284726 249892
rect 284754 249880 284760 249892
rect 284720 249852 284760 249880
rect 284720 249840 284726 249852
rect 284754 249840 284760 249852
rect 284812 249840 284818 249892
rect 324590 249840 324596 249892
rect 324648 249880 324654 249892
rect 324682 249880 324688 249892
rect 324648 249852 324688 249880
rect 324648 249840 324654 249852
rect 324682 249840 324688 249852
rect 324740 249840 324746 249892
rect 327166 249840 327172 249892
rect 327224 249840 327230 249892
rect 250070 249812 250076 249824
rect 250031 249784 250076 249812
rect 250070 249772 250076 249784
rect 250128 249772 250134 249824
rect 285950 249772 285956 249824
rect 286008 249812 286014 249824
rect 286042 249812 286048 249824
rect 286008 249784 286048 249812
rect 286008 249772 286014 249784
rect 286042 249772 286048 249784
rect 286100 249772 286106 249824
rect 306837 249815 306895 249821
rect 306837 249781 306849 249815
rect 306883 249812 306895 249815
rect 306926 249812 306932 249824
rect 306883 249784 306932 249812
rect 306883 249781 306895 249784
rect 306837 249775 306895 249781
rect 306926 249772 306932 249784
rect 306984 249772 306990 249824
rect 325878 249812 325884 249824
rect 325839 249784 325884 249812
rect 325878 249772 325884 249784
rect 325936 249772 325942 249824
rect 358538 249772 358544 249824
rect 358596 249812 358602 249824
rect 358722 249812 358728 249824
rect 358596 249784 358728 249812
rect 358596 249772 358602 249784
rect 358722 249772 358728 249784
rect 358780 249772 358786 249824
rect 421190 249772 421196 249824
rect 421248 249812 421254 249824
rect 421374 249812 421380 249824
rect 421248 249784 421380 249812
rect 421248 249772 421254 249784
rect 421374 249772 421380 249784
rect 421432 249772 421438 249824
rect 284662 249744 284668 249756
rect 284623 249716 284668 249744
rect 284662 249704 284668 249716
rect 284720 249704 284726 249756
rect 327166 249744 327172 249756
rect 327127 249716 327172 249744
rect 327166 249704 327172 249716
rect 327224 249704 327230 249756
rect 289998 248452 290004 248464
rect 289959 248424 290004 248452
rect 289998 248412 290004 248424
rect 290056 248412 290062 248464
rect 294230 248452 294236 248464
rect 294191 248424 294236 248452
rect 294230 248412 294236 248424
rect 294288 248412 294294 248464
rect 291470 248384 291476 248396
rect 291431 248356 291476 248384
rect 291470 248344 291476 248356
rect 291528 248344 291534 248396
rect 289998 245828 290004 245880
rect 290056 245868 290062 245880
rect 290366 245868 290372 245880
rect 290056 245840 290372 245868
rect 290056 245828 290062 245840
rect 290366 245828 290372 245840
rect 290424 245828 290430 245880
rect 285950 244984 285956 244996
rect 285911 244956 285956 244984
rect 285950 244944 285956 244956
rect 286008 244944 286014 244996
rect 272150 244332 272156 244384
rect 272208 244332 272214 244384
rect 341242 244372 341248 244384
rect 341168 244344 341248 244372
rect 236270 244264 236276 244316
rect 236328 244264 236334 244316
rect 270678 244304 270684 244316
rect 270639 244276 270684 244304
rect 270678 244264 270684 244276
rect 270736 244264 270742 244316
rect 236288 244168 236316 244264
rect 272168 244248 272196 244332
rect 339678 244264 339684 244316
rect 339736 244304 339742 244316
rect 339862 244304 339868 244316
rect 339736 244276 339868 244304
rect 339736 244264 339742 244276
rect 339862 244264 339868 244276
rect 339920 244264 339926 244316
rect 341168 244248 341196 244344
rect 341242 244332 341248 244344
rect 341300 244332 341306 244384
rect 360286 244264 360292 244316
rect 360344 244304 360350 244316
rect 360470 244304 360476 244316
rect 360344 244276 360476 244304
rect 360344 244264 360350 244276
rect 360470 244264 360476 244276
rect 360528 244264 360534 244316
rect 272150 244196 272156 244248
rect 272208 244196 272214 244248
rect 341150 244196 341156 244248
rect 341208 244196 341214 244248
rect 236454 244168 236460 244180
rect 236288 244140 236460 244168
rect 236454 244128 236460 244140
rect 236512 244128 236518 244180
rect 259638 242672 259644 242684
rect 259599 242644 259644 242672
rect 259638 242632 259644 242644
rect 259696 242632 259702 242684
rect 358722 241612 358728 241664
rect 358780 241612 358786 241664
rect 270678 241584 270684 241596
rect 270639 241556 270684 241584
rect 270678 241544 270684 241556
rect 270736 241544 270742 241596
rect 358740 241528 358768 241612
rect 388990 241544 388996 241596
rect 389048 241584 389054 241596
rect 389266 241584 389272 241596
rect 389048 241556 389272 241584
rect 389048 241544 389054 241556
rect 389266 241544 389272 241556
rect 389324 241544 389330 241596
rect 250070 241476 250076 241528
rect 250128 241516 250134 241528
rect 250162 241516 250168 241528
rect 250128 241488 250168 241516
rect 250128 241476 250134 241488
rect 250162 241476 250168 241488
rect 250220 241476 250226 241528
rect 251358 241516 251364 241528
rect 251319 241488 251364 241516
rect 251358 241476 251364 241488
rect 251416 241476 251422 241528
rect 310701 241519 310759 241525
rect 310701 241485 310713 241519
rect 310747 241516 310759 241519
rect 310882 241516 310888 241528
rect 310747 241488 310888 241516
rect 310747 241485 310759 241488
rect 310701 241479 310759 241485
rect 310882 241476 310888 241488
rect 310940 241476 310946 241528
rect 323394 241516 323400 241528
rect 323355 241488 323400 241516
rect 323394 241476 323400 241488
rect 323452 241476 323458 241528
rect 358722 241476 358728 241528
rect 358780 241476 358786 241528
rect 359090 241476 359096 241528
rect 359148 241516 359154 241528
rect 359182 241516 359188 241528
rect 359148 241488 359188 241516
rect 359148 241476 359154 241488
rect 359182 241476 359188 241488
rect 359240 241476 359246 241528
rect 367002 241516 367008 241528
rect 366963 241488 367008 241516
rect 367002 241476 367008 241488
rect 367060 241476 367066 241528
rect 470594 241516 470600 241528
rect 470555 241488 470600 241516
rect 470594 241476 470600 241488
rect 470652 241476 470658 241528
rect 270678 241448 270684 241460
rect 270639 241420 270684 241448
rect 270678 241408 270684 241420
rect 270736 241408 270742 241460
rect 299474 241408 299480 241460
rect 299532 241448 299538 241460
rect 362218 241448 362224 241460
rect 299532 241420 299577 241448
rect 362179 241420 362224 241448
rect 299532 241408 299538 241420
rect 362218 241408 362224 241420
rect 362276 241408 362282 241460
rect 375834 241448 375840 241460
rect 375795 241420 375840 241448
rect 375834 241408 375840 241420
rect 375892 241408 375898 241460
rect 389266 241448 389272 241460
rect 389227 241420 389272 241448
rect 389266 241408 389272 241420
rect 389324 241408 389330 241460
rect 327166 240224 327172 240236
rect 327127 240196 327172 240224
rect 327166 240184 327172 240196
rect 327224 240184 327230 240236
rect 232314 240116 232320 240168
rect 232372 240156 232378 240168
rect 232498 240156 232504 240168
rect 232372 240128 232504 240156
rect 232372 240116 232378 240128
rect 232498 240116 232504 240128
rect 232556 240116 232562 240168
rect 244366 240116 244372 240168
rect 244424 240156 244430 240168
rect 244458 240156 244464 240168
rect 244424 240128 244464 240156
rect 244424 240116 244430 240128
rect 244458 240116 244464 240128
rect 244516 240116 244522 240168
rect 245838 240116 245844 240168
rect 245896 240156 245902 240168
rect 245930 240156 245936 240168
rect 245896 240128 245936 240156
rect 245896 240116 245902 240128
rect 245930 240116 245936 240128
rect 245988 240116 245994 240168
rect 251358 240156 251364 240168
rect 251319 240128 251364 240156
rect 251358 240116 251364 240128
rect 251416 240116 251422 240168
rect 284665 240159 284723 240165
rect 284665 240125 284677 240159
rect 284711 240156 284723 240159
rect 284846 240156 284852 240168
rect 284711 240128 284852 240156
rect 284711 240125 284723 240128
rect 284665 240119 284723 240125
rect 284846 240116 284852 240128
rect 284904 240116 284910 240168
rect 299934 240116 299940 240168
rect 299992 240156 299998 240168
rect 300026 240156 300032 240168
rect 299992 240128 300032 240156
rect 299992 240116 299998 240128
rect 300026 240116 300032 240128
rect 300084 240116 300090 240168
rect 302418 240116 302424 240168
rect 302476 240156 302482 240168
rect 302694 240156 302700 240168
rect 302476 240128 302700 240156
rect 302476 240116 302482 240128
rect 302694 240116 302700 240128
rect 302752 240116 302758 240168
rect 306926 240116 306932 240168
rect 306984 240156 306990 240168
rect 307110 240156 307116 240168
rect 306984 240128 307116 240156
rect 306984 240116 306990 240128
rect 307110 240116 307116 240128
rect 307168 240116 307174 240168
rect 324590 240116 324596 240168
rect 324648 240156 324654 240168
rect 324682 240156 324688 240168
rect 324648 240128 324688 240156
rect 324648 240116 324654 240128
rect 324682 240116 324688 240128
rect 324740 240116 324746 240168
rect 325970 240116 325976 240168
rect 326028 240156 326034 240168
rect 326154 240156 326160 240168
rect 326028 240128 326160 240156
rect 326028 240116 326034 240128
rect 326154 240116 326160 240128
rect 326212 240116 326218 240168
rect 337102 240116 337108 240168
rect 337160 240156 337166 240168
rect 337286 240156 337292 240168
rect 337160 240128 337292 240156
rect 337160 240116 337166 240128
rect 337286 240116 337292 240128
rect 337344 240116 337350 240168
rect 291473 240091 291531 240097
rect 291473 240057 291485 240091
rect 291519 240088 291531 240091
rect 291746 240088 291752 240100
rect 291519 240060 291752 240088
rect 291519 240057 291531 240060
rect 291473 240051 291531 240057
rect 291746 240048 291752 240060
rect 291804 240048 291810 240100
rect 327166 240088 327172 240100
rect 327127 240060 327172 240088
rect 327166 240048 327172 240060
rect 327224 240048 327230 240100
rect 330110 240048 330116 240100
rect 330168 240088 330174 240100
rect 330202 240088 330208 240100
rect 330168 240060 330208 240088
rect 330168 240048 330174 240060
rect 330202 240048 330208 240060
rect 330260 240048 330266 240100
rect 330202 238688 330208 238740
rect 330260 238688 330266 238740
rect 330220 238660 330248 238688
rect 330386 238660 330392 238672
rect 330220 238632 330392 238660
rect 330386 238620 330392 238632
rect 330444 238620 330450 238672
rect 3050 237328 3056 237380
rect 3108 237368 3114 237380
rect 15838 237368 15844 237380
rect 3108 237340 15844 237368
rect 3108 237328 3114 237340
rect 15838 237328 15844 237340
rect 15896 237328 15902 237380
rect 244366 234852 244372 234864
rect 244327 234824 244372 234852
rect 244366 234812 244372 234824
rect 244424 234812 244430 234864
rect 310882 234716 310888 234728
rect 310808 234688 310888 234716
rect 250070 234608 250076 234660
rect 250128 234648 250134 234660
rect 250165 234651 250223 234657
rect 250165 234648 250177 234651
rect 250128 234620 250177 234648
rect 250128 234608 250134 234620
rect 250165 234617 250177 234620
rect 250211 234617 250223 234651
rect 250165 234611 250223 234617
rect 310808 234592 310836 234688
rect 310882 234676 310888 234688
rect 310940 234676 310946 234728
rect 323394 234716 323400 234728
rect 323355 234688 323400 234716
rect 323394 234676 323400 234688
rect 323452 234676 323458 234728
rect 389269 234651 389327 234657
rect 389269 234617 389281 234651
rect 389315 234648 389327 234651
rect 389450 234648 389456 234660
rect 389315 234620 389456 234648
rect 389315 234617 389327 234620
rect 389269 234611 389327 234617
rect 389450 234608 389456 234620
rect 389508 234608 389514 234660
rect 310790 234540 310796 234592
rect 310848 234540 310854 234592
rect 285950 234512 285956 234524
rect 285911 234484 285956 234512
rect 285950 234472 285956 234484
rect 286008 234472 286014 234524
rect 270678 232064 270684 232076
rect 270639 232036 270684 232064
rect 270678 232024 270684 232036
rect 270736 232024 270742 232076
rect 302605 231999 302663 232005
rect 302605 231965 302617 231999
rect 302651 231996 302663 231999
rect 302694 231996 302700 232008
rect 302651 231968 302700 231996
rect 302651 231965 302663 231968
rect 302605 231959 302663 231965
rect 302694 231956 302700 231968
rect 302752 231956 302758 232008
rect 236270 231888 236276 231940
rect 236328 231928 236334 231940
rect 236546 231928 236552 231940
rect 236328 231900 236552 231928
rect 236328 231888 236334 231900
rect 236546 231888 236552 231900
rect 236604 231888 236610 231940
rect 266722 231928 266728 231940
rect 266683 231900 266728 231928
rect 266722 231888 266728 231900
rect 266780 231888 266786 231940
rect 301130 231928 301136 231940
rect 301056 231900 301136 231928
rect 262674 231820 262680 231872
rect 262732 231860 262738 231872
rect 262766 231860 262772 231872
rect 262732 231832 262772 231860
rect 262732 231820 262738 231832
rect 262766 231820 262772 231832
rect 262824 231820 262830 231872
rect 265250 231820 265256 231872
rect 265308 231860 265314 231872
rect 265342 231860 265348 231872
rect 265308 231832 265348 231860
rect 265308 231820 265314 231832
rect 265342 231820 265348 231832
rect 265400 231820 265406 231872
rect 299474 231820 299480 231872
rect 299532 231860 299538 231872
rect 299532 231832 299577 231860
rect 299532 231820 299538 231832
rect 301056 231804 301084 231900
rect 301130 231888 301136 231900
rect 301188 231888 301194 231940
rect 366818 231888 366824 231940
rect 366876 231928 366882 231940
rect 367002 231928 367008 231940
rect 366876 231900 367008 231928
rect 366876 231888 366882 231900
rect 367002 231888 367008 231900
rect 367060 231888 367066 231940
rect 306926 231860 306932 231872
rect 306760 231832 306932 231860
rect 306760 231804 306788 231832
rect 306926 231820 306932 231832
rect 306984 231820 306990 231872
rect 357618 231820 357624 231872
rect 357676 231860 357682 231872
rect 357710 231860 357716 231872
rect 357676 231832 357716 231860
rect 357676 231820 357682 231832
rect 357710 231820 357716 231832
rect 357768 231820 357774 231872
rect 359090 231820 359096 231872
rect 359148 231860 359154 231872
rect 359182 231860 359188 231872
rect 359148 231832 359188 231860
rect 359148 231820 359154 231832
rect 359182 231820 359188 231832
rect 359240 231820 359246 231872
rect 372522 231820 372528 231872
rect 372580 231860 372586 231872
rect 372706 231860 372712 231872
rect 372580 231832 372712 231860
rect 372580 231820 372586 231832
rect 372706 231820 372712 231832
rect 372764 231820 372770 231872
rect 375834 231860 375840 231872
rect 375795 231832 375840 231860
rect 375834 231820 375840 231832
rect 375892 231820 375898 231872
rect 376938 231820 376944 231872
rect 376996 231860 377002 231872
rect 377122 231860 377128 231872
rect 376996 231832 377128 231860
rect 376996 231820 377002 231832
rect 377122 231820 377128 231832
rect 377180 231820 377186 231872
rect 301038 231752 301044 231804
rect 301096 231752 301102 231804
rect 306742 231752 306748 231804
rect 306800 231752 306806 231804
rect 310790 231792 310796 231804
rect 310751 231764 310796 231792
rect 310790 231752 310796 231764
rect 310848 231752 310854 231804
rect 323394 231792 323400 231804
rect 323355 231764 323400 231792
rect 323394 231752 323400 231764
rect 323452 231752 323458 231804
rect 324590 231752 324596 231804
rect 324648 231792 324654 231804
rect 324774 231792 324780 231804
rect 324648 231764 324780 231792
rect 324648 231752 324654 231764
rect 324774 231752 324780 231764
rect 324832 231752 324838 231804
rect 367002 231792 367008 231804
rect 366963 231764 367008 231792
rect 367002 231752 367008 231764
rect 367060 231752 367066 231804
rect 327166 230568 327172 230580
rect 327127 230540 327172 230568
rect 327166 230528 327172 230540
rect 327224 230528 327230 230580
rect 337010 230528 337016 230580
rect 337068 230568 337074 230580
rect 337194 230568 337200 230580
rect 337068 230540 337200 230568
rect 337068 230528 337074 230540
rect 337194 230528 337200 230540
rect 337252 230528 337258 230580
rect 244366 230500 244372 230512
rect 244327 230472 244372 230500
rect 244366 230460 244372 230472
rect 244424 230460 244430 230512
rect 245930 230460 245936 230512
rect 245988 230500 245994 230512
rect 246114 230500 246120 230512
rect 245988 230472 246120 230500
rect 245988 230460 245994 230472
rect 246114 230460 246120 230472
rect 246172 230460 246178 230512
rect 250162 230500 250168 230512
rect 250123 230472 250168 230500
rect 250162 230460 250168 230472
rect 250220 230460 250226 230512
rect 251082 230460 251088 230512
rect 251140 230500 251146 230512
rect 251358 230500 251364 230512
rect 251140 230472 251364 230500
rect 251140 230460 251146 230472
rect 251358 230460 251364 230472
rect 251416 230460 251422 230512
rect 259546 230460 259552 230512
rect 259604 230500 259610 230512
rect 259822 230500 259828 230512
rect 259604 230472 259828 230500
rect 259604 230460 259610 230472
rect 259822 230460 259828 230472
rect 259880 230460 259886 230512
rect 266722 230500 266728 230512
rect 266683 230472 266728 230500
rect 266722 230460 266728 230472
rect 266780 230460 266786 230512
rect 267918 230460 267924 230512
rect 267976 230500 267982 230512
rect 268102 230500 268108 230512
rect 267976 230472 268108 230500
rect 267976 230460 267982 230472
rect 268102 230460 268108 230472
rect 268160 230460 268166 230512
rect 302602 230500 302608 230512
rect 302563 230472 302608 230500
rect 302602 230460 302608 230472
rect 302660 230460 302666 230512
rect 341242 230460 341248 230512
rect 341300 230500 341306 230512
rect 341426 230500 341432 230512
rect 341300 230472 341432 230500
rect 341300 230460 341306 230472
rect 341426 230460 341432 230472
rect 341484 230460 341490 230512
rect 358538 230460 358544 230512
rect 358596 230500 358602 230512
rect 358722 230500 358728 230512
rect 358596 230472 358728 230500
rect 358596 230460 358602 230472
rect 358722 230460 358728 230472
rect 358780 230460 358786 230512
rect 362221 230503 362279 230509
rect 362221 230469 362233 230503
rect 362267 230500 362279 230503
rect 362402 230500 362408 230512
rect 362267 230472 362408 230500
rect 362267 230469 362279 230472
rect 362221 230463 362279 230469
rect 362402 230460 362408 230472
rect 362460 230460 362466 230512
rect 421190 230460 421196 230512
rect 421248 230500 421254 230512
rect 421374 230500 421380 230512
rect 421248 230472 421380 230500
rect 421248 230460 421254 230472
rect 421374 230460 421380 230472
rect 421432 230460 421438 230512
rect 244274 229032 244280 229084
rect 244332 229072 244338 229084
rect 244366 229072 244372 229084
rect 244332 229044 244372 229072
rect 244332 229032 244338 229044
rect 244366 229032 244372 229044
rect 244424 229032 244430 229084
rect 284846 225020 284852 225072
rect 284904 225020 284910 225072
rect 341242 225060 341248 225072
rect 341168 225032 341248 225060
rect 236270 224952 236276 225004
rect 236328 224952 236334 225004
rect 270678 224992 270684 225004
rect 270639 224964 270684 224992
rect 270678 224952 270684 224964
rect 270736 224952 270742 225004
rect 236288 224856 236316 224952
rect 284864 224936 284892 225020
rect 339678 224952 339684 225004
rect 339736 224992 339742 225004
rect 339862 224992 339868 225004
rect 339736 224964 339868 224992
rect 339736 224952 339742 224964
rect 339862 224952 339868 224964
rect 339920 224952 339926 225004
rect 341168 224936 341196 225032
rect 341242 225020 341248 225032
rect 341300 225020 341306 225072
rect 360286 224952 360292 225004
rect 360344 224992 360350 225004
rect 360470 224992 360476 225004
rect 360344 224964 360476 224992
rect 360344 224952 360350 224964
rect 360470 224952 360476 224964
rect 360528 224952 360534 225004
rect 284846 224884 284852 224936
rect 284904 224884 284910 224936
rect 341150 224884 341156 224936
rect 341208 224884 341214 224936
rect 236454 224856 236460 224868
rect 236288 224828 236460 224856
rect 236454 224816 236460 224828
rect 236512 224816 236518 224868
rect 329926 224204 329932 224256
rect 329984 224244 329990 224256
rect 330202 224244 330208 224256
rect 329984 224216 330208 224244
rect 329984 224204 329990 224216
rect 330202 224204 330208 224216
rect 330260 224204 330266 224256
rect 358722 222300 358728 222352
rect 358780 222300 358786 222352
rect 265250 222272 265256 222284
rect 265176 222244 265256 222272
rect 265176 222216 265204 222244
rect 265250 222232 265256 222244
rect 265308 222232 265314 222284
rect 270678 222272 270684 222284
rect 270639 222244 270684 222272
rect 270678 222232 270684 222244
rect 270736 222232 270742 222284
rect 358740 222216 358768 222300
rect 245838 222164 245844 222216
rect 245896 222204 245902 222216
rect 246022 222204 246028 222216
rect 245896 222176 246028 222204
rect 245896 222164 245902 222176
rect 246022 222164 246028 222176
rect 246080 222164 246086 222216
rect 265158 222164 265164 222216
rect 265216 222164 265222 222216
rect 295518 222164 295524 222216
rect 295576 222204 295582 222216
rect 295610 222204 295616 222216
rect 295576 222176 295616 222204
rect 295576 222164 295582 222176
rect 295610 222164 295616 222176
rect 295668 222164 295674 222216
rect 296806 222164 296812 222216
rect 296864 222204 296870 222216
rect 296898 222204 296904 222216
rect 296864 222176 296904 222204
rect 296864 222164 296870 222176
rect 296898 222164 296904 222176
rect 296956 222164 296962 222216
rect 306742 222164 306748 222216
rect 306800 222204 306806 222216
rect 306926 222204 306932 222216
rect 306800 222176 306932 222204
rect 306800 222164 306806 222176
rect 306926 222164 306932 222176
rect 306984 222164 306990 222216
rect 310793 222207 310851 222213
rect 310793 222173 310805 222207
rect 310839 222204 310851 222207
rect 310882 222204 310888 222216
rect 310839 222176 310888 222204
rect 310839 222173 310851 222176
rect 310793 222167 310851 222173
rect 310882 222164 310888 222176
rect 310940 222164 310946 222216
rect 358722 222164 358728 222216
rect 358780 222164 358786 222216
rect 362218 222164 362224 222216
rect 362276 222204 362282 222216
rect 362402 222204 362408 222216
rect 362276 222176 362408 222204
rect 362276 222164 362282 222176
rect 362402 222164 362408 222176
rect 362460 222164 362466 222216
rect 367002 222204 367008 222216
rect 366963 222176 367008 222204
rect 367002 222164 367008 222176
rect 367060 222164 367066 222216
rect 389266 222164 389272 222216
rect 389324 222204 389330 222216
rect 389542 222204 389548 222216
rect 389324 222176 389548 222204
rect 389324 222164 389330 222176
rect 389542 222164 389548 222176
rect 389600 222164 389606 222216
rect 463786 222164 463792 222216
rect 463844 222204 463850 222216
rect 464062 222204 464068 222216
rect 463844 222176 464068 222204
rect 463844 222164 463850 222176
rect 464062 222164 464068 222176
rect 464120 222164 464126 222216
rect 470410 222164 470416 222216
rect 470468 222204 470474 222216
rect 470594 222204 470600 222216
rect 470468 222176 470600 222204
rect 470468 222164 470474 222176
rect 470594 222164 470600 222176
rect 470652 222164 470658 222216
rect 270678 222136 270684 222148
rect 270639 222108 270684 222136
rect 270678 222096 270684 222108
rect 270736 222096 270742 222148
rect 299474 222096 299480 222148
rect 299532 222136 299538 222148
rect 375834 222136 375840 222148
rect 299532 222108 299577 222136
rect 375795 222108 375840 222136
rect 299532 222096 299538 222108
rect 375834 222096 375840 222108
rect 375892 222096 375898 222148
rect 337102 220872 337108 220924
rect 337160 220912 337166 220924
rect 337378 220912 337384 220924
rect 337160 220884 337384 220912
rect 337160 220872 337166 220884
rect 337378 220872 337384 220884
rect 337436 220872 337442 220924
rect 232314 220804 232320 220856
rect 232372 220844 232378 220856
rect 232498 220844 232504 220856
rect 232372 220816 232504 220844
rect 232372 220804 232378 220816
rect 232498 220804 232504 220816
rect 232556 220804 232562 220856
rect 251542 220804 251548 220856
rect 251600 220844 251606 220856
rect 251634 220844 251640 220856
rect 251600 220816 251640 220844
rect 251600 220804 251606 220816
rect 251634 220804 251640 220816
rect 251692 220804 251698 220856
rect 267734 220804 267740 220856
rect 267792 220844 267798 220856
rect 267918 220844 267924 220856
rect 267792 220816 267924 220844
rect 267792 220804 267798 220816
rect 267918 220804 267924 220816
rect 267976 220804 267982 220856
rect 290182 220804 290188 220856
rect 290240 220844 290246 220856
rect 290366 220844 290372 220856
rect 290240 220816 290372 220844
rect 290240 220804 290246 220816
rect 290366 220804 290372 220816
rect 290424 220804 290430 220856
rect 291654 220804 291660 220856
rect 291712 220844 291718 220856
rect 291838 220844 291844 220856
rect 291712 220816 291844 220844
rect 291712 220804 291718 220816
rect 291838 220804 291844 220816
rect 291896 220804 291902 220856
rect 294322 220804 294328 220856
rect 294380 220844 294386 220856
rect 294414 220844 294420 220856
rect 294380 220816 294420 220844
rect 294380 220804 294386 220816
rect 294414 220804 294420 220816
rect 294472 220804 294478 220856
rect 325878 220804 325884 220856
rect 325936 220844 325942 220856
rect 326062 220844 326068 220856
rect 325936 220816 326068 220844
rect 325936 220804 325942 220816
rect 326062 220804 326068 220816
rect 326120 220804 326126 220856
rect 327350 220804 327356 220856
rect 327408 220844 327414 220856
rect 327534 220844 327540 220856
rect 327408 220816 327540 220844
rect 327408 220804 327414 220816
rect 327534 220804 327540 220816
rect 327592 220804 327598 220856
rect 337102 220736 337108 220788
rect 337160 220776 337166 220788
rect 337286 220776 337292 220788
rect 337160 220748 337292 220776
rect 337160 220736 337166 220748
rect 337286 220736 337292 220748
rect 337344 220736 337350 220788
rect 341150 220776 341156 220788
rect 341111 220748 341156 220776
rect 341150 220736 341156 220748
rect 341208 220736 341214 220788
rect 244458 219376 244464 219428
rect 244516 219416 244522 219428
rect 244550 219416 244556 219428
rect 244516 219388 244556 219416
rect 244516 219376 244522 219388
rect 244550 219376 244556 219388
rect 244608 219376 244614 219428
rect 317506 219376 317512 219428
rect 317564 219416 317570 219428
rect 317690 219416 317696 219428
rect 317564 219388 317696 219416
rect 317564 219376 317570 219388
rect 317690 219376 317696 219388
rect 317748 219376 317754 219428
rect 330110 219416 330116 219428
rect 330071 219388 330116 219416
rect 330110 219376 330116 219388
rect 330168 219376 330174 219428
rect 244458 217988 244464 218000
rect 244419 217960 244464 217988
rect 244458 217948 244464 217960
rect 244516 217948 244522 218000
rect 310882 215404 310888 215416
rect 310808 215376 310888 215404
rect 310808 215280 310836 215376
rect 310882 215364 310888 215376
rect 310940 215364 310946 215416
rect 389542 215404 389548 215416
rect 389468 215376 389548 215404
rect 362129 215339 362187 215345
rect 362129 215305 362141 215339
rect 362175 215336 362187 215339
rect 362310 215336 362316 215348
rect 362175 215308 362316 215336
rect 362175 215305 362187 215308
rect 362129 215299 362187 215305
rect 362310 215296 362316 215308
rect 362368 215296 362374 215348
rect 389468 215280 389496 215376
rect 389542 215364 389548 215376
rect 389600 215364 389606 215416
rect 464062 215404 464068 215416
rect 463988 215376 464068 215404
rect 463988 215280 464016 215376
rect 464062 215364 464068 215376
rect 464120 215364 464126 215416
rect 310790 215228 310796 215280
rect 310848 215228 310854 215280
rect 341150 215268 341156 215280
rect 341111 215240 341156 215268
rect 341150 215228 341156 215240
rect 341208 215228 341214 215280
rect 357526 215228 357532 215280
rect 357584 215268 357590 215280
rect 357710 215268 357716 215280
rect 357584 215240 357716 215268
rect 357584 215228 357590 215240
rect 357710 215228 357716 215240
rect 357768 215228 357774 215280
rect 358998 215228 359004 215280
rect 359056 215268 359062 215280
rect 359182 215268 359188 215280
rect 359056 215240 359188 215268
rect 359056 215228 359062 215240
rect 359182 215228 359188 215240
rect 359240 215228 359246 215280
rect 389450 215228 389456 215280
rect 389508 215228 389514 215280
rect 463970 215228 463976 215280
rect 464028 215228 464034 215280
rect 270678 212752 270684 212764
rect 270639 212724 270684 212752
rect 270678 212712 270684 212724
rect 270736 212712 270742 212764
rect 236270 212576 236276 212628
rect 236328 212616 236334 212628
rect 236454 212616 236460 212628
rect 236328 212588 236460 212616
rect 236328 212576 236334 212588
rect 236454 212576 236460 212588
rect 236512 212576 236518 212628
rect 239122 212576 239128 212628
rect 239180 212616 239186 212628
rect 239398 212616 239404 212628
rect 239180 212588 239404 212616
rect 239180 212576 239186 212588
rect 239398 212576 239404 212588
rect 239456 212576 239462 212628
rect 290182 212576 290188 212628
rect 290240 212576 290246 212628
rect 291654 212576 291660 212628
rect 291712 212576 291718 212628
rect 301130 212616 301136 212628
rect 301056 212588 301136 212616
rect 245838 212508 245844 212560
rect 245896 212548 245902 212560
rect 245930 212548 245936 212560
rect 245896 212520 245936 212548
rect 245896 212508 245902 212520
rect 245930 212508 245936 212520
rect 245988 212508 245994 212560
rect 250070 212508 250076 212560
rect 250128 212548 250134 212560
rect 250254 212548 250260 212560
rect 250128 212520 250260 212548
rect 250128 212508 250134 212520
rect 250254 212508 250260 212520
rect 250312 212508 250318 212560
rect 265158 212508 265164 212560
rect 265216 212548 265222 212560
rect 265250 212548 265256 212560
rect 265216 212520 265256 212548
rect 265216 212508 265222 212520
rect 265250 212508 265256 212520
rect 265308 212508 265314 212560
rect 266630 212508 266636 212560
rect 266688 212548 266694 212560
rect 266814 212548 266820 212560
rect 266688 212520 266820 212548
rect 266688 212508 266694 212520
rect 266814 212508 266820 212520
rect 266872 212508 266878 212560
rect 267734 212508 267740 212560
rect 267792 212548 267798 212560
rect 267826 212548 267832 212560
rect 267792 212520 267832 212548
rect 267792 212508 267798 212520
rect 267826 212508 267832 212520
rect 267884 212508 267890 212560
rect 272150 212548 272156 212560
rect 272111 212520 272156 212548
rect 272150 212508 272156 212520
rect 272208 212508 272214 212560
rect 290200 212492 290228 212576
rect 291672 212492 291700 212576
rect 299474 212508 299480 212560
rect 299532 212548 299538 212560
rect 299532 212520 299577 212548
rect 299532 212508 299538 212520
rect 301056 212492 301084 212588
rect 301130 212576 301136 212588
rect 301188 212576 301194 212628
rect 306926 212616 306932 212628
rect 306760 212588 306932 212616
rect 306760 212492 306788 212588
rect 306926 212576 306932 212588
rect 306984 212576 306990 212628
rect 324682 212508 324688 212560
rect 324740 212548 324746 212560
rect 324774 212548 324780 212560
rect 324740 212520 324780 212548
rect 324740 212508 324746 212520
rect 324774 212508 324780 212520
rect 324832 212508 324838 212560
rect 325878 212508 325884 212560
rect 325936 212548 325942 212560
rect 325970 212548 325976 212560
rect 325936 212520 325976 212548
rect 325936 212508 325942 212520
rect 325970 212508 325976 212520
rect 326028 212508 326034 212560
rect 372522 212508 372528 212560
rect 372580 212548 372586 212560
rect 372706 212548 372712 212560
rect 372580 212520 372712 212548
rect 372580 212508 372586 212520
rect 372706 212508 372712 212520
rect 372764 212508 372770 212560
rect 375834 212548 375840 212560
rect 375795 212520 375840 212548
rect 375834 212508 375840 212520
rect 375892 212508 375898 212560
rect 376938 212508 376944 212560
rect 376996 212548 377002 212560
rect 377122 212548 377128 212560
rect 376996 212520 377128 212548
rect 376996 212508 377002 212520
rect 377122 212508 377128 212520
rect 377180 212508 377186 212560
rect 284662 212440 284668 212492
rect 284720 212480 284726 212492
rect 284846 212480 284852 212492
rect 284720 212452 284852 212480
rect 284720 212440 284726 212452
rect 284846 212440 284852 212452
rect 284904 212440 284910 212492
rect 290182 212440 290188 212492
rect 290240 212440 290246 212492
rect 291654 212440 291660 212492
rect 291712 212440 291718 212492
rect 301038 212440 301044 212492
rect 301096 212440 301102 212492
rect 306742 212440 306748 212492
rect 306800 212440 306806 212492
rect 310790 212480 310796 212492
rect 310751 212452 310796 212480
rect 310790 212440 310796 212452
rect 310848 212440 310854 212492
rect 232225 211259 232283 211265
rect 232225 211225 232237 211259
rect 232271 211256 232283 211259
rect 232314 211256 232320 211268
rect 232271 211228 232320 211256
rect 232271 211225 232283 211228
rect 232225 211219 232283 211225
rect 232314 211216 232320 211228
rect 232372 211216 232378 211268
rect 272150 211188 272156 211200
rect 272111 211160 272156 211188
rect 272150 211148 272156 211160
rect 272208 211148 272214 211200
rect 358538 211148 358544 211200
rect 358596 211188 358602 211200
rect 358630 211188 358636 211200
rect 358596 211160 358636 211188
rect 358596 211148 358602 211160
rect 358630 211148 358636 211160
rect 358688 211148 358694 211200
rect 362126 211188 362132 211200
rect 362087 211160 362132 211188
rect 362126 211148 362132 211160
rect 362184 211148 362190 211200
rect 239030 211080 239036 211132
rect 239088 211120 239094 211132
rect 239306 211120 239312 211132
rect 239088 211092 239312 211120
rect 239088 211080 239094 211092
rect 239306 211080 239312 211092
rect 239364 211080 239370 211132
rect 265250 211120 265256 211132
rect 265211 211092 265256 211120
rect 265250 211080 265256 211092
rect 265308 211080 265314 211132
rect 284662 211080 284668 211132
rect 284720 211120 284726 211132
rect 284938 211120 284944 211132
rect 284720 211092 284944 211120
rect 284720 211080 284726 211092
rect 284938 211080 284944 211092
rect 284996 211080 285002 211132
rect 294230 211080 294236 211132
rect 294288 211120 294294 211132
rect 294322 211120 294328 211132
rect 294288 211092 294328 211120
rect 294288 211080 294294 211092
rect 294322 211080 294328 211092
rect 294380 211080 294386 211132
rect 288802 210944 288808 210996
rect 288860 210984 288866 210996
rect 289170 210984 289176 210996
rect 288860 210956 289176 210984
rect 288860 210944 288866 210956
rect 289170 210944 289176 210956
rect 289228 210944 289234 210996
rect 232222 209828 232228 209840
rect 232183 209800 232228 209828
rect 232222 209788 232228 209800
rect 232280 209788 232286 209840
rect 317506 209788 317512 209840
rect 317564 209828 317570 209840
rect 317690 209828 317696 209840
rect 317564 209800 317696 209828
rect 317564 209788 317570 209800
rect 317690 209788 317696 209800
rect 317748 209788 317754 209840
rect 330110 209828 330116 209840
rect 330071 209800 330116 209828
rect 330110 209788 330116 209800
rect 330168 209788 330174 209840
rect 284662 209720 284668 209772
rect 284720 209760 284726 209772
rect 284754 209760 284760 209772
rect 284720 209732 284760 209760
rect 284720 209720 284726 209732
rect 284754 209720 284760 209732
rect 284812 209720 284818 209772
rect 330202 209760 330208 209772
rect 330163 209732 330208 209760
rect 330202 209720 330208 209732
rect 330260 209720 330266 209772
rect 250070 205640 250076 205692
rect 250128 205640 250134 205692
rect 323302 205640 323308 205692
rect 323360 205640 323366 205692
rect 339678 205640 339684 205692
rect 339736 205680 339742 205692
rect 339862 205680 339868 205692
rect 339736 205652 339868 205680
rect 339736 205640 339742 205652
rect 339862 205640 339868 205652
rect 339920 205640 339926 205692
rect 360286 205640 360292 205692
rect 360344 205680 360350 205692
rect 360470 205680 360476 205692
rect 360344 205652 360476 205680
rect 360344 205640 360350 205652
rect 360470 205640 360476 205652
rect 360528 205640 360534 205692
rect 250088 205612 250116 205640
rect 250162 205612 250168 205624
rect 250088 205584 250168 205612
rect 250162 205572 250168 205584
rect 250220 205572 250226 205624
rect 323320 205544 323348 205640
rect 323394 205544 323400 205556
rect 323320 205516 323400 205544
rect 323394 205504 323400 205516
rect 323452 205504 323458 205556
rect 245838 202852 245844 202904
rect 245896 202892 245902 202904
rect 245930 202892 245936 202904
rect 245896 202864 245936 202892
rect 245896 202852 245902 202864
rect 245930 202852 245936 202864
rect 245988 202852 245994 202904
rect 267734 202852 267740 202904
rect 267792 202892 267798 202904
rect 267826 202892 267832 202904
rect 267792 202864 267832 202892
rect 267792 202852 267798 202864
rect 267826 202852 267832 202864
rect 267884 202852 267890 202904
rect 285950 202852 285956 202904
rect 286008 202892 286014 202904
rect 286134 202892 286140 202904
rect 286008 202864 286140 202892
rect 286008 202852 286014 202864
rect 286134 202852 286140 202864
rect 286192 202852 286198 202904
rect 295518 202852 295524 202904
rect 295576 202892 295582 202904
rect 295610 202892 295616 202904
rect 295576 202864 295616 202892
rect 295576 202852 295582 202864
rect 295610 202852 295616 202864
rect 295668 202852 295674 202904
rect 296806 202852 296812 202904
rect 296864 202892 296870 202904
rect 296898 202892 296904 202904
rect 296864 202864 296904 202892
rect 296864 202852 296870 202864
rect 296898 202852 296904 202864
rect 296956 202852 296962 202904
rect 306742 202852 306748 202904
rect 306800 202892 306806 202904
rect 306926 202892 306932 202904
rect 306800 202864 306932 202892
rect 306800 202852 306806 202864
rect 306926 202852 306932 202864
rect 306984 202852 306990 202904
rect 310793 202895 310851 202901
rect 310793 202861 310805 202895
rect 310839 202892 310851 202895
rect 310882 202892 310888 202904
rect 310839 202864 310888 202892
rect 310839 202861 310851 202864
rect 310793 202855 310851 202861
rect 310882 202852 310888 202864
rect 310940 202852 310946 202904
rect 324590 202852 324596 202904
rect 324648 202892 324654 202904
rect 324682 202892 324688 202904
rect 324648 202864 324688 202892
rect 324648 202852 324654 202864
rect 324682 202852 324688 202864
rect 324740 202852 324746 202904
rect 325878 202852 325884 202904
rect 325936 202892 325942 202904
rect 325970 202892 325976 202904
rect 325936 202864 325976 202892
rect 325936 202852 325942 202864
rect 325970 202852 325976 202864
rect 326028 202852 326034 202904
rect 341150 202852 341156 202904
rect 341208 202892 341214 202904
rect 341242 202892 341248 202904
rect 341208 202864 341248 202892
rect 341208 202852 341214 202864
rect 341242 202852 341248 202864
rect 341300 202852 341306 202904
rect 358630 202852 358636 202904
rect 358688 202892 358694 202904
rect 358722 202892 358728 202904
rect 358688 202864 358728 202892
rect 358688 202852 358694 202864
rect 358722 202852 358728 202864
rect 358780 202852 358786 202904
rect 359090 202852 359096 202904
rect 359148 202892 359154 202904
rect 359182 202892 359188 202904
rect 359148 202864 359188 202892
rect 359148 202852 359154 202864
rect 359182 202852 359188 202864
rect 359240 202852 359246 202904
rect 362126 202852 362132 202904
rect 362184 202892 362190 202904
rect 362218 202892 362224 202904
rect 362184 202864 362224 202892
rect 362184 202852 362190 202864
rect 362218 202852 362224 202864
rect 362276 202852 362282 202904
rect 389266 202852 389272 202904
rect 389324 202892 389330 202904
rect 389542 202892 389548 202904
rect 389324 202864 389548 202892
rect 389324 202852 389330 202864
rect 389542 202852 389548 202864
rect 389600 202852 389606 202904
rect 421190 202852 421196 202904
rect 421248 202892 421254 202904
rect 421374 202892 421380 202904
rect 421248 202864 421380 202892
rect 421248 202852 421254 202864
rect 421374 202852 421380 202864
rect 421432 202852 421438 202904
rect 424594 202852 424600 202904
rect 424652 202892 424658 202904
rect 424870 202892 424876 202904
rect 424652 202864 424876 202892
rect 424652 202852 424658 202864
rect 424870 202852 424876 202864
rect 424928 202852 424934 202904
rect 463786 202852 463792 202904
rect 463844 202892 463850 202904
rect 464062 202892 464068 202904
rect 463844 202864 464068 202892
rect 463844 202852 463850 202864
rect 464062 202852 464068 202864
rect 464120 202852 464126 202904
rect 470410 202852 470416 202904
rect 470468 202892 470474 202904
rect 470594 202892 470600 202904
rect 470468 202864 470600 202892
rect 470468 202852 470474 202864
rect 470594 202852 470600 202864
rect 470652 202852 470658 202904
rect 299474 202784 299480 202836
rect 299532 202824 299538 202836
rect 299532 202796 299577 202824
rect 299532 202784 299538 202796
rect 330110 202784 330116 202836
rect 330168 202824 330174 202836
rect 330205 202827 330263 202833
rect 330205 202824 330217 202827
rect 330168 202796 330217 202824
rect 330168 202784 330174 202796
rect 330205 202793 330217 202796
rect 330251 202793 330263 202827
rect 336918 202824 336924 202836
rect 336879 202796 336924 202824
rect 330205 202787 330263 202793
rect 336918 202784 336924 202796
rect 336976 202784 336982 202836
rect 375834 202824 375840 202836
rect 375795 202796 375840 202824
rect 375834 202784 375840 202796
rect 375892 202784 375898 202836
rect 265250 202756 265256 202768
rect 265211 202728 265256 202756
rect 265250 202716 265256 202728
rect 265308 202716 265314 202768
rect 264974 201424 264980 201476
rect 265032 201464 265038 201476
rect 265250 201464 265256 201476
rect 265032 201436 265256 201464
rect 265032 201424 265038 201436
rect 265250 201424 265256 201436
rect 265308 201424 265314 201476
rect 266630 201424 266636 201476
rect 266688 201464 266694 201476
rect 266814 201464 266820 201476
rect 266688 201436 266820 201464
rect 266688 201424 266694 201436
rect 266814 201424 266820 201436
rect 266872 201424 266878 201476
rect 358633 201467 358691 201473
rect 358633 201433 358645 201467
rect 358679 201464 358691 201467
rect 358722 201464 358728 201476
rect 358679 201436 358728 201464
rect 358679 201433 358691 201436
rect 358633 201427 358691 201433
rect 358722 201424 358728 201436
rect 358780 201424 358786 201476
rect 421098 201424 421104 201476
rect 421156 201464 421162 201476
rect 421190 201464 421196 201476
rect 421156 201436 421196 201464
rect 421156 201424 421162 201436
rect 421190 201424 421196 201436
rect 421248 201424 421254 201476
rect 244458 200172 244464 200184
rect 244419 200144 244464 200172
rect 244458 200132 244464 200144
rect 244516 200132 244522 200184
rect 284662 200064 284668 200116
rect 284720 200104 284726 200116
rect 284846 200104 284852 200116
rect 284720 200076 284852 200104
rect 284720 200064 284726 200076
rect 284846 200064 284852 200076
rect 284904 200064 284910 200116
rect 291473 200107 291531 200113
rect 291473 200073 291485 200107
rect 291519 200104 291531 200107
rect 291654 200104 291660 200116
rect 291519 200076 291660 200104
rect 291519 200073 291531 200076
rect 291473 200067 291531 200073
rect 291654 200064 291660 200076
rect 291712 200064 291718 200116
rect 317506 200064 317512 200116
rect 317564 200104 317570 200116
rect 317690 200104 317696 200116
rect 317564 200076 317696 200104
rect 317564 200064 317570 200076
rect 317690 200064 317696 200076
rect 317748 200064 317754 200116
rect 284662 198676 284668 198688
rect 284623 198648 284668 198676
rect 284662 198636 284668 198648
rect 284720 198636 284726 198688
rect 285766 198024 285772 198076
rect 285824 198064 285830 198076
rect 285950 198064 285956 198076
rect 285824 198036 285956 198064
rect 285824 198024 285830 198036
rect 285950 198024 285956 198036
rect 286008 198024 286014 198076
rect 294230 198024 294236 198076
rect 294288 198064 294294 198076
rect 294414 198064 294420 198076
rect 294288 198036 294420 198064
rect 294288 198024 294294 198036
rect 294414 198024 294420 198036
rect 294472 198024 294478 198076
rect 362218 198064 362224 198076
rect 362179 198036 362224 198064
rect 362218 198024 362224 198036
rect 362276 198024 362282 198076
rect 289998 196596 290004 196648
rect 290056 196636 290062 196648
rect 290182 196636 290188 196648
rect 290056 196608 290188 196636
rect 290056 196596 290062 196608
rect 290182 196596 290188 196608
rect 290240 196596 290246 196648
rect 310882 196092 310888 196104
rect 310808 196064 310888 196092
rect 262582 195984 262588 196036
rect 262640 195984 262646 196036
rect 262600 195956 262628 195984
rect 310808 195968 310836 196064
rect 310882 196052 310888 196064
rect 310940 196052 310946 196104
rect 389542 196092 389548 196104
rect 389468 196064 389548 196092
rect 389468 195968 389496 196064
rect 389542 196052 389548 196064
rect 389600 196052 389606 196104
rect 464062 196092 464068 196104
rect 463988 196064 464068 196092
rect 424686 195984 424692 196036
rect 424744 196024 424750 196036
rect 424870 196024 424876 196036
rect 424744 195996 424876 196024
rect 424744 195984 424750 195996
rect 424870 195984 424876 195996
rect 424928 195984 424934 196036
rect 463988 195968 464016 196064
rect 464062 196052 464068 196064
rect 464120 196052 464126 196104
rect 262674 195956 262680 195968
rect 262600 195928 262680 195956
rect 262674 195916 262680 195928
rect 262732 195916 262738 195968
rect 310790 195916 310796 195968
rect 310848 195916 310854 195968
rect 389450 195916 389456 195968
rect 389508 195916 389514 195968
rect 463970 195916 463976 195968
rect 464028 195916 464034 195968
rect 236270 193332 236276 193384
rect 236328 193332 236334 193384
rect 245838 193332 245844 193384
rect 245896 193332 245902 193384
rect 236288 193248 236316 193332
rect 236270 193196 236276 193248
rect 236328 193196 236334 193248
rect 239122 193196 239128 193248
rect 239180 193236 239186 193248
rect 239214 193236 239220 193248
rect 239180 193208 239220 193236
rect 239180 193196 239186 193208
rect 239214 193196 239220 193208
rect 239272 193196 239278 193248
rect 245856 193180 245884 193332
rect 302694 193304 302700 193316
rect 302528 193276 302700 193304
rect 250070 193196 250076 193248
rect 250128 193236 250134 193248
rect 250254 193236 250260 193248
rect 250128 193208 250260 193236
rect 250128 193196 250134 193208
rect 250254 193196 250260 193208
rect 250312 193196 250318 193248
rect 259730 193196 259736 193248
rect 259788 193236 259794 193248
rect 259914 193236 259920 193248
rect 259788 193208 259920 193236
rect 259788 193196 259794 193208
rect 259914 193196 259920 193208
rect 259972 193196 259978 193248
rect 299474 193196 299480 193248
rect 299532 193236 299538 193248
rect 299532 193208 299577 193236
rect 299532 193196 299538 193208
rect 302528 193180 302556 193276
rect 302694 193264 302700 193276
rect 302752 193264 302758 193316
rect 366818 193264 366824 193316
rect 366876 193304 366882 193316
rect 367002 193304 367008 193316
rect 366876 193276 367008 193304
rect 366876 193264 366882 193276
rect 367002 193264 367008 193276
rect 367060 193264 367066 193316
rect 323302 193196 323308 193248
rect 323360 193236 323366 193248
rect 323486 193236 323492 193248
rect 323360 193208 323492 193236
rect 323360 193196 323366 193208
rect 323486 193196 323492 193208
rect 323544 193196 323550 193248
rect 324590 193196 324596 193248
rect 324648 193236 324654 193248
rect 324682 193236 324688 193248
rect 324648 193208 324688 193236
rect 324648 193196 324654 193208
rect 324682 193196 324688 193208
rect 324740 193196 324746 193248
rect 336918 193236 336924 193248
rect 336879 193208 336924 193236
rect 336918 193196 336924 193208
rect 336976 193196 336982 193248
rect 337194 193196 337200 193248
rect 337252 193236 337258 193248
rect 337378 193236 337384 193248
rect 337252 193208 337384 193236
rect 337252 193196 337258 193208
rect 337378 193196 337384 193208
rect 337436 193196 337442 193248
rect 341242 193196 341248 193248
rect 341300 193236 341306 193248
rect 341426 193236 341432 193248
rect 341300 193208 341432 193236
rect 341300 193196 341306 193208
rect 341426 193196 341432 193208
rect 341484 193196 341490 193248
rect 357618 193196 357624 193248
rect 357676 193236 357682 193248
rect 357710 193236 357716 193248
rect 357676 193208 357716 193236
rect 357676 193196 357682 193208
rect 357710 193196 357716 193208
rect 357768 193196 357774 193248
rect 359090 193196 359096 193248
rect 359148 193236 359154 193248
rect 359182 193236 359188 193248
rect 359148 193208 359188 193236
rect 359148 193196 359154 193208
rect 359182 193196 359188 193208
rect 359240 193196 359246 193248
rect 362221 193239 362279 193245
rect 362221 193205 362233 193239
rect 362267 193236 362279 193239
rect 362310 193236 362316 193248
rect 362267 193208 362316 193236
rect 362267 193205 362279 193208
rect 362221 193199 362279 193205
rect 362310 193196 362316 193208
rect 362368 193196 362374 193248
rect 372522 193196 372528 193248
rect 372580 193236 372586 193248
rect 372706 193236 372712 193248
rect 372580 193208 372712 193236
rect 372580 193196 372586 193208
rect 372706 193196 372712 193208
rect 372764 193196 372770 193248
rect 375834 193236 375840 193248
rect 375795 193208 375840 193236
rect 375834 193196 375840 193208
rect 375892 193196 375898 193248
rect 376938 193196 376944 193248
rect 376996 193236 377002 193248
rect 377122 193236 377128 193248
rect 376996 193208 377128 193236
rect 376996 193196 377002 193208
rect 377122 193196 377128 193208
rect 377180 193196 377186 193248
rect 245838 193128 245844 193180
rect 245896 193128 245902 193180
rect 302510 193128 302516 193180
rect 302568 193128 302574 193180
rect 367002 193168 367008 193180
rect 366963 193140 367008 193168
rect 367002 193128 367008 193140
rect 367060 193128 367066 193180
rect 358630 191876 358636 191888
rect 358591 191848 358636 191876
rect 358630 191836 358636 191848
rect 358688 191836 358694 191888
rect 239122 191768 239128 191820
rect 239180 191808 239186 191820
rect 239398 191808 239404 191820
rect 239180 191780 239404 191808
rect 239180 191768 239186 191780
rect 239398 191768 239404 191780
rect 239456 191768 239462 191820
rect 251542 191768 251548 191820
rect 251600 191808 251606 191820
rect 251634 191808 251640 191820
rect 251600 191780 251640 191808
rect 251600 191768 251606 191780
rect 251634 191768 251640 191780
rect 251692 191768 251698 191820
rect 324682 191768 324688 191820
rect 324740 191808 324746 191820
rect 324866 191808 324872 191820
rect 324740 191780 324872 191808
rect 324740 191768 324746 191780
rect 324866 191768 324872 191780
rect 324924 191768 324930 191820
rect 288802 190476 288808 190528
rect 288860 190516 288866 190528
rect 288894 190516 288900 190528
rect 288860 190488 288900 190516
rect 288860 190476 288866 190488
rect 288894 190476 288900 190488
rect 288952 190476 288958 190528
rect 291470 190516 291476 190528
rect 291431 190488 291476 190516
rect 291470 190476 291476 190488
rect 291528 190476 291534 190528
rect 317506 190476 317512 190528
rect 317564 190516 317570 190528
rect 317690 190516 317696 190528
rect 317564 190488 317696 190516
rect 317564 190476 317570 190488
rect 317690 190476 317696 190488
rect 317748 190476 317754 190528
rect 288802 190340 288808 190392
rect 288860 190380 288866 190392
rect 288986 190380 288992 190392
rect 288860 190352 288992 190380
rect 288860 190340 288866 190352
rect 288986 190340 288992 190352
rect 289044 190340 289050 190392
rect 264974 189932 264980 189984
rect 265032 189972 265038 189984
rect 265158 189972 265164 189984
rect 265032 189944 265164 189972
rect 265032 189932 265038 189944
rect 265158 189932 265164 189944
rect 265216 189932 265222 189984
rect 299842 188476 299848 188488
rect 299803 188448 299848 188476
rect 299842 188436 299848 188448
rect 299900 188436 299906 188488
rect 306834 188476 306840 188488
rect 306795 188448 306840 188476
rect 306834 188436 306840 188448
rect 306892 188436 306898 188488
rect 244369 186983 244427 186989
rect 244369 186949 244381 186983
rect 244415 186980 244427 186983
rect 244458 186980 244464 186992
rect 244415 186952 244464 186980
rect 244415 186949 244427 186952
rect 244369 186943 244427 186949
rect 244458 186940 244464 186952
rect 244516 186940 244522 186992
rect 295610 186436 295616 186448
rect 295536 186408 295616 186436
rect 267734 186368 267740 186380
rect 267695 186340 267740 186368
rect 267734 186328 267740 186340
rect 267792 186328 267798 186380
rect 270678 186368 270684 186380
rect 270639 186340 270684 186368
rect 270678 186328 270684 186340
rect 270736 186328 270742 186380
rect 295536 186312 295564 186408
rect 295610 186396 295616 186408
rect 295668 186396 295674 186448
rect 296898 186436 296904 186448
rect 296824 186408 296904 186436
rect 296824 186312 296852 186408
rect 296898 186396 296904 186408
rect 296956 186396 296962 186448
rect 325970 186436 325976 186448
rect 325896 186408 325976 186436
rect 325896 186312 325924 186408
rect 325970 186396 325976 186408
rect 326028 186396 326034 186448
rect 330110 186328 330116 186380
rect 330168 186328 330174 186380
rect 295518 186260 295524 186312
rect 295576 186260 295582 186312
rect 296806 186260 296812 186312
rect 296864 186260 296870 186312
rect 325878 186260 325884 186312
rect 325936 186260 325942 186312
rect 330128 186244 330156 186328
rect 330110 186192 330116 186244
rect 330168 186192 330174 186244
rect 285950 183676 285956 183728
rect 286008 183676 286014 183728
rect 285968 183592 285996 183676
rect 302510 183608 302516 183660
rect 302568 183648 302574 183660
rect 302568 183620 302648 183648
rect 302568 183608 302574 183620
rect 302620 183592 302648 183620
rect 267734 183580 267740 183592
rect 267695 183552 267740 183580
rect 267734 183540 267740 183552
rect 267792 183540 267798 183592
rect 270678 183580 270684 183592
rect 270639 183552 270684 183580
rect 270678 183540 270684 183552
rect 270736 183540 270742 183592
rect 272150 183540 272156 183592
rect 272208 183580 272214 183592
rect 272208 183552 272288 183580
rect 272208 183540 272214 183552
rect 272260 183524 272288 183552
rect 285950 183540 285956 183592
rect 286008 183540 286014 183592
rect 294230 183540 294236 183592
rect 294288 183580 294294 183592
rect 294414 183580 294420 183592
rect 294288 183552 294420 183580
rect 294288 183540 294294 183552
rect 294414 183540 294420 183552
rect 294472 183540 294478 183592
rect 299842 183580 299848 183592
rect 299803 183552 299848 183580
rect 299842 183540 299848 183552
rect 299900 183540 299906 183592
rect 301038 183540 301044 183592
rect 301096 183580 301102 183592
rect 301222 183580 301228 183592
rect 301096 183552 301228 183580
rect 301096 183540 301102 183552
rect 301222 183540 301228 183552
rect 301280 183540 301286 183592
rect 302602 183540 302608 183592
rect 302660 183540 302666 183592
rect 306834 183580 306840 183592
rect 306795 183552 306840 183580
rect 306834 183540 306840 183552
rect 306892 183540 306898 183592
rect 310882 183540 310888 183592
rect 310940 183580 310946 183592
rect 311066 183580 311072 183592
rect 310940 183552 311072 183580
rect 310940 183540 310946 183552
rect 311066 183540 311072 183552
rect 311124 183540 311130 183592
rect 358630 183540 358636 183592
rect 358688 183580 358694 183592
rect 358722 183580 358728 183592
rect 358688 183552 358728 183580
rect 358688 183540 358694 183552
rect 358722 183540 358728 183552
rect 358780 183540 358786 183592
rect 367002 183580 367008 183592
rect 366963 183552 367008 183580
rect 367002 183540 367008 183552
rect 367060 183540 367066 183592
rect 389266 183540 389272 183592
rect 389324 183580 389330 183592
rect 389542 183580 389548 183592
rect 389324 183552 389548 183580
rect 389324 183540 389330 183552
rect 389542 183540 389548 183552
rect 389600 183540 389606 183592
rect 424042 183540 424048 183592
rect 424100 183580 424106 183592
rect 424686 183580 424692 183592
rect 424100 183552 424692 183580
rect 424100 183540 424106 183552
rect 424686 183540 424692 183552
rect 424744 183540 424750 183592
rect 463786 183540 463792 183592
rect 463844 183580 463850 183592
rect 464062 183580 464068 183592
rect 463844 183552 464068 183580
rect 463844 183540 463850 183552
rect 464062 183540 464068 183552
rect 464120 183540 464126 183592
rect 470410 183540 470416 183592
rect 470468 183580 470474 183592
rect 470594 183580 470600 183592
rect 470468 183552 470600 183580
rect 470468 183540 470474 183552
rect 470594 183540 470600 183552
rect 470652 183540 470658 183592
rect 272242 183472 272248 183524
rect 272300 183472 272306 183524
rect 284662 183512 284668 183524
rect 284623 183484 284668 183512
rect 284662 183472 284668 183484
rect 284720 183472 284726 183524
rect 337102 183512 337108 183524
rect 337063 183484 337108 183512
rect 337102 183472 337108 183484
rect 337160 183472 337166 183524
rect 375834 183512 375840 183524
rect 375795 183484 375840 183512
rect 375834 183472 375840 183484
rect 375892 183472 375898 183524
rect 424042 183444 424048 183456
rect 424003 183416 424048 183444
rect 424042 183404 424048 183416
rect 424100 183404 424106 183456
rect 339678 182996 339684 183048
rect 339736 183036 339742 183048
rect 339862 183036 339868 183048
rect 339736 183008 339868 183036
rect 339736 182996 339742 183008
rect 339862 182996 339868 183008
rect 339920 182996 339926 183048
rect 362218 182180 362224 182232
rect 362276 182220 362282 182232
rect 362310 182220 362316 182232
rect 362276 182192 362316 182220
rect 362276 182180 362282 182192
rect 362310 182180 362316 182192
rect 362368 182180 362374 182232
rect 251450 182112 251456 182164
rect 251508 182152 251514 182164
rect 251726 182152 251732 182164
rect 251508 182124 251732 182152
rect 251508 182112 251514 182124
rect 251726 182112 251732 182124
rect 251784 182112 251790 182164
rect 299842 182112 299848 182164
rect 299900 182152 299906 182164
rect 299934 182152 299940 182164
rect 299900 182124 299940 182152
rect 299900 182112 299906 182124
rect 299934 182112 299940 182124
rect 299992 182112 299998 182164
rect 327350 182112 327356 182164
rect 327408 182152 327414 182164
rect 327534 182152 327540 182164
rect 327408 182124 327540 182152
rect 327408 182112 327414 182124
rect 327534 182112 327540 182124
rect 327592 182112 327598 182164
rect 329926 182112 329932 182164
rect 329984 182152 329990 182164
rect 330110 182152 330116 182164
rect 329984 182124 330116 182152
rect 329984 182112 329990 182124
rect 330110 182112 330116 182124
rect 330168 182112 330174 182164
rect 339494 182112 339500 182164
rect 339552 182152 339558 182164
rect 339678 182152 339684 182164
rect 339552 182124 339684 182152
rect 339552 182112 339558 182124
rect 339678 182112 339684 182124
rect 339736 182112 339742 182164
rect 341150 182112 341156 182164
rect 341208 182152 341214 182164
rect 341426 182152 341432 182164
rect 341208 182124 341432 182152
rect 341208 182112 341214 182124
rect 341426 182112 341432 182124
rect 341484 182112 341490 182164
rect 358538 182112 358544 182164
rect 358596 182152 358602 182164
rect 358722 182152 358728 182164
rect 358596 182124 358728 182152
rect 358596 182112 358602 182124
rect 358722 182112 358728 182124
rect 358780 182112 358786 182164
rect 421190 182112 421196 182164
rect 421248 182152 421254 182164
rect 421374 182152 421380 182164
rect 421248 182124 421380 182152
rect 421248 182112 421254 182124
rect 421374 182112 421380 182124
rect 421432 182112 421438 182164
rect 244366 180860 244372 180872
rect 244327 180832 244372 180860
rect 244366 180820 244372 180832
rect 244424 180820 244430 180872
rect 251174 180752 251180 180804
rect 251232 180792 251238 180804
rect 251450 180792 251456 180804
rect 251232 180764 251456 180792
rect 251232 180752 251238 180764
rect 251450 180752 251456 180764
rect 251508 180752 251514 180804
rect 265158 180752 265164 180804
rect 265216 180792 265222 180804
rect 265250 180792 265256 180804
rect 265216 180764 265256 180792
rect 265216 180752 265222 180764
rect 265250 180752 265256 180764
rect 265308 180752 265314 180804
rect 284662 180792 284668 180804
rect 284623 180764 284668 180792
rect 284662 180752 284668 180764
rect 284720 180752 284726 180804
rect 285950 180792 285956 180804
rect 285911 180764 285956 180792
rect 285950 180752 285956 180764
rect 286008 180752 286014 180804
rect 288710 180792 288716 180804
rect 288671 180764 288716 180792
rect 288710 180752 288716 180764
rect 288768 180752 288774 180804
rect 317506 180752 317512 180804
rect 317564 180792 317570 180804
rect 317690 180792 317696 180804
rect 317564 180764 317696 180792
rect 317564 180752 317570 180764
rect 317690 180752 317696 180764
rect 317748 180752 317754 180804
rect 265161 179367 265219 179373
rect 265161 179333 265173 179367
rect 265207 179364 265219 179367
rect 265250 179364 265256 179376
rect 265207 179336 265256 179364
rect 265207 179333 265219 179336
rect 265161 179327 265219 179333
rect 265250 179324 265256 179336
rect 265308 179324 265314 179376
rect 358998 179364 359004 179376
rect 358959 179336 359004 179364
rect 358998 179324 359004 179336
rect 359056 179324 359062 179376
rect 294230 178712 294236 178764
rect 294288 178752 294294 178764
rect 294414 178752 294420 178764
rect 294288 178724 294420 178752
rect 294288 178712 294294 178724
rect 294414 178712 294420 178724
rect 294472 178712 294478 178764
rect 295518 178712 295524 178764
rect 295576 178752 295582 178764
rect 295702 178752 295708 178764
rect 295576 178724 295708 178752
rect 295576 178712 295582 178724
rect 295702 178712 295708 178724
rect 295760 178712 295766 178764
rect 337105 178755 337163 178761
rect 337105 178721 337117 178755
rect 337151 178752 337163 178755
rect 337194 178752 337200 178764
rect 337151 178724 337200 178752
rect 337151 178721 337163 178724
rect 337105 178715 337163 178721
rect 337194 178712 337200 178724
rect 337252 178712 337258 178764
rect 288713 177871 288771 177877
rect 288713 177837 288725 177871
rect 288759 177868 288771 177871
rect 289078 177868 289084 177880
rect 288759 177840 289084 177868
rect 288759 177837 288771 177840
rect 288713 177831 288771 177837
rect 289078 177828 289084 177840
rect 289136 177828 289142 177880
rect 302602 176780 302608 176792
rect 302528 176752 302608 176780
rect 232222 176672 232228 176724
rect 232280 176672 232286 176724
rect 301038 176672 301044 176724
rect 301096 176672 301102 176724
rect 232240 176644 232268 176672
rect 232314 176644 232320 176656
rect 232240 176616 232320 176644
rect 232314 176604 232320 176616
rect 232372 176604 232378 176656
rect 301056 176576 301084 176672
rect 302528 176656 302556 176752
rect 302602 176740 302608 176752
rect 302660 176740 302666 176792
rect 306834 176780 306840 176792
rect 306760 176752 306840 176780
rect 306760 176656 306788 176752
rect 306834 176740 306840 176752
rect 306892 176740 306898 176792
rect 310882 176780 310888 176792
rect 310808 176752 310888 176780
rect 310808 176656 310836 176752
rect 310882 176740 310888 176752
rect 310940 176740 310946 176792
rect 389542 176780 389548 176792
rect 389468 176752 389548 176780
rect 389468 176656 389496 176752
rect 389542 176740 389548 176752
rect 389600 176740 389606 176792
rect 463878 176672 463884 176724
rect 463936 176712 463942 176724
rect 464062 176712 464068 176724
rect 463936 176684 464068 176712
rect 463936 176672 463942 176684
rect 464062 176672 464068 176684
rect 464120 176672 464126 176724
rect 302510 176604 302516 176656
rect 302568 176604 302574 176656
rect 306742 176604 306748 176656
rect 306800 176604 306806 176656
rect 310790 176604 310796 176656
rect 310848 176604 310854 176656
rect 389450 176604 389456 176656
rect 389508 176604 389514 176656
rect 301130 176576 301136 176588
rect 301056 176548 301136 176576
rect 301130 176536 301136 176548
rect 301188 176536 301194 176588
rect 424045 176579 424103 176585
rect 424045 176545 424057 176579
rect 424091 176576 424103 176579
rect 424226 176576 424232 176588
rect 424091 176548 424232 176576
rect 424091 176545 424103 176548
rect 424045 176539 424103 176545
rect 424226 176536 424232 176548
rect 424284 176536 424290 176588
rect 285950 175964 285956 175976
rect 285911 175936 285956 175964
rect 285950 175924 285956 175936
rect 286008 175924 286014 175976
rect 266722 174060 266728 174072
rect 266648 174032 266728 174060
rect 236270 173952 236276 174004
rect 236328 173952 236334 174004
rect 236288 173868 236316 173952
rect 266648 173936 266676 174032
rect 266722 174020 266728 174032
rect 266780 174020 266786 174072
rect 270494 173952 270500 174004
rect 270552 173992 270558 174004
rect 270678 173992 270684 174004
rect 270552 173964 270684 173992
rect 270552 173952 270558 173964
rect 270678 173952 270684 173964
rect 270736 173952 270742 174004
rect 372614 173952 372620 174004
rect 372672 173992 372678 174004
rect 372798 173992 372804 174004
rect 372672 173964 372804 173992
rect 372672 173952 372678 173964
rect 372798 173952 372804 173964
rect 372856 173952 372862 174004
rect 244366 173884 244372 173936
rect 244424 173924 244430 173936
rect 244458 173924 244464 173936
rect 244424 173896 244464 173924
rect 244424 173884 244430 173896
rect 244458 173884 244464 173896
rect 244516 173884 244522 173936
rect 245838 173884 245844 173936
rect 245896 173924 245902 173936
rect 245930 173924 245936 173936
rect 245896 173896 245936 173924
rect 245896 173884 245902 173896
rect 245930 173884 245936 173896
rect 245988 173884 245994 173936
rect 250070 173884 250076 173936
rect 250128 173924 250134 173936
rect 250254 173924 250260 173936
rect 250128 173896 250260 173924
rect 250128 173884 250134 173896
rect 250254 173884 250260 173896
rect 250312 173884 250318 173936
rect 259638 173924 259644 173936
rect 259599 173896 259644 173924
rect 259638 173884 259644 173896
rect 259696 173884 259702 173936
rect 262582 173884 262588 173936
rect 262640 173924 262646 173936
rect 262674 173924 262680 173936
rect 262640 173896 262680 173924
rect 262640 173884 262646 173896
rect 262674 173884 262680 173896
rect 262732 173884 262738 173936
rect 266630 173884 266636 173936
rect 266688 173884 266694 173936
rect 267826 173884 267832 173936
rect 267884 173924 267890 173936
rect 267918 173924 267924 173936
rect 267884 173896 267924 173924
rect 267884 173884 267890 173896
rect 267918 173884 267924 173896
rect 267976 173884 267982 173936
rect 323302 173884 323308 173936
rect 323360 173924 323366 173936
rect 323486 173924 323492 173936
rect 323360 173896 323492 173924
rect 323360 173884 323366 173896
rect 323486 173884 323492 173896
rect 323544 173884 323550 173936
rect 325878 173884 325884 173936
rect 325936 173924 325942 173936
rect 325970 173924 325976 173936
rect 325936 173896 325976 173924
rect 325936 173884 325942 173896
rect 325970 173884 325976 173896
rect 326028 173884 326034 173936
rect 336734 173884 336740 173936
rect 336792 173924 336798 173936
rect 336918 173924 336924 173936
rect 336792 173896 336924 173924
rect 336792 173884 336798 173896
rect 336918 173884 336924 173896
rect 336976 173884 336982 173936
rect 375834 173924 375840 173936
rect 375795 173896 375840 173924
rect 375834 173884 375840 173896
rect 375892 173884 375898 173936
rect 376938 173884 376944 173936
rect 376996 173924 377002 173936
rect 377122 173924 377128 173936
rect 376996 173896 377128 173924
rect 376996 173884 377002 173896
rect 377122 173884 377128 173896
rect 377180 173884 377186 173936
rect 236270 173816 236276 173868
rect 236328 173816 236334 173868
rect 239122 172592 239128 172644
rect 239180 172632 239186 172644
rect 239398 172632 239404 172644
rect 239180 172604 239404 172632
rect 239180 172592 239186 172604
rect 239398 172592 239404 172604
rect 239456 172592 239462 172644
rect 259638 172564 259644 172576
rect 259599 172536 259644 172564
rect 259638 172524 259644 172536
rect 259696 172524 259702 172576
rect 296898 172456 296904 172508
rect 296956 172496 296962 172508
rect 296990 172496 296996 172508
rect 296956 172468 296996 172496
rect 296956 172456 296962 172468
rect 296990 172456 296996 172468
rect 297048 172456 297054 172508
rect 324593 172499 324651 172505
rect 324593 172465 324605 172499
rect 324639 172496 324651 172499
rect 324682 172496 324688 172508
rect 324639 172468 324688 172496
rect 324639 172465 324651 172468
rect 324593 172459 324651 172465
rect 324682 172456 324688 172468
rect 324740 172456 324746 172508
rect 360286 171068 360292 171080
rect 360247 171040 360292 171068
rect 360286 171028 360292 171040
rect 360344 171028 360350 171080
rect 362221 171071 362279 171077
rect 362221 171037 362233 171071
rect 362267 171068 362279 171071
rect 362310 171068 362316 171080
rect 362267 171040 362316 171068
rect 362267 171037 362279 171040
rect 362221 171031 362279 171037
rect 362310 171028 362316 171040
rect 362368 171028 362374 171080
rect 359001 169779 359059 169785
rect 359001 169745 359013 169779
rect 359047 169776 359059 169779
rect 359090 169776 359096 169788
rect 359047 169748 359096 169776
rect 359047 169745 359059 169748
rect 359001 169739 359059 169745
rect 359090 169736 359096 169748
rect 359148 169736 359154 169788
rect 289078 169708 289084 169720
rect 289039 169680 289084 169708
rect 289078 169668 289084 169680
rect 289136 169668 289142 169720
rect 302510 169532 302516 169584
rect 302568 169572 302574 169584
rect 302786 169572 302792 169584
rect 302568 169544 302792 169572
rect 302568 169532 302574 169544
rect 302786 169532 302792 169544
rect 302844 169532 302850 169584
rect 306742 169532 306748 169584
rect 306800 169572 306806 169584
rect 307018 169572 307024 169584
rect 306800 169544 307024 169572
rect 306800 169532 306806 169544
rect 307018 169532 307024 169544
rect 307076 169532 307082 169584
rect 270494 169056 270500 169108
rect 270552 169096 270558 169108
rect 270678 169096 270684 169108
rect 270552 169068 270684 169096
rect 270552 169056 270558 169068
rect 270678 169056 270684 169068
rect 270736 169056 270742 169108
rect 272150 167016 272156 167068
rect 272208 167056 272214 167068
rect 272208 167028 272288 167056
rect 272208 167016 272214 167028
rect 272260 167000 272288 167028
rect 310790 167016 310796 167068
rect 310848 167016 310854 167068
rect 272242 166948 272248 167000
rect 272300 166948 272306 167000
rect 310808 166920 310836 167016
rect 424226 166948 424232 167000
rect 424284 166948 424290 167000
rect 310882 166920 310888 166932
rect 310808 166892 310888 166920
rect 310882 166880 310888 166892
rect 310940 166880 310946 166932
rect 424244 166920 424272 166948
rect 424410 166920 424416 166932
rect 424244 166892 424416 166920
rect 424410 166880 424416 166892
rect 424468 166880 424474 166932
rect 2774 165452 2780 165504
rect 2832 165492 2838 165504
rect 5166 165492 5172 165504
rect 2832 165464 5172 165492
rect 2832 165452 2838 165464
rect 5166 165452 5172 165464
rect 5224 165452 5230 165504
rect 330110 164296 330116 164348
rect 330168 164336 330174 164348
rect 330202 164336 330208 164348
rect 330168 164308 330208 164336
rect 330168 164296 330174 164308
rect 330202 164296 330208 164308
rect 330260 164296 330266 164348
rect 239122 164228 239128 164280
rect 239180 164228 239186 164280
rect 239140 164132 239168 164228
rect 244366 164160 244372 164212
rect 244424 164200 244430 164212
rect 244550 164200 244556 164212
rect 244424 164172 244556 164200
rect 244424 164160 244430 164172
rect 244550 164160 244556 164172
rect 244608 164160 244614 164212
rect 372798 164200 372804 164212
rect 372759 164172 372804 164200
rect 372798 164160 372804 164172
rect 372856 164160 372862 164212
rect 375834 164200 375840 164212
rect 375795 164172 375840 164200
rect 375834 164160 375840 164172
rect 375892 164160 375898 164212
rect 376938 164160 376944 164212
rect 376996 164200 377002 164212
rect 377122 164200 377128 164212
rect 376996 164172 377128 164200
rect 376996 164160 377002 164172
rect 377122 164160 377128 164172
rect 377180 164160 377186 164212
rect 424410 164160 424416 164212
rect 424468 164200 424474 164212
rect 424502 164200 424508 164212
rect 424468 164172 424508 164200
rect 424468 164160 424474 164172
rect 424502 164160 424508 164172
rect 424560 164160 424566 164212
rect 463786 164160 463792 164212
rect 463844 164200 463850 164212
rect 464062 164200 464068 164212
rect 463844 164172 464068 164200
rect 463844 164160 463850 164172
rect 464062 164160 464068 164172
rect 464120 164160 464126 164212
rect 239306 164132 239312 164144
rect 239140 164104 239312 164132
rect 239306 164092 239312 164104
rect 239364 164092 239370 164144
rect 284662 162908 284668 162920
rect 284623 162880 284668 162908
rect 284662 162868 284668 162880
rect 284720 162868 284726 162920
rect 294322 162868 294328 162920
rect 294380 162908 294386 162920
rect 294414 162908 294420 162920
rect 294380 162880 294420 162908
rect 294380 162868 294386 162880
rect 294414 162868 294420 162880
rect 294472 162868 294478 162920
rect 324590 162908 324596 162920
rect 324551 162880 324596 162908
rect 324590 162868 324596 162880
rect 324648 162868 324654 162920
rect 236270 162800 236276 162852
rect 236328 162840 236334 162852
rect 236454 162840 236460 162852
rect 236328 162812 236460 162840
rect 236328 162800 236334 162812
rect 236454 162800 236460 162812
rect 236512 162800 236518 162852
rect 245838 162840 245844 162852
rect 245799 162812 245844 162840
rect 245838 162800 245844 162812
rect 245896 162800 245902 162852
rect 250070 162800 250076 162852
rect 250128 162800 250134 162852
rect 272058 162840 272064 162852
rect 272019 162812 272064 162840
rect 272058 162800 272064 162812
rect 272116 162800 272122 162852
rect 302513 162843 302571 162849
rect 302513 162809 302525 162843
rect 302559 162840 302571 162843
rect 302602 162840 302608 162852
rect 302559 162812 302608 162840
rect 302559 162809 302571 162812
rect 302513 162803 302571 162809
rect 302602 162800 302608 162812
rect 302660 162800 302666 162852
rect 306742 162800 306748 162852
rect 306800 162840 306806 162852
rect 306834 162840 306840 162852
rect 306800 162812 306840 162840
rect 306800 162800 306806 162812
rect 306834 162800 306840 162812
rect 306892 162800 306898 162852
rect 327166 162800 327172 162852
rect 327224 162840 327230 162852
rect 327442 162840 327448 162852
rect 327224 162812 327448 162840
rect 327224 162800 327230 162812
rect 327442 162800 327448 162812
rect 327500 162800 327506 162852
rect 358630 162800 358636 162852
rect 358688 162840 358694 162852
rect 358722 162840 358728 162852
rect 358688 162812 358728 162840
rect 358688 162800 358694 162812
rect 358722 162800 358728 162812
rect 358780 162800 358786 162852
rect 358998 162800 359004 162852
rect 359056 162840 359062 162852
rect 359090 162840 359096 162852
rect 359056 162812 359096 162840
rect 359056 162800 359062 162812
rect 359090 162800 359096 162812
rect 359148 162800 359154 162852
rect 421190 162840 421196 162852
rect 421151 162812 421196 162840
rect 421190 162800 421196 162812
rect 421248 162800 421254 162852
rect 239030 162732 239036 162784
rect 239088 162772 239094 162784
rect 239306 162772 239312 162784
rect 239088 162744 239312 162772
rect 239088 162732 239094 162744
rect 239306 162732 239312 162744
rect 239364 162732 239370 162784
rect 250088 162772 250116 162800
rect 250346 162772 250352 162784
rect 250088 162744 250352 162772
rect 250346 162732 250352 162744
rect 250404 162732 250410 162784
rect 259546 161440 259552 161492
rect 259604 161480 259610 161492
rect 259638 161480 259644 161492
rect 259604 161452 259644 161480
rect 259604 161440 259610 161452
rect 259638 161440 259644 161452
rect 259696 161440 259702 161492
rect 265158 161480 265164 161492
rect 265119 161452 265164 161480
rect 265158 161440 265164 161452
rect 265216 161440 265222 161492
rect 360289 161483 360347 161489
rect 360289 161449 360301 161483
rect 360335 161480 360347 161483
rect 360470 161480 360476 161492
rect 360335 161452 360476 161480
rect 360335 161449 360347 161452
rect 360289 161443 360347 161449
rect 360470 161440 360476 161452
rect 360528 161440 360534 161492
rect 362218 161480 362224 161492
rect 362179 161452 362224 161480
rect 362218 161440 362224 161452
rect 362276 161440 362282 161492
rect 250346 161412 250352 161424
rect 250307 161384 250352 161412
rect 250346 161372 250352 161384
rect 250404 161372 250410 161424
rect 359090 161412 359096 161424
rect 359051 161384 359096 161412
rect 359090 161372 359096 161384
rect 359148 161372 359154 161424
rect 289078 160120 289084 160132
rect 289039 160092 289084 160120
rect 289078 160080 289084 160092
rect 289136 160080 289142 160132
rect 299750 159332 299756 159384
rect 299808 159372 299814 159384
rect 299934 159372 299940 159384
rect 299808 159344 299940 159372
rect 299808 159332 299814 159344
rect 299934 159332 299940 159344
rect 299992 159332 299998 159384
rect 341058 159332 341064 159384
rect 341116 159372 341122 159384
rect 341242 159372 341248 159384
rect 341116 159344 341248 159372
rect 341116 159332 341122 159344
rect 341242 159332 341248 159344
rect 341300 159332 341306 159384
rect 417878 157564 417884 157616
rect 417936 157604 417942 157616
rect 418246 157604 418252 157616
rect 417936 157576 418252 157604
rect 417936 157564 417942 157576
rect 418246 157564 418252 157576
rect 418304 157564 418310 157616
rect 298002 157496 298008 157548
rect 298060 157536 298066 157548
rect 306282 157536 306288 157548
rect 298060 157508 306288 157536
rect 298060 157496 298066 157508
rect 306282 157496 306288 157508
rect 306340 157496 306346 157548
rect 437198 157496 437204 157548
rect 437256 157536 437262 157548
rect 437474 157536 437480 157548
rect 437256 157508 437480 157536
rect 437256 157496 437262 157508
rect 437474 157496 437480 157508
rect 437532 157496 437538 157548
rect 456518 157496 456524 157548
rect 456576 157536 456582 157548
rect 456886 157536 456892 157548
rect 456576 157508 456892 157536
rect 456576 157496 456582 157508
rect 456886 157496 456892 157508
rect 456944 157496 456950 157548
rect 273530 157428 273536 157480
rect 273588 157428 273594 157480
rect 307570 157428 307576 157480
rect 307628 157468 307634 157480
rect 315942 157468 315948 157480
rect 307628 157440 315948 157468
rect 307628 157428 307634 157440
rect 315942 157428 315948 157440
rect 316000 157428 316006 157480
rect 267734 157360 267740 157412
rect 267792 157360 267798 157412
rect 267752 157276 267780 157360
rect 273548 157344 273576 157428
rect 295518 157360 295524 157412
rect 295576 157400 295582 157412
rect 295702 157400 295708 157412
rect 295576 157372 295708 157400
rect 295576 157360 295582 157372
rect 295702 157360 295708 157372
rect 295760 157360 295766 157412
rect 296806 157360 296812 157412
rect 296864 157400 296870 157412
rect 296990 157400 296996 157412
rect 296864 157372 296996 157400
rect 296864 157360 296870 157372
rect 296990 157360 296996 157372
rect 297048 157360 297054 157412
rect 337102 157360 337108 157412
rect 337160 157360 337166 157412
rect 273530 157292 273536 157344
rect 273588 157292 273594 157344
rect 267734 157224 267740 157276
rect 267792 157224 267798 157276
rect 325970 157224 325976 157276
rect 326028 157224 326034 157276
rect 337120 157264 337148 157360
rect 372798 157332 372804 157344
rect 372759 157304 372804 157332
rect 372798 157292 372804 157304
rect 372856 157292 372862 157344
rect 337194 157264 337200 157276
rect 337120 157236 337200 157264
rect 337194 157224 337200 157236
rect 337252 157224 337258 157276
rect 270678 157156 270684 157208
rect 270736 157156 270742 157208
rect 270696 157128 270724 157156
rect 325988 157140 326016 157224
rect 270770 157128 270776 157140
rect 270696 157100 270776 157128
rect 270770 157088 270776 157100
rect 270828 157088 270834 157140
rect 325970 157088 325976 157140
rect 326028 157088 326034 157140
rect 375834 154612 375840 154624
rect 375795 154584 375840 154612
rect 375834 154572 375840 154584
rect 375892 154572 375898 154624
rect 232314 154544 232320 154556
rect 232275 154516 232320 154544
rect 232314 154504 232320 154516
rect 232372 154504 232378 154556
rect 272061 154547 272119 154553
rect 272061 154513 272073 154547
rect 272107 154544 272119 154547
rect 272242 154544 272248 154556
rect 272107 154516 272248 154544
rect 272107 154513 272119 154516
rect 272061 154507 272119 154513
rect 272242 154504 272248 154516
rect 272300 154504 272306 154556
rect 341058 154504 341064 154556
rect 341116 154544 341122 154556
rect 341242 154544 341248 154556
rect 341116 154516 341248 154544
rect 341116 154504 341122 154516
rect 341242 154504 341248 154516
rect 341300 154504 341306 154556
rect 389450 154504 389456 154556
rect 389508 154544 389514 154556
rect 389634 154544 389640 154556
rect 389508 154516 389640 154544
rect 389508 154504 389514 154516
rect 389634 154504 389640 154516
rect 389692 154504 389698 154556
rect 470410 154504 470416 154556
rect 470468 154544 470474 154556
rect 470594 154544 470600 154556
rect 470468 154516 470600 154544
rect 470468 154504 470474 154516
rect 470594 154504 470600 154516
rect 470652 154504 470658 154556
rect 245841 154479 245899 154485
rect 245841 154445 245853 154479
rect 245887 154476 245899 154479
rect 245930 154476 245936 154488
rect 245887 154448 245936 154476
rect 245887 154445 245899 154448
rect 245841 154439 245899 154445
rect 245930 154436 245936 154448
rect 245988 154436 245994 154488
rect 301038 154436 301044 154488
rect 301096 154476 301102 154488
rect 301222 154476 301228 154488
rect 301096 154448 301228 154476
rect 301096 154436 301102 154448
rect 301222 154436 301228 154448
rect 301280 154436 301286 154488
rect 302510 153252 302516 153264
rect 302471 153224 302516 153252
rect 302510 153212 302516 153224
rect 302568 153212 302574 153264
rect 421190 153252 421196 153264
rect 421151 153224 421196 153252
rect 421190 153212 421196 153224
rect 421248 153212 421254 153264
rect 245930 153184 245936 153196
rect 245891 153156 245936 153184
rect 245930 153144 245936 153156
rect 245988 153144 245994 153196
rect 265158 153144 265164 153196
rect 265216 153184 265222 153196
rect 265342 153184 265348 153196
rect 265216 153156 265348 153184
rect 265216 153144 265222 153156
rect 265342 153144 265348 153156
rect 265400 153144 265406 153196
rect 266630 153184 266636 153196
rect 266591 153156 266636 153184
rect 266630 153144 266636 153156
rect 266688 153144 266694 153196
rect 285950 153144 285956 153196
rect 286008 153184 286014 153196
rect 286042 153184 286048 153196
rect 286008 153156 286048 153184
rect 286008 153144 286014 153156
rect 286042 153144 286048 153156
rect 286100 153144 286106 153196
rect 310790 153184 310796 153196
rect 310751 153156 310796 153184
rect 310790 153144 310796 153156
rect 310848 153144 310854 153196
rect 337105 153187 337163 153193
rect 337105 153153 337117 153187
rect 337151 153184 337163 153187
rect 337194 153184 337200 153196
rect 337151 153156 337200 153184
rect 337151 153153 337163 153156
rect 337105 153147 337163 153153
rect 337194 153144 337200 153156
rect 337252 153144 337258 153196
rect 302510 153076 302516 153128
rect 302568 153116 302574 153128
rect 302786 153116 302792 153128
rect 302568 153088 302792 153116
rect 302568 153076 302574 153088
rect 302786 153076 302792 153088
rect 302844 153076 302850 153128
rect 250346 151824 250352 151836
rect 250307 151796 250352 151824
rect 250346 151784 250352 151796
rect 250404 151784 250410 151836
rect 359093 151827 359151 151833
rect 359093 151793 359105 151827
rect 359139 151824 359151 151827
rect 359182 151824 359188 151836
rect 359139 151796 359188 151824
rect 359139 151793 359151 151796
rect 359093 151787 359151 151793
rect 359182 151784 359188 151796
rect 359240 151784 359246 151836
rect 3326 151716 3332 151768
rect 3384 151756 3390 151768
rect 17218 151756 17224 151768
rect 3384 151728 17224 151756
rect 3384 151716 3390 151728
rect 17218 151716 17224 151728
rect 17276 151716 17282 151768
rect 288805 150399 288863 150405
rect 288805 150365 288817 150399
rect 288851 150396 288863 150399
rect 288986 150396 288992 150408
rect 288851 150368 288992 150396
rect 288851 150365 288863 150368
rect 288805 150359 288863 150365
rect 288986 150356 288992 150368
rect 289044 150356 289050 150408
rect 284662 147704 284668 147756
rect 284720 147704 284726 147756
rect 284680 147620 284708 147704
rect 284662 147568 284668 147620
rect 284720 147568 284726 147620
rect 310790 147608 310796 147620
rect 310751 147580 310796 147608
rect 310790 147568 310796 147580
rect 310848 147568 310854 147620
rect 232314 144956 232320 144968
rect 232275 144928 232320 144956
rect 232314 144916 232320 144928
rect 232372 144916 232378 144968
rect 250346 144956 250352 144968
rect 250180 144928 250352 144956
rect 250180 144900 250208 144928
rect 250346 144916 250352 144928
rect 250404 144916 250410 144968
rect 250162 144848 250168 144900
rect 250220 144848 250226 144900
rect 262582 144848 262588 144900
rect 262640 144888 262646 144900
rect 262766 144888 262772 144900
rect 262640 144860 262772 144888
rect 262640 144848 262646 144860
rect 262766 144848 262772 144860
rect 262824 144848 262830 144900
rect 266630 144888 266636 144900
rect 266591 144860 266636 144888
rect 266630 144848 266636 144860
rect 266688 144848 266694 144900
rect 267734 144848 267740 144900
rect 267792 144888 267798 144900
rect 267918 144888 267924 144900
rect 267792 144860 267924 144888
rect 267792 144848 267798 144860
rect 267918 144848 267924 144860
rect 267976 144848 267982 144900
rect 270678 144848 270684 144900
rect 270736 144888 270742 144900
rect 270954 144888 270960 144900
rect 270736 144860 270960 144888
rect 270736 144848 270742 144860
rect 270954 144848 270960 144860
rect 271012 144848 271018 144900
rect 272150 144848 272156 144900
rect 272208 144888 272214 144900
rect 272426 144888 272432 144900
rect 272208 144860 272432 144888
rect 272208 144848 272214 144860
rect 272426 144848 272432 144860
rect 272484 144848 272490 144900
rect 273530 144888 273536 144900
rect 273491 144860 273536 144888
rect 273530 144848 273536 144860
rect 273588 144848 273594 144900
rect 323302 144848 323308 144900
rect 323360 144888 323366 144900
rect 323394 144888 323400 144900
rect 323360 144860 323400 144888
rect 323360 144848 323366 144860
rect 323394 144848 323400 144860
rect 323452 144848 323458 144900
rect 324590 144848 324596 144900
rect 324648 144888 324654 144900
rect 324774 144888 324780 144900
rect 324648 144860 324780 144888
rect 324648 144848 324654 144860
rect 324774 144848 324780 144860
rect 324832 144848 324838 144900
rect 325878 144848 325884 144900
rect 325936 144888 325942 144900
rect 326062 144888 326068 144900
rect 325936 144860 326068 144888
rect 325936 144848 325942 144860
rect 326062 144848 326068 144860
rect 326120 144848 326126 144900
rect 327166 144848 327172 144900
rect 327224 144888 327230 144900
rect 327258 144888 327264 144900
rect 327224 144860 327264 144888
rect 327224 144848 327230 144860
rect 327258 144848 327264 144860
rect 327316 144848 327322 144900
rect 359182 144848 359188 144900
rect 359240 144888 359246 144900
rect 359274 144888 359280 144900
rect 359240 144860 359280 144888
rect 359240 144848 359246 144860
rect 359274 144848 359280 144860
rect 359332 144848 359338 144900
rect 362126 144848 362132 144900
rect 362184 144888 362190 144900
rect 362310 144888 362316 144900
rect 362184 144860 362316 144888
rect 362184 144848 362190 144860
rect 362310 144848 362316 144860
rect 362368 144848 362374 144900
rect 367002 144888 367008 144900
rect 366963 144860 367008 144888
rect 367002 144848 367008 144860
rect 367060 144848 367066 144900
rect 375834 144888 375840 144900
rect 375795 144860 375840 144888
rect 375834 144848 375840 144860
rect 375892 144848 375898 144900
rect 376938 144848 376944 144900
rect 376996 144888 377002 144900
rect 377122 144888 377128 144900
rect 376996 144860 377128 144888
rect 376996 144848 377002 144860
rect 377122 144848 377128 144860
rect 377180 144848 377186 144900
rect 329926 144304 329932 144356
rect 329984 144344 329990 144356
rect 330386 144344 330392 144356
rect 329984 144316 330392 144344
rect 329984 144304 329990 144316
rect 330386 144304 330392 144316
rect 330444 144304 330450 144356
rect 245930 143596 245936 143608
rect 245891 143568 245936 143596
rect 245930 143556 245936 143568
rect 245988 143556 245994 143608
rect 337102 143596 337108 143608
rect 337063 143568 337108 143596
rect 337102 143556 337108 143568
rect 337160 143556 337166 143608
rect 232314 143528 232320 143540
rect 232275 143500 232320 143528
rect 232314 143488 232320 143500
rect 232372 143488 232378 143540
rect 244458 143528 244464 143540
rect 244419 143500 244464 143528
rect 244458 143488 244464 143500
rect 244516 143488 244522 143540
rect 250162 143488 250168 143540
rect 250220 143528 250226 143540
rect 250254 143528 250260 143540
rect 250220 143500 250260 143528
rect 250220 143488 250226 143500
rect 250254 143488 250260 143500
rect 250312 143488 250318 143540
rect 270954 143528 270960 143540
rect 270915 143500 270960 143528
rect 270954 143488 270960 143500
rect 271012 143488 271018 143540
rect 272334 143488 272340 143540
rect 272392 143528 272398 143540
rect 272426 143528 272432 143540
rect 272392 143500 272432 143528
rect 272392 143488 272398 143500
rect 272426 143488 272432 143500
rect 272484 143488 272490 143540
rect 302418 143488 302424 143540
rect 302476 143528 302482 143540
rect 302602 143528 302608 143540
rect 302476 143500 302608 143528
rect 302476 143488 302482 143500
rect 302602 143488 302608 143500
rect 302660 143488 302666 143540
rect 323302 143488 323308 143540
rect 323360 143528 323366 143540
rect 323486 143528 323492 143540
rect 323360 143500 323492 143528
rect 323360 143488 323366 143500
rect 323486 143488 323492 143500
rect 323544 143488 323550 143540
rect 327258 143528 327264 143540
rect 327219 143500 327264 143528
rect 327258 143488 327264 143500
rect 327316 143488 327322 143540
rect 358722 143528 358728 143540
rect 358683 143500 358728 143528
rect 358722 143488 358728 143500
rect 358780 143488 358786 143540
rect 362310 143488 362316 143540
rect 362368 143528 362374 143540
rect 362494 143528 362500 143540
rect 362368 143500 362500 143528
rect 362368 143488 362374 143500
rect 362494 143488 362500 143500
rect 362552 143488 362558 143540
rect 421190 143528 421196 143540
rect 421151 143500 421196 143528
rect 421190 143488 421196 143500
rect 421248 143488 421254 143540
rect 424134 142808 424140 142860
rect 424192 142848 424198 142860
rect 424594 142848 424600 142860
rect 424192 142820 424600 142848
rect 424192 142808 424198 142820
rect 424594 142808 424600 142820
rect 424652 142808 424658 142860
rect 317506 142128 317512 142180
rect 317564 142168 317570 142180
rect 317690 142168 317696 142180
rect 317564 142140 317696 142168
rect 317564 142128 317570 142140
rect 317690 142128 317696 142140
rect 317748 142128 317754 142180
rect 249981 142103 250039 142109
rect 249981 142069 249993 142103
rect 250027 142100 250039 142103
rect 250254 142100 250260 142112
rect 250027 142072 250260 142100
rect 250027 142069 250039 142072
rect 249981 142063 250039 142069
rect 250254 142060 250260 142072
rect 250312 142060 250318 142112
rect 259638 142100 259644 142112
rect 259599 142072 259644 142100
rect 259638 142060 259644 142072
rect 259696 142060 259702 142112
rect 286045 142103 286103 142109
rect 286045 142069 286057 142103
rect 286091 142100 286103 142103
rect 286134 142100 286140 142112
rect 286091 142072 286140 142100
rect 286091 142069 286103 142072
rect 286045 142063 286103 142069
rect 286134 142060 286140 142072
rect 286192 142060 286198 142112
rect 296901 142103 296959 142109
rect 296901 142069 296913 142103
rect 296947 142100 296959 142103
rect 296990 142100 296996 142112
rect 296947 142072 296996 142100
rect 296947 142069 296959 142072
rect 296901 142063 296959 142069
rect 296990 142060 296996 142072
rect 297048 142060 297054 142112
rect 288802 140808 288808 140820
rect 288763 140780 288808 140808
rect 288802 140768 288808 140780
rect 288860 140768 288866 140820
rect 295702 140740 295708 140752
rect 295663 140712 295708 140740
rect 295702 140700 295708 140712
rect 295760 140700 295766 140752
rect 291562 139340 291568 139392
rect 291620 139380 291626 139392
rect 291746 139380 291752 139392
rect 291620 139352 291752 139380
rect 291620 139340 291626 139352
rect 291746 139340 291752 139352
rect 291804 139340 291810 139392
rect 310793 138703 310851 138709
rect 310793 138669 310805 138703
rect 310839 138700 310851 138703
rect 310882 138700 310888 138712
rect 310839 138672 310888 138700
rect 310839 138669 310851 138672
rect 310793 138663 310851 138669
rect 310882 138660 310888 138672
rect 310940 138660 310946 138712
rect 372709 138159 372767 138165
rect 372709 138125 372721 138159
rect 372755 138156 372767 138159
rect 372798 138156 372804 138168
rect 372755 138128 372804 138156
rect 372755 138125 372767 138128
rect 372709 138119 372767 138125
rect 372798 138116 372804 138128
rect 372856 138116 372862 138168
rect 251450 138020 251456 138032
rect 251411 137992 251456 138020
rect 251450 137980 251456 137992
rect 251508 137980 251514 138032
rect 301038 137980 301044 138032
rect 301096 137980 301102 138032
rect 337102 137980 337108 138032
rect 337160 137980 337166 138032
rect 389358 137980 389364 138032
rect 389416 137980 389422 138032
rect 244458 137952 244464 137964
rect 244419 137924 244464 137952
rect 244458 137912 244464 137924
rect 244516 137912 244522 137964
rect 273530 137952 273536 137964
rect 273491 137924 273536 137952
rect 273530 137912 273536 137924
rect 273588 137912 273594 137964
rect 291565 137955 291623 137961
rect 291565 137921 291577 137955
rect 291611 137952 291623 137955
rect 291746 137952 291752 137964
rect 291611 137924 291752 137952
rect 291611 137921 291623 137924
rect 291565 137915 291623 137921
rect 291746 137912 291752 137924
rect 291804 137912 291810 137964
rect 301056 137952 301084 137980
rect 301130 137952 301136 137964
rect 301056 137924 301136 137952
rect 301130 137912 301136 137924
rect 301188 137912 301194 137964
rect 317506 137912 317512 137964
rect 317564 137952 317570 137964
rect 317782 137952 317788 137964
rect 317564 137924 317788 137952
rect 317564 137912 317570 137924
rect 317782 137912 317788 137924
rect 317840 137912 317846 137964
rect 329926 137912 329932 137964
rect 329984 137952 329990 137964
rect 330202 137952 330208 137964
rect 329984 137924 330208 137952
rect 329984 137912 329990 137924
rect 330202 137912 330208 137924
rect 330260 137912 330266 137964
rect 337120 137952 337148 137980
rect 337194 137952 337200 137964
rect 337120 137924 337200 137952
rect 337194 137912 337200 137924
rect 337252 137912 337258 137964
rect 389376 137952 389404 137980
rect 389450 137952 389456 137964
rect 389376 137924 389456 137952
rect 389450 137912 389456 137924
rect 389508 137912 389514 137964
rect 2774 136484 2780 136536
rect 2832 136524 2838 136536
rect 5074 136524 5080 136536
rect 2832 136496 5080 136524
rect 2832 136484 2838 136496
rect 5074 136484 5080 136496
rect 5132 136484 5138 136536
rect 367002 135300 367008 135312
rect 366963 135272 367008 135300
rect 367002 135260 367008 135272
rect 367060 135260 367066 135312
rect 372706 135300 372712 135312
rect 372667 135272 372712 135300
rect 372706 135260 372712 135272
rect 372764 135260 372770 135312
rect 375834 135300 375840 135312
rect 375795 135272 375840 135300
rect 375834 135260 375840 135272
rect 375892 135260 375898 135312
rect 239122 135192 239128 135244
rect 239180 135232 239186 135244
rect 239306 135232 239312 135244
rect 239180 135204 239312 135232
rect 239180 135192 239186 135204
rect 239306 135192 239312 135204
rect 239364 135192 239370 135244
rect 267734 135192 267740 135244
rect 267792 135232 267798 135244
rect 267826 135232 267832 135244
rect 267792 135204 267832 135232
rect 267792 135192 267798 135204
rect 267826 135192 267832 135204
rect 267884 135192 267890 135244
rect 324590 135192 324596 135244
rect 324648 135232 324654 135244
rect 324682 135232 324688 135244
rect 324648 135204 324688 135232
rect 324648 135192 324654 135204
rect 324682 135192 324688 135204
rect 324740 135192 324746 135244
rect 327258 135232 327264 135244
rect 327219 135204 327264 135232
rect 327258 135192 327264 135204
rect 327316 135192 327322 135244
rect 340874 135192 340880 135244
rect 340932 135232 340938 135244
rect 341242 135232 341248 135244
rect 340932 135204 341248 135232
rect 340932 135192 340938 135204
rect 341242 135192 341248 135204
rect 341300 135192 341306 135244
rect 357434 135192 357440 135244
rect 357492 135232 357498 135244
rect 357492 135204 357537 135232
rect 357492 135192 357498 135204
rect 470410 135192 470416 135244
rect 470468 135232 470474 135244
rect 470594 135232 470600 135244
rect 470468 135204 470600 135232
rect 470468 135192 470474 135204
rect 470594 135192 470600 135204
rect 470652 135192 470658 135244
rect 270954 135096 270960 135108
rect 270915 135068 270960 135096
rect 270954 135056 270960 135068
rect 271012 135056 271018 135108
rect 251450 133940 251456 133952
rect 251411 133912 251456 133940
rect 251450 133900 251456 133912
rect 251508 133900 251514 133952
rect 358722 133900 358728 133952
rect 358780 133940 358786 133952
rect 421190 133940 421196 133952
rect 358780 133912 358825 133940
rect 421151 133912 421196 133940
rect 358780 133900 358786 133912
rect 421190 133900 421196 133912
rect 421248 133900 421254 133952
rect 337194 133872 337200 133884
rect 337155 133844 337200 133872
rect 337194 133832 337200 133844
rect 337252 133832 337258 133884
rect 389450 133872 389456 133884
rect 389411 133844 389456 133872
rect 389450 133832 389456 133844
rect 389508 133832 389514 133884
rect 249978 132512 249984 132524
rect 249939 132484 249984 132512
rect 249978 132472 249984 132484
rect 250036 132472 250042 132524
rect 259641 132515 259699 132521
rect 259641 132481 259653 132515
rect 259687 132512 259699 132515
rect 259730 132512 259736 132524
rect 259687 132484 259736 132512
rect 259687 132481 259699 132484
rect 259641 132475 259699 132481
rect 259730 132472 259736 132484
rect 259788 132472 259794 132524
rect 286042 132512 286048 132524
rect 286003 132484 286048 132512
rect 286042 132472 286048 132484
rect 286100 132472 286106 132524
rect 296898 132512 296904 132524
rect 296859 132484 296904 132512
rect 296898 132472 296904 132484
rect 296956 132472 296962 132524
rect 299750 132472 299756 132524
rect 299808 132512 299814 132524
rect 299842 132512 299848 132524
rect 299808 132484 299848 132512
rect 299808 132472 299814 132484
rect 299842 132472 299848 132484
rect 299900 132472 299906 132524
rect 302418 132472 302424 132524
rect 302476 132512 302482 132524
rect 302602 132512 302608 132524
rect 302476 132484 302608 132512
rect 302476 132472 302482 132484
rect 302602 132472 302608 132484
rect 302660 132472 302666 132524
rect 284662 132444 284668 132456
rect 284623 132416 284668 132444
rect 284662 132404 284668 132416
rect 284720 132404 284726 132456
rect 306742 132444 306748 132456
rect 306703 132416 306748 132444
rect 306742 132404 306748 132416
rect 306800 132404 306806 132456
rect 288802 131220 288808 131232
rect 288728 131192 288808 131220
rect 288728 131164 288756 131192
rect 288802 131180 288808 131192
rect 288860 131180 288866 131232
rect 288710 131112 288716 131164
rect 288768 131112 288774 131164
rect 295610 131112 295616 131164
rect 295668 131152 295674 131164
rect 295705 131155 295763 131161
rect 295705 131152 295717 131155
rect 295668 131124 295717 131152
rect 295668 131112 295674 131124
rect 295705 131121 295717 131124
rect 295751 131121 295763 131155
rect 295705 131115 295763 131121
rect 463878 130364 463884 130416
rect 463936 130404 463942 130416
rect 464062 130404 464068 130416
rect 463936 130376 464068 130404
rect 463936 130364 463942 130376
rect 464062 130364 464068 130376
rect 464120 130364 464126 130416
rect 306745 129931 306803 129937
rect 306745 129897 306757 129931
rect 306791 129928 306803 129931
rect 306834 129928 306840 129940
rect 306791 129900 306840 129928
rect 306791 129897 306803 129900
rect 306745 129891 306803 129897
rect 306834 129888 306840 129900
rect 306892 129888 306898 129940
rect 325970 128432 325976 128444
rect 325896 128404 325976 128432
rect 325896 128308 325924 128404
rect 325970 128392 325976 128404
rect 326028 128392 326034 128444
rect 339678 128324 339684 128376
rect 339736 128364 339742 128376
rect 339862 128364 339868 128376
rect 339736 128336 339868 128364
rect 339736 128324 339742 128336
rect 339862 128324 339868 128336
rect 339920 128324 339926 128376
rect 360286 128324 360292 128376
rect 360344 128364 360350 128376
rect 360470 128364 360476 128376
rect 360344 128336 360476 128364
rect 360344 128324 360350 128336
rect 360470 128324 360476 128336
rect 360528 128324 360534 128376
rect 424134 128324 424140 128376
rect 424192 128364 424198 128376
rect 424502 128364 424508 128376
rect 424192 128336 424508 128364
rect 424192 128324 424198 128336
rect 424502 128324 424508 128336
rect 424560 128324 424566 128376
rect 310790 128296 310796 128308
rect 310751 128268 310796 128296
rect 310790 128256 310796 128268
rect 310848 128256 310854 128308
rect 325878 128256 325884 128308
rect 325936 128256 325942 128308
rect 357437 128231 357495 128237
rect 357437 128197 357449 128231
rect 357483 128228 357495 128231
rect 357526 128228 357532 128240
rect 357483 128200 357532 128228
rect 357483 128197 357495 128200
rect 357437 128191 357495 128197
rect 357526 128188 357532 128200
rect 357584 128188 357590 128240
rect 232314 125712 232320 125724
rect 232275 125684 232320 125712
rect 232314 125672 232320 125684
rect 232372 125672 232378 125724
rect 265158 125536 265164 125588
rect 265216 125576 265222 125588
rect 265342 125576 265348 125588
rect 265216 125548 265348 125576
rect 265216 125536 265222 125548
rect 265342 125536 265348 125548
rect 265400 125536 265406 125588
rect 267734 125536 267740 125588
rect 267792 125576 267798 125588
rect 267918 125576 267924 125588
rect 267792 125548 267924 125576
rect 267792 125536 267798 125548
rect 267918 125536 267924 125548
rect 267976 125536 267982 125588
rect 270678 125536 270684 125588
rect 270736 125576 270742 125588
rect 270954 125576 270960 125588
rect 270736 125548 270960 125576
rect 270736 125536 270742 125548
rect 270954 125536 270960 125548
rect 271012 125536 271018 125588
rect 272150 125536 272156 125588
rect 272208 125576 272214 125588
rect 272426 125576 272432 125588
rect 272208 125548 272432 125576
rect 272208 125536 272214 125548
rect 272426 125536 272432 125548
rect 272484 125536 272490 125588
rect 273530 125576 273536 125588
rect 273491 125548 273536 125576
rect 273530 125536 273536 125548
rect 273588 125536 273594 125588
rect 323210 125536 323216 125588
rect 323268 125576 323274 125588
rect 323394 125576 323400 125588
rect 323268 125548 323400 125576
rect 323268 125536 323274 125548
rect 323394 125536 323400 125548
rect 323452 125536 323458 125588
rect 324590 125536 324596 125588
rect 324648 125576 324654 125588
rect 324774 125576 324780 125588
rect 324648 125548 324780 125576
rect 324648 125536 324654 125548
rect 324774 125536 324780 125548
rect 324832 125536 324838 125588
rect 325878 125536 325884 125588
rect 325936 125576 325942 125588
rect 326062 125576 326068 125588
rect 325936 125548 326068 125576
rect 325936 125536 325942 125548
rect 326062 125536 326068 125548
rect 326120 125536 326126 125588
rect 327166 125536 327172 125588
rect 327224 125536 327230 125588
rect 341058 125536 341064 125588
rect 341116 125576 341122 125588
rect 341153 125579 341211 125585
rect 341153 125576 341165 125579
rect 341116 125548 341165 125576
rect 341116 125536 341122 125548
rect 341153 125545 341165 125548
rect 341199 125545 341211 125579
rect 341153 125539 341211 125545
rect 357526 125536 357532 125588
rect 357584 125536 357590 125588
rect 367002 125576 367008 125588
rect 366963 125548 367008 125576
rect 367002 125536 367008 125548
rect 367060 125536 367066 125588
rect 310793 125511 310851 125517
rect 310793 125477 310805 125511
rect 310839 125508 310851 125511
rect 310882 125508 310888 125520
rect 310839 125480 310888 125508
rect 310839 125477 310851 125480
rect 310793 125471 310851 125477
rect 310882 125468 310888 125480
rect 310940 125468 310946 125520
rect 327184 125508 327212 125536
rect 327258 125508 327264 125520
rect 327184 125480 327264 125508
rect 327258 125468 327264 125480
rect 327316 125468 327322 125520
rect 357544 125508 357572 125536
rect 357618 125508 357624 125520
rect 357544 125480 357624 125508
rect 357618 125468 357624 125480
rect 357676 125468 357682 125520
rect 337197 124219 337255 124225
rect 337197 124185 337209 124219
rect 337243 124216 337255 124219
rect 337286 124216 337292 124228
rect 337243 124188 337292 124216
rect 337243 124185 337255 124188
rect 337197 124179 337255 124185
rect 337286 124176 337292 124188
rect 337344 124176 337350 124228
rect 232314 124148 232320 124160
rect 232275 124120 232320 124148
rect 232314 124108 232320 124120
rect 232372 124108 232378 124160
rect 249978 124148 249984 124160
rect 249939 124120 249984 124148
rect 249978 124108 249984 124120
rect 250036 124108 250042 124160
rect 272153 124151 272211 124157
rect 272153 124117 272165 124151
rect 272199 124148 272211 124151
rect 272426 124148 272432 124160
rect 272199 124120 272432 124148
rect 272199 124117 272211 124120
rect 272153 124111 272211 124117
rect 272426 124108 272432 124120
rect 272484 124108 272490 124160
rect 358722 124148 358728 124160
rect 358683 124120 358728 124148
rect 358722 124108 358728 124120
rect 358780 124108 358786 124160
rect 421190 124148 421196 124160
rect 421151 124120 421196 124148
rect 421190 124108 421196 124120
rect 421248 124108 421254 124160
rect 284665 122859 284723 122865
rect 284665 122825 284677 122859
rect 284711 122856 284723 122859
rect 284846 122856 284852 122868
rect 284711 122828 284852 122856
rect 284711 122825 284723 122828
rect 284665 122819 284723 122825
rect 284846 122816 284852 122828
rect 284904 122816 284910 122868
rect 289998 122816 290004 122868
rect 290056 122816 290062 122868
rect 296898 122816 296904 122868
rect 296956 122856 296962 122868
rect 297082 122856 297088 122868
rect 296956 122828 297088 122856
rect 296956 122816 296962 122828
rect 297082 122816 297088 122828
rect 297140 122816 297146 122868
rect 389174 122816 389180 122868
rect 389232 122856 389238 122868
rect 389453 122859 389511 122865
rect 389453 122856 389465 122859
rect 389232 122828 389465 122856
rect 389232 122816 389238 122828
rect 389453 122825 389465 122828
rect 389499 122825 389511 122859
rect 389453 122819 389511 122825
rect 290016 122720 290044 122816
rect 290090 122720 290096 122732
rect 290016 122692 290096 122720
rect 290090 122680 290096 122692
rect 290148 122680 290154 122732
rect 2774 122272 2780 122324
rect 2832 122312 2838 122324
rect 4982 122312 4988 122324
rect 2832 122284 4988 122312
rect 2832 122272 2838 122284
rect 4982 122272 4988 122284
rect 5040 122272 5046 122324
rect 306834 121388 306840 121440
rect 306892 121388 306898 121440
rect 330202 121388 330208 121440
rect 330260 121428 330266 121440
rect 330570 121428 330576 121440
rect 330260 121400 330576 121428
rect 330260 121388 330266 121400
rect 330570 121388 330576 121400
rect 330628 121388 330634 121440
rect 306852 121301 306880 121388
rect 306837 121295 306895 121301
rect 306837 121261 306849 121295
rect 306883 121261 306895 121295
rect 306837 121255 306895 121261
rect 324593 120615 324651 120621
rect 324593 120581 324605 120615
rect 324639 120612 324651 120615
rect 324774 120612 324780 120624
rect 324639 120584 324780 120612
rect 324639 120581 324651 120584
rect 324593 120575 324651 120581
rect 324774 120572 324780 120584
rect 324832 120572 324838 120624
rect 291562 120136 291568 120148
rect 291523 120108 291568 120136
rect 291562 120096 291568 120108
rect 291620 120096 291626 120148
rect 330570 120068 330576 120080
rect 330531 120040 330576 120068
rect 330570 120028 330576 120040
rect 330628 120028 330634 120080
rect 251450 118736 251456 118788
rect 251508 118736 251514 118788
rect 299842 118736 299848 118788
rect 299900 118736 299906 118788
rect 339773 118779 339831 118785
rect 339773 118745 339785 118779
rect 339819 118776 339831 118779
rect 339862 118776 339868 118788
rect 339819 118748 339868 118776
rect 339819 118745 339831 118748
rect 339773 118739 339831 118745
rect 339862 118736 339868 118748
rect 339920 118736 339926 118788
rect 251468 118652 251496 118736
rect 299860 118652 299888 118736
rect 337102 118668 337108 118720
rect 337160 118708 337166 118720
rect 337286 118708 337292 118720
rect 337160 118680 337292 118708
rect 337160 118668 337166 118680
rect 337286 118668 337292 118680
rect 337344 118668 337350 118720
rect 377122 118668 377128 118720
rect 377180 118668 377186 118720
rect 463878 118668 463884 118720
rect 463936 118668 463942 118720
rect 251450 118600 251456 118652
rect 251508 118600 251514 118652
rect 299842 118600 299848 118652
rect 299900 118600 299906 118652
rect 341150 118640 341156 118652
rect 341111 118612 341156 118640
rect 341150 118600 341156 118612
rect 341208 118600 341214 118652
rect 377140 118584 377168 118668
rect 463896 118640 463924 118668
rect 463970 118640 463976 118652
rect 463896 118612 463976 118640
rect 463970 118600 463976 118612
rect 464028 118600 464034 118652
rect 377122 118532 377128 118584
rect 377180 118532 377186 118584
rect 326062 118396 326068 118448
rect 326120 118396 326126 118448
rect 326080 118312 326108 118396
rect 326062 118260 326068 118312
rect 326120 118260 326126 118312
rect 273530 115988 273536 116000
rect 273491 115960 273536 115988
rect 273530 115948 273536 115960
rect 273588 115948 273594 116000
rect 339770 115988 339776 116000
rect 339731 115960 339776 115988
rect 339770 115948 339776 115960
rect 339828 115948 339834 116000
rect 367002 115988 367008 116000
rect 366963 115960 367008 115988
rect 367002 115948 367008 115960
rect 367060 115948 367066 116000
rect 270678 115880 270684 115932
rect 270736 115920 270742 115932
rect 270954 115920 270960 115932
rect 270736 115892 270960 115920
rect 270736 115880 270742 115892
rect 270954 115880 270960 115892
rect 271012 115880 271018 115932
rect 341242 115880 341248 115932
rect 341300 115920 341306 115932
rect 341426 115920 341432 115932
rect 341300 115892 341432 115920
rect 341300 115880 341306 115892
rect 341426 115880 341432 115892
rect 341484 115880 341490 115932
rect 377033 115923 377091 115929
rect 377033 115889 377045 115923
rect 377079 115920 377091 115923
rect 377122 115920 377128 115932
rect 377079 115892 377128 115920
rect 377079 115889 377091 115892
rect 377033 115883 377091 115889
rect 377122 115880 377128 115892
rect 377180 115880 377186 115932
rect 424594 115880 424600 115932
rect 424652 115920 424658 115932
rect 424686 115920 424692 115932
rect 424652 115892 424692 115920
rect 424652 115880 424658 115892
rect 424686 115880 424692 115892
rect 424744 115880 424750 115932
rect 366818 115812 366824 115864
rect 366876 115852 366882 115864
rect 367002 115852 367008 115864
rect 366876 115824 367008 115852
rect 366876 115812 366882 115824
rect 367002 115812 367008 115824
rect 367060 115812 367066 115864
rect 291473 115243 291531 115249
rect 291473 115209 291485 115243
rect 291519 115240 291531 115243
rect 291562 115240 291568 115252
rect 291519 115212 291568 115240
rect 291519 115209 291531 115212
rect 291473 115203 291531 115209
rect 291562 115200 291568 115212
rect 291620 115200 291626 115252
rect 310793 114631 310851 114637
rect 310793 114597 310805 114631
rect 310839 114628 310851 114631
rect 310882 114628 310888 114640
rect 310839 114600 310888 114628
rect 310839 114597 310851 114600
rect 310793 114591 310851 114597
rect 310882 114588 310888 114600
rect 310940 114588 310946 114640
rect 232314 114560 232320 114572
rect 232275 114532 232320 114560
rect 232314 114520 232320 114532
rect 232372 114520 232378 114572
rect 249981 114563 250039 114569
rect 249981 114529 249993 114563
rect 250027 114560 250039 114563
rect 250254 114560 250260 114572
rect 250027 114532 250260 114560
rect 250027 114529 250039 114532
rect 249981 114523 250039 114529
rect 250254 114520 250260 114532
rect 250312 114520 250318 114572
rect 272150 114560 272156 114572
rect 272111 114532 272156 114560
rect 272150 114520 272156 114532
rect 272208 114520 272214 114572
rect 358722 114560 358728 114572
rect 358683 114532 358728 114560
rect 358722 114520 358728 114532
rect 358780 114520 358786 114572
rect 421190 114560 421196 114572
rect 421151 114532 421196 114560
rect 421190 114520 421196 114532
rect 421248 114520 421254 114572
rect 267826 114492 267832 114504
rect 267787 114464 267832 114492
rect 267826 114452 267832 114464
rect 267884 114452 267890 114504
rect 285950 114452 285956 114504
rect 286008 114492 286014 114504
rect 286226 114492 286232 114504
rect 286008 114464 286232 114492
rect 286008 114452 286014 114464
rect 286226 114452 286232 114464
rect 286284 114452 286290 114504
rect 310790 114492 310796 114504
rect 310751 114464 310796 114492
rect 310790 114452 310796 114464
rect 310848 114452 310854 114504
rect 424505 114495 424563 114501
rect 424505 114461 424517 114495
rect 424551 114492 424563 114495
rect 424594 114492 424600 114504
rect 424551 114464 424600 114492
rect 424551 114461 424563 114464
rect 424505 114455 424563 114461
rect 424594 114452 424600 114464
rect 424652 114452 424658 114504
rect 301038 113228 301044 113280
rect 301096 113228 301102 113280
rect 259638 113160 259644 113212
rect 259696 113200 259702 113212
rect 259730 113200 259736 113212
rect 259696 113172 259736 113200
rect 259696 113160 259702 113172
rect 259730 113160 259736 113172
rect 259788 113160 259794 113212
rect 296990 113160 296996 113212
rect 297048 113200 297054 113212
rect 297082 113200 297088 113212
rect 297048 113172 297088 113200
rect 297048 113160 297054 113172
rect 297082 113160 297088 113172
rect 297140 113160 297146 113212
rect 301056 113200 301084 113228
rect 301130 113200 301136 113212
rect 301056 113172 301136 113200
rect 301130 113160 301136 113172
rect 301188 113160 301194 113212
rect 324590 113200 324596 113212
rect 324551 113172 324596 113200
rect 324590 113160 324596 113172
rect 324648 113160 324654 113212
rect 267829 113135 267887 113141
rect 267829 113101 267841 113135
rect 267875 113132 267887 113135
rect 268013 113135 268071 113141
rect 268013 113132 268025 113135
rect 267875 113104 268025 113132
rect 267875 113101 267887 113104
rect 267829 113095 267887 113101
rect 268013 113101 268025 113104
rect 268059 113101 268071 113135
rect 268013 113095 268071 113101
rect 299842 113092 299848 113144
rect 299900 113132 299906 113144
rect 299934 113132 299940 113144
rect 299900 113104 299940 113132
rect 299900 113092 299906 113104
rect 299934 113092 299940 113104
rect 299992 113092 299998 113144
rect 306834 111840 306840 111852
rect 306795 111812 306840 111840
rect 306834 111800 306840 111812
rect 306892 111800 306898 111852
rect 330570 111772 330576 111784
rect 330531 111744 330576 111772
rect 330570 111732 330576 111744
rect 330628 111732 330634 111784
rect 368198 110644 368204 110696
rect 368256 110684 368262 110696
rect 376662 110684 376668 110696
rect 368256 110656 376668 110684
rect 368256 110644 368262 110656
rect 376662 110644 376668 110656
rect 376720 110644 376726 110696
rect 456518 110644 456524 110696
rect 456576 110684 456582 110696
rect 458818 110684 458824 110696
rect 456576 110656 458824 110684
rect 456576 110644 456582 110656
rect 458818 110644 458824 110656
rect 458876 110644 458882 110696
rect 414014 110576 414020 110628
rect 414072 110616 414078 110628
rect 423490 110616 423496 110628
rect 414072 110588 423496 110616
rect 414072 110576 414078 110588
rect 423490 110576 423496 110588
rect 423548 110576 423554 110628
rect 437198 110576 437204 110628
rect 437256 110616 437262 110628
rect 437474 110616 437480 110628
rect 437256 110588 437480 110616
rect 437256 110576 437262 110588
rect 437474 110576 437480 110588
rect 437532 110576 437538 110628
rect 347774 110508 347780 110560
rect 347832 110548 347838 110560
rect 357342 110548 357348 110560
rect 347832 110520 357348 110548
rect 347832 110508 347838 110520
rect 357342 110508 357348 110520
rect 357400 110508 357406 110560
rect 324590 109692 324596 109744
rect 324648 109692 324654 109744
rect 324608 109608 324636 109692
rect 324590 109556 324596 109608
rect 324648 109556 324654 109608
rect 362218 109120 362224 109132
rect 362144 109092 362224 109120
rect 266630 109012 266636 109064
rect 266688 109012 266694 109064
rect 266648 108984 266676 109012
rect 362144 108996 362172 109092
rect 362218 109080 362224 109092
rect 362276 109080 362282 109132
rect 463786 109012 463792 109064
rect 463844 109052 463850 109064
rect 463970 109052 463976 109064
rect 463844 109024 463976 109052
rect 463844 109012 463850 109024
rect 463970 109012 463976 109024
rect 464028 109012 464034 109064
rect 266722 108984 266728 108996
rect 266648 108956 266728 108984
rect 266722 108944 266728 108956
rect 266780 108944 266786 108996
rect 278774 108944 278780 108996
rect 278832 108984 278838 108996
rect 279050 108984 279056 108996
rect 278832 108956 279056 108984
rect 278832 108944 278838 108956
rect 279050 108944 279056 108956
rect 279108 108944 279114 108996
rect 362126 108944 362132 108996
rect 362184 108944 362190 108996
rect 330205 106743 330263 106749
rect 330205 106709 330217 106743
rect 330251 106740 330263 106743
rect 330570 106740 330576 106752
rect 330251 106712 330576 106740
rect 330251 106709 330263 106712
rect 330205 106703 330263 106709
rect 330570 106700 330576 106712
rect 330628 106700 330634 106752
rect 284846 106332 284852 106344
rect 284772 106304 284852 106332
rect 284772 106276 284800 106304
rect 284846 106292 284852 106304
rect 284904 106292 284910 106344
rect 358722 106332 358728 106344
rect 358683 106304 358728 106332
rect 358722 106292 358728 106304
rect 358780 106292 358786 106344
rect 377030 106332 377036 106344
rect 376991 106304 377036 106332
rect 377030 106292 377036 106304
rect 377088 106292 377094 106344
rect 236454 106224 236460 106276
rect 236512 106264 236518 106276
rect 236638 106264 236644 106276
rect 236512 106236 236644 106264
rect 236512 106224 236518 106236
rect 236638 106224 236644 106236
rect 236696 106224 236702 106276
rect 239122 106224 239128 106276
rect 239180 106264 239186 106276
rect 239306 106264 239312 106276
rect 239180 106236 239312 106264
rect 239180 106224 239186 106236
rect 239306 106224 239312 106236
rect 239364 106224 239370 106276
rect 259546 106224 259552 106276
rect 259604 106264 259610 106276
rect 259822 106264 259828 106276
rect 259604 106236 259828 106264
rect 259604 106224 259610 106236
rect 259822 106224 259828 106236
rect 259880 106224 259886 106276
rect 270678 106224 270684 106276
rect 270736 106264 270742 106276
rect 270954 106264 270960 106276
rect 270736 106236 270960 106264
rect 270736 106224 270742 106236
rect 270954 106224 270960 106236
rect 271012 106224 271018 106276
rect 272150 106224 272156 106276
rect 272208 106264 272214 106276
rect 272426 106264 272432 106276
rect 272208 106236 272432 106264
rect 272208 106224 272214 106236
rect 272426 106224 272432 106236
rect 272484 106224 272490 106276
rect 273530 106264 273536 106276
rect 273491 106236 273536 106264
rect 273530 106224 273536 106236
rect 273588 106224 273594 106276
rect 284754 106224 284760 106276
rect 284812 106224 284818 106276
rect 375834 106264 375840 106276
rect 375795 106236 375840 106264
rect 375834 106224 375840 106236
rect 375892 106224 375898 106276
rect 377122 106264 377128 106276
rect 377083 106236 377128 106264
rect 377122 106224 377128 106236
rect 377180 106224 377186 106276
rect 358722 104972 358728 104984
rect 358683 104944 358728 104972
rect 358722 104932 358728 104944
rect 358780 104932 358786 104984
rect 265250 104864 265256 104916
rect 265308 104904 265314 104916
rect 265342 104904 265348 104916
rect 265308 104876 265348 104904
rect 265308 104864 265314 104876
rect 265342 104864 265348 104876
rect 265400 104864 265406 104916
rect 288802 104864 288808 104916
rect 288860 104904 288866 104916
rect 288986 104904 288992 104916
rect 288860 104876 288992 104904
rect 288860 104864 288866 104876
rect 288986 104864 288992 104876
rect 289044 104864 289050 104916
rect 310793 104907 310851 104913
rect 310793 104873 310805 104907
rect 310839 104904 310851 104907
rect 310882 104904 310888 104916
rect 310839 104876 310888 104904
rect 310839 104873 310851 104876
rect 310793 104867 310851 104873
rect 310882 104864 310888 104876
rect 310940 104864 310946 104916
rect 424502 104904 424508 104916
rect 424463 104876 424508 104904
rect 424502 104864 424508 104876
rect 424560 104864 424566 104916
rect 232314 104836 232320 104848
rect 232275 104808 232320 104836
rect 232314 104796 232320 104808
rect 232372 104796 232378 104848
rect 295518 104796 295524 104848
rect 295576 104836 295582 104848
rect 295610 104836 295616 104848
rect 295576 104808 295616 104836
rect 295576 104796 295582 104808
rect 295610 104796 295616 104808
rect 295668 104796 295674 104848
rect 302602 104836 302608 104848
rect 302563 104808 302608 104836
rect 302602 104796 302608 104808
rect 302660 104796 302666 104848
rect 323394 104836 323400 104848
rect 323355 104808 323400 104836
rect 323394 104796 323400 104808
rect 323452 104796 323458 104848
rect 324590 104836 324596 104848
rect 324551 104808 324596 104836
rect 324590 104796 324596 104808
rect 324648 104796 324654 104848
rect 337197 104839 337255 104845
rect 337197 104805 337209 104839
rect 337243 104836 337255 104839
rect 337286 104836 337292 104848
rect 337243 104808 337292 104836
rect 337243 104805 337255 104808
rect 337197 104799 337255 104805
rect 337286 104796 337292 104808
rect 337344 104796 337350 104848
rect 339494 104796 339500 104848
rect 339552 104836 339558 104848
rect 339770 104836 339776 104848
rect 339552 104808 339776 104836
rect 339552 104796 339558 104808
rect 339770 104796 339776 104808
rect 339828 104796 339834 104848
rect 358633 104839 358691 104845
rect 358633 104805 358645 104839
rect 358679 104836 358691 104839
rect 358722 104836 358728 104848
rect 358679 104808 358728 104836
rect 358679 104805 358691 104808
rect 358633 104799 358691 104805
rect 358722 104796 358728 104808
rect 358780 104796 358786 104848
rect 421190 104836 421196 104848
rect 421151 104808 421196 104836
rect 421190 104796 421196 104808
rect 421248 104796 421254 104848
rect 268013 103615 268071 103621
rect 268013 103612 268025 103615
rect 267844 103584 268025 103612
rect 267844 103485 267872 103584
rect 268013 103581 268025 103584
rect 268059 103581 268071 103615
rect 268013 103575 268071 103581
rect 291470 103544 291476 103556
rect 291431 103516 291476 103544
rect 291470 103504 291476 103516
rect 291528 103504 291534 103556
rect 267829 103479 267887 103485
rect 267829 103445 267841 103479
rect 267875 103445 267887 103479
rect 267829 103439 267887 103445
rect 272426 103436 272432 103488
rect 272484 103476 272490 103488
rect 327166 103476 327172 103488
rect 272484 103448 272529 103476
rect 327127 103448 327172 103476
rect 272484 103436 272490 103448
rect 327166 103436 327172 103448
rect 327224 103436 327230 103488
rect 339405 103479 339463 103485
rect 339405 103445 339417 103479
rect 339451 103476 339463 103479
rect 339494 103476 339500 103488
rect 339451 103448 339500 103476
rect 339451 103445 339463 103448
rect 339405 103439 339463 103445
rect 339494 103436 339500 103448
rect 339552 103436 339558 103488
rect 330202 102184 330208 102196
rect 330163 102156 330208 102184
rect 330202 102144 330208 102156
rect 330260 102144 330266 102196
rect 288713 102119 288771 102125
rect 288713 102085 288725 102119
rect 288759 102116 288771 102119
rect 288802 102116 288808 102128
rect 288759 102088 288808 102116
rect 288759 102085 288771 102088
rect 288713 102079 288771 102085
rect 288802 102076 288808 102088
rect 288860 102076 288866 102128
rect 294230 100036 294236 100088
rect 294288 100076 294294 100088
rect 294414 100076 294420 100088
rect 294288 100048 294420 100076
rect 294288 100036 294294 100048
rect 294414 100036 294420 100048
rect 294472 100036 294478 100088
rect 244458 99424 244464 99476
rect 244516 99424 244522 99476
rect 245930 99424 245936 99476
rect 245988 99424 245994 99476
rect 310882 99424 310888 99476
rect 310940 99424 310946 99476
rect 244476 99340 244504 99424
rect 245948 99340 245976 99424
rect 251450 99396 251456 99408
rect 251411 99368 251456 99396
rect 251450 99356 251456 99368
rect 251508 99356 251514 99408
rect 278866 99356 278872 99408
rect 278924 99396 278930 99408
rect 279050 99396 279056 99408
rect 278924 99368 279056 99396
rect 278924 99356 278930 99368
rect 279050 99356 279056 99368
rect 279108 99356 279114 99408
rect 310900 99340 310928 99424
rect 424502 99356 424508 99408
rect 424560 99356 424566 99408
rect 244458 99288 244464 99340
rect 244516 99288 244522 99340
rect 245930 99288 245936 99340
rect 245988 99288 245994 99340
rect 273530 99328 273536 99340
rect 273491 99300 273536 99328
rect 273530 99288 273536 99300
rect 273588 99288 273594 99340
rect 310882 99288 310888 99340
rect 310940 99288 310946 99340
rect 377122 99328 377128 99340
rect 377083 99300 377128 99328
rect 377122 99288 377128 99300
rect 377180 99288 377186 99340
rect 424520 99328 424548 99356
rect 424686 99328 424692 99340
rect 424520 99300 424692 99328
rect 424686 99288 424692 99300
rect 424744 99288 424750 99340
rect 389361 99195 389419 99201
rect 389361 99161 389373 99195
rect 389407 99192 389419 99195
rect 389450 99192 389456 99204
rect 389407 99164 389456 99192
rect 389407 99161 389419 99164
rect 389361 99155 389419 99161
rect 389450 99152 389456 99164
rect 389508 99152 389514 99204
rect 327166 98716 327172 98728
rect 327127 98688 327172 98716
rect 327166 98676 327172 98688
rect 327224 98676 327230 98728
rect 270494 98064 270500 98116
rect 270552 98104 270558 98116
rect 270954 98104 270960 98116
rect 270552 98076 270960 98104
rect 270552 98064 270558 98076
rect 270954 98064 270960 98076
rect 271012 98064 271018 98116
rect 375834 97832 375840 97844
rect 375795 97804 375840 97832
rect 375834 97792 375840 97804
rect 375892 97792 375898 97844
rect 330113 97291 330171 97297
rect 330113 97257 330125 97291
rect 330159 97288 330171 97291
rect 330202 97288 330208 97300
rect 330159 97260 330208 97288
rect 330159 97257 330171 97260
rect 330113 97251 330171 97257
rect 330202 97248 330208 97260
rect 330260 97248 330266 97300
rect 250070 96636 250076 96688
rect 250128 96676 250134 96688
rect 250254 96676 250260 96688
rect 250128 96648 250260 96676
rect 250128 96636 250134 96648
rect 250254 96636 250260 96648
rect 250312 96636 250318 96688
rect 251450 96676 251456 96688
rect 251411 96648 251456 96676
rect 251450 96636 251456 96648
rect 251508 96636 251514 96688
rect 367002 96608 367008 96620
rect 366963 96580 367008 96608
rect 367002 96568 367008 96580
rect 367060 96568 367066 96620
rect 372614 96568 372620 96620
rect 372672 96608 372678 96620
rect 372706 96608 372712 96620
rect 372672 96580 372712 96608
rect 372672 96568 372678 96580
rect 372706 96568 372712 96580
rect 372764 96568 372770 96620
rect 232314 95248 232320 95260
rect 232275 95220 232320 95248
rect 232314 95208 232320 95220
rect 232372 95208 232378 95260
rect 285950 95208 285956 95260
rect 286008 95248 286014 95260
rect 286042 95248 286048 95260
rect 286008 95220 286048 95248
rect 286008 95208 286014 95220
rect 286042 95208 286048 95220
rect 286100 95208 286106 95260
rect 302602 95248 302608 95260
rect 302563 95220 302608 95248
rect 302602 95208 302608 95220
rect 302660 95208 302666 95260
rect 323394 95248 323400 95260
rect 323355 95220 323400 95248
rect 323394 95208 323400 95220
rect 323452 95208 323458 95260
rect 324590 95248 324596 95260
rect 324551 95220 324596 95248
rect 324590 95208 324596 95220
rect 324648 95208 324654 95260
rect 325878 95208 325884 95260
rect 325936 95248 325942 95260
rect 325970 95248 325976 95260
rect 325936 95220 325976 95248
rect 325936 95208 325942 95220
rect 325970 95208 325976 95220
rect 326028 95208 326034 95260
rect 337194 95248 337200 95260
rect 337155 95220 337200 95248
rect 337194 95208 337200 95220
rect 337252 95208 337258 95260
rect 339405 95251 339463 95257
rect 339405 95217 339417 95251
rect 339451 95248 339463 95251
rect 339494 95248 339500 95260
rect 339451 95220 339500 95248
rect 339451 95217 339463 95220
rect 339405 95211 339463 95217
rect 339494 95208 339500 95220
rect 339552 95208 339558 95260
rect 358630 95248 358636 95260
rect 358591 95220 358636 95248
rect 358630 95208 358636 95220
rect 358688 95208 358694 95260
rect 266630 95180 266636 95192
rect 266591 95152 266636 95180
rect 266630 95140 266636 95152
rect 266688 95140 266694 95192
rect 284754 95180 284760 95192
rect 284715 95152 284760 95180
rect 284754 95140 284760 95152
rect 284812 95140 284818 95192
rect 310790 95180 310796 95192
rect 310751 95152 310796 95180
rect 310790 95140 310796 95152
rect 310848 95140 310854 95192
rect 362310 95180 362316 95192
rect 362271 95152 362316 95180
rect 362310 95140 362316 95152
rect 362368 95140 362374 95192
rect 267734 93848 267740 93900
rect 267792 93888 267798 93900
rect 267829 93891 267887 93897
rect 267829 93888 267841 93891
rect 267792 93860 267841 93888
rect 267792 93848 267798 93860
rect 267829 93857 267841 93860
rect 267875 93857 267887 93891
rect 267829 93851 267887 93857
rect 272334 93848 272340 93900
rect 272392 93888 272398 93900
rect 272429 93891 272487 93897
rect 272429 93888 272441 93891
rect 272392 93860 272441 93888
rect 272392 93848 272398 93860
rect 272429 93857 272441 93860
rect 272475 93857 272487 93891
rect 284754 93888 284760 93900
rect 284715 93860 284760 93888
rect 272429 93851 272487 93857
rect 284754 93848 284760 93860
rect 284812 93848 284818 93900
rect 463694 93848 463700 93900
rect 463752 93888 463758 93900
rect 463878 93888 463884 93900
rect 463752 93860 463884 93888
rect 463752 93848 463758 93860
rect 463878 93848 463884 93860
rect 463936 93848 463942 93900
rect 291381 93823 291439 93829
rect 291381 93789 291393 93823
rect 291427 93820 291439 93823
rect 291470 93820 291476 93832
rect 291427 93792 291476 93820
rect 291427 93789 291439 93792
rect 291381 93783 291439 93789
rect 291470 93780 291476 93792
rect 291528 93780 291534 93832
rect 306834 92596 306840 92608
rect 306760 92568 306840 92596
rect 306760 92540 306788 92568
rect 306834 92556 306840 92568
rect 306892 92556 306898 92608
rect 288710 92528 288716 92540
rect 288671 92500 288716 92528
rect 288710 92488 288716 92500
rect 288768 92488 288774 92540
rect 306742 92488 306748 92540
rect 306800 92488 306806 92540
rect 317782 89700 317788 89752
rect 317840 89700 317846 89752
rect 424502 89700 424508 89752
rect 424560 89740 424566 89752
rect 424686 89740 424692 89752
rect 424560 89712 424692 89740
rect 424560 89700 424566 89712
rect 424686 89700 424692 89712
rect 424744 89700 424750 89752
rect 317800 89604 317828 89700
rect 317874 89604 317880 89616
rect 317800 89576 317880 89604
rect 317874 89564 317880 89576
rect 317932 89564 317938 89616
rect 291378 88992 291384 89004
rect 291339 88964 291384 88992
rect 291378 88952 291384 88964
rect 291436 88952 291442 89004
rect 389358 87904 389364 87916
rect 389319 87876 389364 87904
rect 389358 87864 389364 87876
rect 389416 87864 389422 87916
rect 395890 87184 395896 87236
rect 395948 87184 395954 87236
rect 395982 87184 395988 87236
rect 396040 87184 396046 87236
rect 251174 87048 251180 87100
rect 251232 87088 251238 87100
rect 260650 87088 260656 87100
rect 251232 87060 260656 87088
rect 251232 87048 251238 87060
rect 260650 87048 260656 87060
rect 260708 87048 260714 87100
rect 297542 87048 297548 87100
rect 297600 87088 297606 87100
rect 306282 87088 306288 87100
rect 297600 87060 306288 87088
rect 297600 87048 297606 87060
rect 306282 87048 306288 87060
rect 306340 87048 306346 87100
rect 376754 87048 376760 87100
rect 376812 87088 376818 87100
rect 386230 87088 386236 87100
rect 376812 87060 386236 87088
rect 376812 87048 376818 87060
rect 386230 87048 386236 87060
rect 386288 87048 386294 87100
rect 386414 87048 386420 87100
rect 386472 87088 386478 87100
rect 395798 87088 395804 87100
rect 386472 87060 395804 87088
rect 386472 87048 386478 87060
rect 395798 87048 395804 87060
rect 395856 87048 395862 87100
rect 395908 87032 395936 87184
rect 396000 87032 396028 87184
rect 437198 87116 437204 87168
rect 437256 87156 437262 87168
rect 437474 87156 437480 87168
rect 437256 87128 437480 87156
rect 437256 87116 437262 87128
rect 437474 87116 437480 87128
rect 437532 87116 437538 87168
rect 456518 87116 456524 87168
rect 456576 87156 456582 87168
rect 456978 87156 456984 87168
rect 456576 87128 456984 87156
rect 456576 87116 456582 87128
rect 456978 87116 456984 87128
rect 457036 87116 457042 87168
rect 494606 87116 494612 87168
rect 494664 87156 494670 87168
rect 502242 87156 502248 87168
rect 494664 87128 502248 87156
rect 494664 87116 494670 87128
rect 502242 87116 502248 87128
rect 502300 87116 502306 87168
rect 262582 86980 262588 87032
rect 262640 87020 262646 87032
rect 262674 87020 262680 87032
rect 262640 86992 262680 87020
rect 262640 86980 262646 86992
rect 262674 86980 262680 86992
rect 262732 86980 262738 87032
rect 294414 86980 294420 87032
rect 294472 86980 294478 87032
rect 347774 86980 347780 87032
rect 347832 87020 347838 87032
rect 357342 87020 357348 87032
rect 347832 86992 357348 87020
rect 347832 86980 347838 86992
rect 357342 86980 357348 86992
rect 357400 86980 357406 87032
rect 367002 87020 367008 87032
rect 366963 86992 367008 87020
rect 367002 86980 367008 86992
rect 367060 86980 367066 87032
rect 395890 86980 395896 87032
rect 395948 86980 395954 87032
rect 395982 86980 395988 87032
rect 396040 86980 396046 87032
rect 421190 87020 421196 87032
rect 421151 86992 421196 87020
rect 421190 86980 421196 86992
rect 421248 86980 421254 87032
rect 251450 86952 251456 86964
rect 251411 86924 251456 86952
rect 251450 86912 251456 86924
rect 251508 86912 251514 86964
rect 294432 86896 294460 86980
rect 324590 86912 324596 86964
rect 324648 86912 324654 86964
rect 327166 86912 327172 86964
rect 327224 86952 327230 86964
rect 327258 86952 327264 86964
rect 327224 86924 327264 86952
rect 327224 86912 327230 86924
rect 327258 86912 327264 86924
rect 327316 86912 327322 86964
rect 336918 86912 336924 86964
rect 336976 86912 336982 86964
rect 341061 86955 341119 86961
rect 341061 86921 341073 86955
rect 341107 86952 341119 86955
rect 341150 86952 341156 86964
rect 341107 86924 341156 86952
rect 341107 86921 341119 86924
rect 341061 86915 341119 86921
rect 341150 86912 341156 86924
rect 341208 86912 341214 86964
rect 294414 86844 294420 86896
rect 294472 86844 294478 86896
rect 324608 86884 324636 86912
rect 324682 86884 324688 86896
rect 324608 86856 324688 86884
rect 324682 86844 324688 86856
rect 324740 86844 324746 86896
rect 336936 86828 336964 86912
rect 336918 86776 336924 86828
rect 336976 86776 336982 86828
rect 265250 85552 265256 85604
rect 265308 85592 265314 85604
rect 265342 85592 265348 85604
rect 265308 85564 265348 85592
rect 265308 85552 265314 85564
rect 265342 85552 265348 85564
rect 265400 85552 265406 85604
rect 266633 85595 266691 85601
rect 266633 85561 266645 85595
rect 266679 85592 266691 85595
rect 266722 85592 266728 85604
rect 266679 85564 266728 85592
rect 266679 85561 266691 85564
rect 266633 85555 266691 85561
rect 266722 85552 266728 85564
rect 266780 85552 266786 85604
rect 267734 85552 267740 85604
rect 267792 85592 267798 85604
rect 267826 85592 267832 85604
rect 267792 85564 267832 85592
rect 267792 85552 267798 85564
rect 267826 85552 267832 85564
rect 267884 85552 267890 85604
rect 272150 85552 272156 85604
rect 272208 85592 272214 85604
rect 272334 85592 272340 85604
rect 272208 85564 272340 85592
rect 272208 85552 272214 85564
rect 272334 85552 272340 85564
rect 272392 85552 272398 85604
rect 299842 85552 299848 85604
rect 299900 85592 299906 85604
rect 299934 85592 299940 85604
rect 299900 85564 299940 85592
rect 299900 85552 299906 85564
rect 299934 85552 299940 85564
rect 299992 85552 299998 85604
rect 301130 85552 301136 85604
rect 301188 85592 301194 85604
rect 301222 85592 301228 85604
rect 301188 85564 301228 85592
rect 301188 85552 301194 85564
rect 301222 85552 301228 85564
rect 301280 85552 301286 85604
rect 306742 85552 306748 85604
rect 306800 85592 306806 85604
rect 306834 85592 306840 85604
rect 306800 85564 306840 85592
rect 306800 85552 306806 85564
rect 306834 85552 306840 85564
rect 306892 85552 306898 85604
rect 310790 85592 310796 85604
rect 310751 85564 310796 85592
rect 310790 85552 310796 85564
rect 310848 85552 310854 85604
rect 323026 85552 323032 85604
rect 323084 85592 323090 85604
rect 323394 85592 323400 85604
rect 323084 85564 323400 85592
rect 323084 85552 323090 85564
rect 323394 85552 323400 85564
rect 323452 85552 323458 85604
rect 325878 85552 325884 85604
rect 325936 85592 325942 85604
rect 325970 85592 325976 85604
rect 325936 85564 325976 85592
rect 325936 85552 325942 85564
rect 325970 85552 325976 85564
rect 326028 85552 326034 85604
rect 339494 85552 339500 85604
rect 339552 85592 339558 85604
rect 339862 85592 339868 85604
rect 339552 85564 339868 85592
rect 339552 85552 339558 85564
rect 339862 85552 339868 85564
rect 339920 85552 339926 85604
rect 362313 85595 362371 85601
rect 362313 85561 362325 85595
rect 362359 85592 362371 85595
rect 362402 85592 362408 85604
rect 362359 85564 362408 85592
rect 362359 85561 362371 85564
rect 362313 85555 362371 85561
rect 362402 85552 362408 85564
rect 362460 85552 362466 85604
rect 232225 85527 232283 85533
rect 232225 85493 232237 85527
rect 232271 85524 232283 85527
rect 232314 85524 232320 85536
rect 232271 85496 232320 85524
rect 232271 85493 232283 85496
rect 232225 85487 232283 85493
rect 232314 85484 232320 85496
rect 232372 85484 232378 85536
rect 317693 85527 317751 85533
rect 317693 85493 317705 85527
rect 317739 85524 317751 85527
rect 317874 85524 317880 85536
rect 317739 85496 317880 85524
rect 317739 85493 317751 85496
rect 317693 85487 317751 85493
rect 317874 85484 317880 85496
rect 317932 85484 317938 85536
rect 360197 85527 360255 85533
rect 360197 85493 360209 85527
rect 360243 85524 360255 85527
rect 360378 85524 360384 85536
rect 360243 85496 360384 85524
rect 360243 85493 360255 85496
rect 360197 85487 360255 85493
rect 360378 85484 360384 85496
rect 360436 85484 360442 85536
rect 421009 85527 421067 85533
rect 421009 85493 421021 85527
rect 421055 85524 421067 85527
rect 421190 85524 421196 85536
rect 421055 85496 421196 85524
rect 421055 85493 421067 85496
rect 421009 85487 421067 85493
rect 421190 85484 421196 85496
rect 421248 85484 421254 85536
rect 266722 84164 266728 84176
rect 266683 84136 266728 84164
rect 266722 84124 266728 84136
rect 266780 84124 266786 84176
rect 267737 84167 267795 84173
rect 267737 84133 267749 84167
rect 267783 84164 267795 84167
rect 267826 84164 267832 84176
rect 267783 84136 267832 84164
rect 267783 84133 267795 84136
rect 267737 84127 267795 84133
rect 267826 84124 267832 84136
rect 267884 84124 267890 84176
rect 284665 84167 284723 84173
rect 284665 84133 284677 84167
rect 284711 84164 284723 84167
rect 284754 84164 284760 84176
rect 284711 84136 284760 84164
rect 284711 84133 284723 84136
rect 284665 84127 284723 84133
rect 284754 84124 284760 84136
rect 284812 84124 284818 84176
rect 285953 84167 286011 84173
rect 285953 84133 285965 84167
rect 285999 84164 286011 84167
rect 286042 84164 286048 84176
rect 285999 84136 286048 84164
rect 285999 84133 286011 84136
rect 285953 84127 286011 84133
rect 286042 84124 286048 84136
rect 286100 84124 286106 84176
rect 288710 84164 288716 84176
rect 288671 84136 288716 84164
rect 288710 84124 288716 84136
rect 288768 84124 288774 84176
rect 289906 84164 289912 84176
rect 289867 84136 289912 84164
rect 289906 84124 289912 84136
rect 289964 84124 289970 84176
rect 296990 84164 296996 84176
rect 296951 84136 296996 84164
rect 296990 84124 296996 84136
rect 297048 84124 297054 84176
rect 306745 84167 306803 84173
rect 306745 84133 306757 84167
rect 306791 84164 306803 84167
rect 306834 84164 306840 84176
rect 306791 84136 306840 84164
rect 306791 84133 306803 84136
rect 306745 84127 306803 84133
rect 306834 84124 306840 84136
rect 306892 84124 306898 84176
rect 330113 82943 330171 82949
rect 330113 82909 330125 82943
rect 330159 82940 330171 82943
rect 330294 82940 330300 82952
rect 330159 82912 330300 82940
rect 330159 82909 330171 82912
rect 330113 82903 330171 82909
rect 330294 82900 330300 82912
rect 330352 82900 330358 82952
rect 357710 80152 357716 80164
rect 357636 80124 357716 80152
rect 357636 80096 357664 80124
rect 357710 80112 357716 80124
rect 357768 80112 357774 80164
rect 372890 80152 372896 80164
rect 372724 80124 372896 80152
rect 303890 80044 303896 80096
rect 303948 80044 303954 80096
rect 357618 80044 357624 80096
rect 357676 80044 357682 80096
rect 303908 79960 303936 80044
rect 372724 80028 372752 80124
rect 372890 80112 372896 80124
rect 372948 80112 372954 80164
rect 389358 80044 389364 80096
rect 389416 80044 389422 80096
rect 463786 80044 463792 80096
rect 463844 80044 463850 80096
rect 372706 79976 372712 80028
rect 372764 79976 372770 80028
rect 375834 79976 375840 80028
rect 375892 79976 375898 80028
rect 377122 79976 377128 80028
rect 377180 79976 377186 80028
rect 303890 79908 303896 79960
rect 303948 79908 303954 79960
rect 375852 79948 375880 79976
rect 375926 79948 375932 79960
rect 375852 79920 375932 79948
rect 375926 79908 375932 79920
rect 375984 79908 375990 79960
rect 377140 79948 377168 79976
rect 377214 79948 377220 79960
rect 377140 79920 377220 79948
rect 377214 79908 377220 79920
rect 377272 79908 377278 79960
rect 389376 79948 389404 80044
rect 463804 79960 463832 80044
rect 389450 79948 389456 79960
rect 389376 79920 389456 79948
rect 389450 79908 389456 79920
rect 389508 79908 389514 79960
rect 463786 79908 463792 79960
rect 463844 79908 463850 79960
rect 2774 79772 2780 79824
rect 2832 79812 2838 79824
rect 4890 79812 4896 79824
rect 2832 79784 4896 79812
rect 2832 79772 2838 79784
rect 4890 79772 4896 79784
rect 4948 79772 4954 79824
rect 250070 77392 250076 77444
rect 250128 77392 250134 77444
rect 236270 77256 236276 77308
rect 236328 77296 236334 77308
rect 236454 77296 236460 77308
rect 236328 77268 236460 77296
rect 236328 77256 236334 77268
rect 236454 77256 236460 77268
rect 236512 77256 236518 77308
rect 249978 77256 249984 77308
rect 250036 77296 250042 77308
rect 250088 77296 250116 77392
rect 301222 77364 301228 77376
rect 301183 77336 301228 77364
rect 301222 77324 301228 77336
rect 301280 77324 301286 77376
rect 251450 77296 251456 77308
rect 250036 77268 250116 77296
rect 251411 77268 251456 77296
rect 250036 77256 250042 77268
rect 251450 77256 251456 77268
rect 251508 77256 251514 77308
rect 262582 77256 262588 77308
rect 262640 77296 262646 77308
rect 262674 77296 262680 77308
rect 262640 77268 262680 77296
rect 262640 77256 262646 77268
rect 262674 77256 262680 77268
rect 262732 77256 262738 77308
rect 299750 77256 299756 77308
rect 299808 77296 299814 77308
rect 299842 77296 299848 77308
rect 299808 77268 299848 77296
rect 299808 77256 299814 77268
rect 299842 77256 299848 77268
rect 299900 77256 299906 77308
rect 302510 77256 302516 77308
rect 302568 77296 302574 77308
rect 302602 77296 302608 77308
rect 302568 77268 302608 77296
rect 302568 77256 302574 77268
rect 302602 77256 302608 77268
rect 302660 77256 302666 77308
rect 341058 77296 341064 77308
rect 341019 77268 341064 77296
rect 341058 77256 341064 77268
rect 341116 77256 341122 77308
rect 303890 77188 303896 77240
rect 303948 77228 303954 77240
rect 303982 77228 303988 77240
rect 303948 77200 303988 77228
rect 303948 77188 303954 77200
rect 303982 77188 303988 77200
rect 304040 77188 304046 77240
rect 389361 77231 389419 77237
rect 389361 77197 389373 77231
rect 389407 77228 389419 77231
rect 389450 77228 389456 77240
rect 389407 77200 389456 77228
rect 389407 77197 389419 77200
rect 389361 77191 389419 77197
rect 389450 77188 389456 77200
rect 389508 77188 389514 77240
rect 341058 77160 341064 77172
rect 341019 77132 341064 77160
rect 341058 77120 341064 77132
rect 341116 77120 341122 77172
rect 294230 76440 294236 76492
rect 294288 76480 294294 76492
rect 294414 76480 294420 76492
rect 294288 76452 294420 76480
rect 294288 76440 294294 76452
rect 294414 76440 294420 76452
rect 294472 76440 294478 76492
rect 367094 76168 367100 76220
rect 367152 76208 367158 76220
rect 376662 76208 376668 76220
rect 367152 76180 376668 76208
rect 367152 76168 367158 76180
rect 376662 76168 376668 76180
rect 376720 76168 376726 76220
rect 396074 76032 396080 76084
rect 396132 76072 396138 76084
rect 399386 76072 399392 76084
rect 396132 76044 399392 76072
rect 396132 76032 396138 76044
rect 399386 76032 399392 76044
rect 399444 76032 399450 76084
rect 437198 76032 437204 76084
rect 437256 76072 437262 76084
rect 437474 76072 437480 76084
rect 437256 76044 437480 76072
rect 437256 76032 437262 76044
rect 437474 76032 437480 76044
rect 437532 76032 437538 76084
rect 456518 76032 456524 76084
rect 456576 76072 456582 76084
rect 456794 76072 456800 76084
rect 456576 76044 456800 76072
rect 456576 76032 456582 76044
rect 456794 76032 456800 76044
rect 456852 76032 456858 76084
rect 232222 75936 232228 75948
rect 232183 75908 232228 75936
rect 232222 75896 232228 75908
rect 232280 75896 232286 75948
rect 270494 75896 270500 75948
rect 270552 75936 270558 75948
rect 270678 75936 270684 75948
rect 270552 75908 270684 75936
rect 270552 75896 270558 75908
rect 270678 75896 270684 75908
rect 270736 75896 270742 75948
rect 306374 75896 306380 75948
rect 306432 75936 306438 75948
rect 311250 75936 311256 75948
rect 306432 75908 311256 75936
rect 306432 75896 306438 75908
rect 311250 75896 311256 75908
rect 311308 75896 311314 75948
rect 317690 75936 317696 75948
rect 317651 75908 317696 75936
rect 317690 75896 317696 75908
rect 317748 75896 317754 75948
rect 323026 75896 323032 75948
rect 323084 75936 323090 75948
rect 323302 75936 323308 75948
rect 323084 75908 323308 75936
rect 323084 75896 323090 75908
rect 323302 75896 323308 75908
rect 323360 75896 323366 75948
rect 358722 75896 358728 75948
rect 358780 75936 358786 75948
rect 358998 75936 359004 75948
rect 358780 75908 359004 75936
rect 358780 75896 358786 75908
rect 358998 75896 359004 75908
rect 359056 75896 359062 75948
rect 360194 75936 360200 75948
rect 360155 75908 360200 75936
rect 360194 75896 360200 75908
rect 360252 75896 360258 75948
rect 362218 75896 362224 75948
rect 362276 75936 362282 75948
rect 362402 75936 362408 75948
rect 362276 75908 362408 75936
rect 362276 75896 362282 75908
rect 362402 75896 362408 75908
rect 362460 75896 362466 75948
rect 421006 75936 421012 75948
rect 420967 75908 421012 75936
rect 421006 75896 421012 75908
rect 421064 75896 421070 75948
rect 301222 75868 301228 75880
rect 301183 75840 301228 75868
rect 301222 75828 301228 75840
rect 301280 75828 301286 75880
rect 310790 75868 310796 75880
rect 310751 75840 310796 75868
rect 310790 75828 310796 75840
rect 310848 75828 310854 75880
rect 330202 75868 330208 75880
rect 330163 75840 330208 75868
rect 330202 75828 330208 75840
rect 330260 75828 330266 75880
rect 288713 75803 288771 75809
rect 288713 75769 288725 75803
rect 288759 75800 288771 75803
rect 288894 75800 288900 75812
rect 288759 75772 288900 75800
rect 288759 75769 288771 75772
rect 288713 75763 288771 75769
rect 288894 75760 288900 75772
rect 288952 75760 288958 75812
rect 306742 75800 306748 75812
rect 306703 75772 306748 75800
rect 306742 75760 306748 75772
rect 306800 75760 306806 75812
rect 266725 74579 266783 74585
rect 266725 74545 266737 74579
rect 266771 74576 266783 74579
rect 266814 74576 266820 74588
rect 266771 74548 266820 74576
rect 266771 74545 266783 74548
rect 266725 74539 266783 74545
rect 266814 74536 266820 74548
rect 266872 74536 266878 74588
rect 267734 74536 267740 74588
rect 267792 74576 267798 74588
rect 289909 74579 289967 74585
rect 267792 74548 267837 74576
rect 267792 74536 267798 74548
rect 289909 74545 289921 74579
rect 289955 74576 289967 74579
rect 289998 74576 290004 74588
rect 289955 74548 290004 74576
rect 289955 74545 289967 74548
rect 289909 74539 289967 74545
rect 289998 74536 290004 74548
rect 290056 74536 290062 74588
rect 296898 74536 296904 74588
rect 296956 74576 296962 74588
rect 296993 74579 297051 74585
rect 296993 74576 297005 74579
rect 296956 74548 297005 74576
rect 296956 74536 296962 74548
rect 296993 74545 297005 74548
rect 297039 74545 297051 74579
rect 296993 74539 297051 74545
rect 359090 74536 359096 74588
rect 359148 74576 359154 74588
rect 359182 74576 359188 74588
rect 359148 74548 359188 74576
rect 359148 74536 359154 74548
rect 359182 74536 359188 74548
rect 359240 74536 359246 74588
rect 362218 74468 362224 74520
rect 362276 74508 362282 74520
rect 362402 74508 362408 74520
rect 362276 74480 362408 74508
rect 362276 74468 362282 74480
rect 362402 74468 362408 74480
rect 362460 74468 362466 74520
rect 296809 74443 296867 74449
rect 296809 74409 296821 74443
rect 296855 74440 296867 74443
rect 296898 74440 296904 74452
rect 296855 74412 296904 74440
rect 296855 74409 296867 74412
rect 296809 74403 296867 74409
rect 296898 74400 296904 74412
rect 296956 74400 296962 74452
rect 272153 72471 272211 72477
rect 272153 72437 272165 72471
rect 272199 72468 272211 72471
rect 272242 72468 272248 72480
rect 272199 72440 272248 72468
rect 272199 72437 272211 72440
rect 272153 72431 272211 72437
rect 272242 72428 272248 72440
rect 272300 72428 272306 72480
rect 357618 70496 357624 70508
rect 357579 70468 357624 70496
rect 357618 70456 357624 70468
rect 357676 70456 357682 70508
rect 341061 70295 341119 70301
rect 341061 70261 341073 70295
rect 341107 70292 341119 70295
rect 341150 70292 341156 70304
rect 341107 70264 341156 70292
rect 341107 70261 341119 70264
rect 341061 70255 341119 70261
rect 341150 70252 341156 70264
rect 341208 70252 341214 70304
rect 330202 69952 330208 69964
rect 330163 69924 330208 69952
rect 330202 69912 330208 69924
rect 330260 69912 330266 69964
rect 302510 67708 302516 67720
rect 302436 67680 302516 67708
rect 302436 67652 302464 67680
rect 302510 67668 302516 67680
rect 302568 67668 302574 67720
rect 272150 67640 272156 67652
rect 272111 67612 272156 67640
rect 272150 67600 272156 67612
rect 272208 67600 272214 67652
rect 302418 67600 302424 67652
rect 302476 67600 302482 67652
rect 325878 67600 325884 67652
rect 325936 67640 325942 67652
rect 325970 67640 325976 67652
rect 325936 67612 325976 67640
rect 325936 67600 325942 67612
rect 325970 67600 325976 67612
rect 326028 67600 326034 67652
rect 389358 67640 389364 67652
rect 389319 67612 389364 67640
rect 389358 67600 389364 67612
rect 389416 67600 389422 67652
rect 236270 67572 236276 67584
rect 236231 67544 236276 67572
rect 236270 67532 236276 67544
rect 236328 67532 236334 67584
rect 273622 67572 273628 67584
rect 273583 67544 273628 67572
rect 273622 67532 273628 67544
rect 273680 67532 273686 67584
rect 270678 66308 270684 66360
rect 270736 66348 270742 66360
rect 310790 66348 310796 66360
rect 270736 66320 270816 66348
rect 310751 66320 310796 66348
rect 270736 66308 270742 66320
rect 270788 66292 270816 66320
rect 310790 66308 310796 66320
rect 310848 66308 310854 66360
rect 266630 66240 266636 66292
rect 266688 66280 266694 66292
rect 266814 66280 266820 66292
rect 266688 66252 266820 66280
rect 266688 66240 266694 66252
rect 266814 66240 266820 66252
rect 266872 66240 266878 66292
rect 270770 66240 270776 66292
rect 270828 66240 270834 66292
rect 284662 66280 284668 66292
rect 284623 66252 284668 66280
rect 284662 66240 284668 66252
rect 284720 66240 284726 66292
rect 285950 66280 285956 66292
rect 285911 66252 285956 66280
rect 285950 66240 285956 66252
rect 286008 66240 286014 66292
rect 301038 66240 301044 66292
rect 301096 66280 301102 66292
rect 301222 66280 301228 66292
rect 301096 66252 301228 66280
rect 301096 66240 301102 66252
rect 301222 66240 301228 66252
rect 301280 66240 301286 66292
rect 306650 66240 306656 66292
rect 306708 66280 306714 66292
rect 306742 66280 306748 66292
rect 306708 66252 306748 66280
rect 306708 66240 306714 66252
rect 306742 66240 306748 66252
rect 306800 66240 306806 66292
rect 357618 66280 357624 66292
rect 357579 66252 357624 66280
rect 357618 66240 357624 66252
rect 357676 66240 357682 66292
rect 232225 66215 232283 66221
rect 232225 66181 232237 66215
rect 232271 66212 232283 66215
rect 232314 66212 232320 66224
rect 232271 66184 232320 66212
rect 232271 66181 232283 66184
rect 232225 66175 232283 66181
rect 232314 66172 232320 66184
rect 232372 66172 232378 66224
rect 250070 66212 250076 66224
rect 250031 66184 250076 66212
rect 250070 66172 250076 66184
rect 250128 66172 250134 66224
rect 265158 66172 265164 66224
rect 265216 66212 265222 66224
rect 265253 66215 265311 66221
rect 265253 66212 265265 66215
rect 265216 66184 265265 66212
rect 265216 66172 265222 66184
rect 265253 66181 265265 66184
rect 265299 66181 265311 66215
rect 310790 66212 310796 66224
rect 310751 66184 310796 66212
rect 265253 66175 265311 66181
rect 310790 66172 310796 66184
rect 310848 66172 310854 66224
rect 325878 66172 325884 66224
rect 325936 66212 325942 66224
rect 325973 66215 326031 66221
rect 325973 66212 325985 66215
rect 325936 66184 325985 66212
rect 325936 66172 325942 66184
rect 325973 66181 325985 66184
rect 326019 66181 326031 66215
rect 327166 66212 327172 66224
rect 327127 66184 327172 66212
rect 325973 66175 326031 66181
rect 327166 66172 327172 66184
rect 327224 66172 327230 66224
rect 336918 66212 336924 66224
rect 336879 66184 336924 66212
rect 336918 66172 336924 66184
rect 336976 66172 336982 66224
rect 421101 66215 421159 66221
rect 421101 66181 421113 66215
rect 421147 66212 421159 66215
rect 421190 66212 421196 66224
rect 421147 66184 421196 66212
rect 421147 66181 421159 66184
rect 421101 66175 421159 66181
rect 421190 66172 421196 66184
rect 421248 66172 421254 66224
rect 296806 64920 296812 64932
rect 296767 64892 296812 64920
rect 296806 64880 296812 64892
rect 296864 64880 296870 64932
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 24118 64852 24124 64864
rect 3384 64824 24124 64852
rect 3384 64812 3390 64824
rect 24118 64812 24124 64824
rect 24176 64812 24182 64864
rect 267734 64812 267740 64864
rect 267792 64852 267798 64864
rect 294230 64852 294236 64864
rect 267792 64824 267837 64852
rect 294191 64824 294236 64852
rect 267792 64812 267798 64824
rect 294230 64812 294236 64824
rect 294288 64812 294294 64864
rect 324866 64812 324872 64864
rect 324924 64852 324930 64864
rect 324958 64852 324964 64864
rect 324924 64824 324964 64852
rect 324924 64812 324930 64824
rect 324958 64812 324964 64824
rect 325016 64812 325022 64864
rect 359090 64852 359096 64864
rect 359051 64824 359096 64852
rect 359090 64812 359096 64824
rect 359148 64812 359154 64864
rect 362221 64855 362279 64861
rect 362221 64821 362233 64855
rect 362267 64852 362279 64855
rect 362494 64852 362500 64864
rect 362267 64824 362500 64852
rect 362267 64821 362279 64824
rect 362221 64815 362279 64821
rect 362494 64812 362500 64824
rect 362552 64812 362558 64864
rect 414014 63724 414020 63776
rect 414072 63764 414078 63776
rect 418890 63764 418896 63776
rect 414072 63736 418896 63764
rect 414072 63724 414078 63736
rect 418890 63724 418896 63736
rect 418948 63724 418954 63776
rect 437198 63656 437204 63708
rect 437256 63696 437262 63708
rect 437474 63696 437480 63708
rect 437256 63668 437480 63696
rect 437256 63656 437262 63668
rect 437474 63656 437480 63668
rect 437532 63656 437538 63708
rect 456518 63656 456524 63708
rect 456576 63696 456582 63708
rect 456886 63696 456892 63708
rect 456576 63668 456892 63696
rect 456576 63656 456582 63668
rect 456886 63656 456892 63668
rect 456944 63656 456950 63708
rect 266630 61452 266636 61464
rect 266591 61424 266636 61452
rect 266630 61412 266636 61424
rect 266688 61412 266694 61464
rect 323302 61452 323308 61464
rect 323263 61424 323308 61452
rect 323302 61412 323308 61424
rect 323360 61412 323366 61464
rect 250070 60704 250076 60716
rect 250031 60676 250076 60704
rect 250070 60664 250076 60676
rect 250128 60664 250134 60716
rect 259638 60664 259644 60716
rect 259696 60704 259702 60716
rect 259822 60704 259828 60716
rect 259696 60676 259828 60704
rect 259696 60664 259702 60676
rect 259822 60664 259828 60676
rect 259880 60664 259886 60716
rect 262582 60664 262588 60716
rect 262640 60704 262646 60716
rect 262766 60704 262772 60716
rect 262640 60676 262772 60704
rect 262640 60664 262646 60676
rect 262766 60664 262772 60676
rect 262824 60664 262830 60716
rect 339678 60664 339684 60716
rect 339736 60704 339742 60716
rect 339862 60704 339868 60716
rect 339736 60676 339868 60704
rect 339736 60664 339742 60676
rect 339862 60664 339868 60676
rect 339920 60664 339926 60716
rect 341150 60664 341156 60716
rect 341208 60704 341214 60716
rect 341334 60704 341340 60716
rect 341208 60676 341340 60704
rect 341208 60664 341214 60676
rect 341334 60664 341340 60676
rect 341392 60664 341398 60716
rect 360286 60664 360292 60716
rect 360344 60704 360350 60716
rect 360470 60704 360476 60716
rect 360344 60676 360476 60704
rect 360344 60664 360350 60676
rect 360470 60664 360476 60676
rect 360528 60664 360534 60716
rect 306650 59984 306656 60036
rect 306708 60024 306714 60036
rect 306745 60027 306803 60033
rect 306745 60024 306757 60027
rect 306708 59996 306757 60024
rect 306708 59984 306714 59996
rect 306745 59993 306757 59996
rect 306791 59993 306803 60027
rect 306745 59987 306803 59993
rect 310793 60027 310851 60033
rect 310793 59993 310805 60027
rect 310839 60024 310851 60027
rect 311066 60024 311072 60036
rect 310839 59996 311072 60024
rect 310839 59993 310851 59996
rect 310793 59987 310851 59993
rect 311066 59984 311072 59996
rect 311124 59984 311130 60036
rect 272150 58012 272156 58064
rect 272208 58012 272214 58064
rect 236270 57984 236276 57996
rect 236231 57956 236276 57984
rect 236270 57944 236276 57956
rect 236328 57944 236334 57996
rect 272168 57928 272196 58012
rect 273622 57984 273628 57996
rect 273583 57956 273628 57984
rect 273622 57944 273628 57956
rect 273680 57944 273686 57996
rect 299750 57944 299756 57996
rect 299808 57984 299814 57996
rect 299842 57984 299848 57996
rect 299808 57956 299848 57984
rect 299808 57944 299814 57956
rect 299842 57944 299848 57956
rect 299900 57944 299906 57996
rect 302418 57944 302424 57996
rect 302476 57984 302482 57996
rect 302510 57984 302516 57996
rect 302476 57956 302516 57984
rect 302476 57944 302482 57956
rect 302510 57944 302516 57956
rect 302568 57944 302574 57996
rect 303890 57944 303896 57996
rect 303948 57984 303954 57996
rect 303982 57984 303988 57996
rect 303948 57956 303988 57984
rect 303948 57944 303954 57956
rect 303982 57944 303988 57956
rect 304040 57944 304046 57996
rect 245562 57876 245568 57928
rect 245620 57916 245626 57928
rect 245930 57916 245936 57928
rect 245620 57888 245936 57916
rect 245620 57876 245626 57888
rect 245930 57876 245936 57888
rect 245988 57876 245994 57928
rect 272150 57876 272156 57928
rect 272208 57876 272214 57928
rect 289998 57876 290004 57928
rect 290056 57916 290062 57928
rect 290090 57916 290096 57928
rect 290056 57888 290096 57916
rect 290056 57876 290062 57888
rect 290090 57876 290096 57888
rect 290148 57876 290154 57928
rect 291470 57876 291476 57928
rect 291528 57916 291534 57928
rect 291562 57916 291568 57928
rect 291528 57888 291568 57916
rect 291528 57876 291534 57888
rect 291562 57876 291568 57888
rect 291620 57876 291626 57928
rect 301038 57916 301044 57928
rect 300999 57888 301044 57916
rect 301038 57876 301044 57888
rect 301096 57876 301102 57928
rect 339773 57919 339831 57925
rect 339773 57885 339785 57919
rect 339819 57916 339831 57919
rect 339862 57916 339868 57928
rect 339819 57888 339868 57916
rect 339819 57885 339831 57888
rect 339773 57879 339831 57885
rect 339862 57876 339868 57888
rect 339920 57876 339926 57928
rect 367002 57916 367008 57928
rect 366963 57888 367008 57916
rect 367002 57876 367008 57888
rect 367060 57876 367066 57928
rect 389174 57916 389180 57928
rect 389135 57888 389180 57916
rect 389174 57876 389180 57888
rect 389232 57876 389238 57928
rect 470594 57916 470600 57928
rect 470555 57888 470600 57916
rect 470594 57876 470600 57888
rect 470652 57876 470658 57928
rect 284662 57032 284668 57044
rect 284623 57004 284668 57032
rect 284662 56992 284668 57004
rect 284720 56992 284726 57044
rect 421098 56692 421104 56704
rect 421059 56664 421104 56692
rect 421098 56652 421104 56664
rect 421156 56652 421162 56704
rect 327169 56627 327227 56633
rect 327169 56593 327181 56627
rect 327215 56624 327227 56627
rect 327258 56624 327264 56636
rect 327215 56596 327264 56624
rect 327215 56593 327227 56596
rect 327169 56587 327227 56593
rect 327258 56584 327264 56596
rect 327316 56584 327322 56636
rect 336918 56624 336924 56636
rect 336879 56596 336924 56624
rect 336918 56584 336924 56596
rect 336976 56584 336982 56636
rect 286042 56516 286048 56568
rect 286100 56556 286106 56568
rect 337286 56556 337292 56568
rect 286100 56528 286145 56556
rect 337247 56528 337292 56556
rect 286100 56516 286106 56528
rect 337286 56516 337292 56528
rect 337344 56516 337350 56568
rect 359090 56556 359096 56568
rect 359051 56528 359096 56556
rect 359090 56516 359096 56528
rect 359148 56516 359154 56568
rect 421009 56559 421067 56565
rect 421009 56525 421021 56559
rect 421055 56556 421067 56559
rect 421098 56556 421104 56568
rect 421055 56528 421104 56556
rect 421055 56525 421067 56528
rect 421009 56519 421067 56525
rect 421098 56516 421104 56528
rect 421156 56516 421162 56568
rect 267737 55267 267795 55273
rect 267737 55233 267749 55267
rect 267783 55264 267795 55267
rect 268102 55264 268108 55276
rect 267783 55236 268108 55264
rect 267783 55233 267795 55236
rect 267737 55227 267795 55233
rect 268102 55224 268108 55236
rect 268160 55224 268166 55276
rect 294230 55264 294236 55276
rect 294191 55236 294236 55264
rect 294230 55224 294236 55236
rect 294288 55224 294294 55276
rect 317506 55224 317512 55276
rect 317564 55264 317570 55276
rect 317690 55264 317696 55276
rect 317564 55236 317696 55264
rect 317564 55224 317570 55236
rect 317690 55224 317696 55236
rect 317748 55224 317754 55276
rect 362218 55264 362224 55276
rect 362179 55236 362224 55264
rect 362218 55224 362224 55236
rect 362276 55224 362282 55276
rect 424502 53836 424508 53848
rect 424463 53808 424508 53836
rect 424502 53796 424508 53808
rect 424560 53796 424566 53848
rect 262582 52232 262588 52284
rect 262640 52272 262646 52284
rect 262766 52272 262772 52284
rect 262640 52244 262772 52272
rect 262640 52232 262646 52244
rect 262766 52232 262772 52244
rect 262824 52232 262830 52284
rect 306745 52003 306803 52009
rect 306745 51969 306757 52003
rect 306791 52000 306803 52003
rect 307018 52000 307024 52012
rect 306791 51972 307024 52000
rect 306791 51969 306803 51972
rect 306745 51963 306803 51969
rect 307018 51960 307024 51972
rect 307076 51960 307082 52012
rect 301038 51796 301044 51808
rect 300999 51768 301044 51796
rect 301038 51756 301044 51768
rect 301096 51756 301102 51808
rect 244458 51116 244464 51128
rect 244384 51088 244464 51116
rect 244384 51060 244412 51088
rect 244458 51076 244464 51088
rect 244516 51076 244522 51128
rect 244366 51008 244372 51060
rect 244424 51008 244430 51060
rect 250070 50980 250076 50992
rect 250031 50952 250076 50980
rect 250070 50940 250076 50952
rect 250128 50940 250134 50992
rect 2774 50464 2780 50516
rect 2832 50504 2838 50516
rect 4798 50504 4804 50516
rect 2832 50476 4804 50504
rect 2832 50464 2838 50476
rect 4798 50464 4804 50476
rect 4856 50464 4862 50516
rect 232222 48328 232228 48340
rect 232183 48300 232228 48328
rect 232222 48288 232228 48300
rect 232280 48288 232286 48340
rect 250070 48328 250076 48340
rect 250031 48300 250076 48328
rect 250070 48288 250076 48300
rect 250128 48288 250134 48340
rect 266630 48328 266636 48340
rect 266591 48300 266636 48328
rect 266630 48288 266636 48300
rect 266688 48288 266694 48340
rect 284665 48331 284723 48337
rect 284665 48297 284677 48331
rect 284711 48328 284723 48331
rect 284754 48328 284760 48340
rect 284711 48300 284760 48328
rect 284711 48297 284723 48300
rect 284665 48291 284723 48297
rect 284754 48288 284760 48300
rect 284812 48288 284818 48340
rect 323302 48328 323308 48340
rect 323263 48300 323308 48328
rect 323302 48288 323308 48300
rect 323360 48288 323366 48340
rect 339770 48328 339776 48340
rect 339731 48300 339776 48328
rect 339770 48288 339776 48300
rect 339828 48288 339834 48340
rect 358630 48288 358636 48340
rect 358688 48328 358694 48340
rect 358722 48328 358728 48340
rect 358688 48300 358728 48328
rect 358688 48288 358694 48300
rect 358722 48288 358728 48300
rect 358780 48288 358786 48340
rect 367002 48328 367008 48340
rect 366963 48300 367008 48328
rect 367002 48288 367008 48300
rect 367060 48288 367066 48340
rect 389177 48331 389235 48337
rect 389177 48297 389189 48331
rect 389223 48328 389235 48331
rect 389266 48328 389272 48340
rect 389223 48300 389272 48328
rect 389223 48297 389235 48300
rect 389177 48291 389235 48297
rect 389266 48288 389272 48300
rect 389324 48288 389330 48340
rect 424505 48331 424563 48337
rect 424505 48297 424517 48331
rect 424551 48328 424563 48331
rect 424686 48328 424692 48340
rect 424551 48300 424692 48328
rect 424551 48297 424563 48300
rect 424505 48291 424563 48297
rect 424686 48288 424692 48300
rect 424744 48288 424750 48340
rect 470594 48328 470600 48340
rect 470555 48300 470600 48328
rect 470594 48288 470600 48300
rect 470652 48288 470658 48340
rect 236270 48260 236276 48272
rect 236231 48232 236276 48260
rect 236270 48220 236276 48232
rect 236328 48220 236334 48272
rect 273530 48260 273536 48272
rect 273491 48232 273536 48260
rect 273530 48220 273536 48232
rect 273588 48220 273594 48272
rect 325973 48195 326031 48201
rect 325973 48161 325985 48195
rect 326019 48192 326031 48195
rect 326062 48192 326068 48204
rect 326019 48164 326068 48192
rect 326019 48161 326031 48164
rect 325973 48155 326031 48161
rect 326062 48152 326068 48164
rect 326120 48152 326126 48204
rect 265250 46968 265256 46980
rect 265211 46940 265256 46968
rect 265250 46928 265256 46940
rect 265308 46928 265314 46980
rect 285950 46928 285956 46980
rect 286008 46968 286014 46980
rect 286045 46971 286103 46977
rect 286045 46968 286057 46971
rect 286008 46940 286057 46968
rect 286008 46928 286014 46940
rect 286045 46937 286057 46940
rect 286091 46937 286103 46971
rect 286045 46931 286103 46937
rect 337102 46928 337108 46980
rect 337160 46968 337166 46980
rect 337289 46971 337347 46977
rect 337289 46968 337301 46971
rect 337160 46940 337301 46968
rect 337160 46928 337166 46940
rect 337289 46937 337301 46940
rect 337335 46937 337347 46971
rect 421006 46968 421012 46980
rect 420967 46940 421012 46968
rect 337289 46931 337347 46937
rect 421006 46928 421012 46940
rect 421064 46928 421070 46980
rect 234982 46900 234988 46912
rect 234943 46872 234988 46900
rect 234982 46860 234988 46872
rect 235040 46860 235046 46912
rect 259638 46860 259644 46912
rect 259696 46900 259702 46912
rect 259730 46900 259736 46912
rect 259696 46872 259736 46900
rect 259696 46860 259702 46872
rect 259730 46860 259736 46872
rect 259788 46860 259794 46912
rect 301038 46860 301044 46912
rect 301096 46900 301102 46912
rect 301314 46900 301320 46912
rect 301096 46872 301320 46900
rect 301096 46860 301102 46872
rect 301314 46860 301320 46872
rect 301372 46860 301378 46912
rect 302510 46860 302516 46912
rect 302568 46900 302574 46912
rect 302602 46900 302608 46912
rect 302568 46872 302608 46900
rect 302568 46860 302574 46872
rect 302602 46860 302608 46872
rect 302660 46860 302666 46912
rect 327258 46900 327264 46912
rect 327219 46872 327264 46900
rect 327258 46860 327264 46872
rect 327316 46860 327322 46912
rect 330110 46900 330116 46912
rect 330071 46872 330116 46900
rect 330110 46860 330116 46872
rect 330168 46860 330174 46912
rect 336918 46900 336924 46912
rect 336879 46872 336924 46900
rect 336918 46860 336924 46872
rect 336976 46860 336982 46912
rect 341245 46903 341303 46909
rect 341245 46869 341257 46903
rect 341291 46900 341303 46903
rect 341426 46900 341432 46912
rect 341291 46872 341432 46900
rect 341291 46869 341303 46872
rect 341245 46863 341303 46869
rect 341426 46860 341432 46872
rect 341484 46860 341490 46912
rect 358633 46903 358691 46909
rect 358633 46869 358645 46903
rect 358679 46900 358691 46903
rect 358722 46900 358728 46912
rect 358679 46872 358728 46900
rect 358679 46869 358691 46872
rect 358633 46863 358691 46869
rect 358722 46860 358728 46872
rect 358780 46860 358786 46912
rect 359090 46900 359096 46912
rect 359051 46872 359096 46900
rect 359090 46860 359096 46872
rect 359148 46860 359154 46912
rect 267829 45951 267887 45957
rect 267829 45917 267841 45951
rect 267875 45948 267887 45951
rect 268102 45948 268108 45960
rect 267875 45920 268108 45948
rect 267875 45917 267887 45920
rect 267829 45911 267887 45917
rect 268102 45908 268108 45920
rect 268160 45908 268166 45960
rect 310882 45636 310888 45688
rect 310940 45676 310946 45688
rect 311066 45676 311072 45688
rect 310940 45648 311072 45676
rect 310940 45636 310946 45648
rect 311066 45636 311072 45648
rect 311124 45636 311130 45688
rect 267826 45608 267832 45620
rect 267787 45580 267832 45608
rect 267826 45568 267832 45580
rect 267884 45568 267890 45620
rect 265250 45540 265256 45552
rect 265211 45512 265256 45540
rect 265250 45500 265256 45512
rect 265308 45500 265314 45552
rect 290090 45500 290096 45552
rect 290148 45500 290154 45552
rect 291562 45500 291568 45552
rect 291620 45500 291626 45552
rect 296806 45540 296812 45552
rect 296767 45512 296812 45540
rect 296806 45500 296812 45512
rect 296864 45500 296870 45552
rect 301314 45540 301320 45552
rect 301275 45512 301320 45540
rect 301314 45500 301320 45512
rect 301372 45500 301378 45552
rect 307018 45540 307024 45552
rect 306979 45512 307024 45540
rect 307018 45500 307024 45512
rect 307076 45500 307082 45552
rect 310882 45500 310888 45552
rect 310940 45540 310946 45552
rect 311066 45540 311072 45552
rect 310940 45512 311072 45540
rect 310940 45500 310946 45512
rect 311066 45500 311072 45512
rect 311124 45500 311130 45552
rect 317506 45500 317512 45552
rect 317564 45540 317570 45552
rect 317690 45540 317696 45552
rect 317564 45512 317696 45540
rect 317564 45500 317570 45512
rect 317690 45500 317696 45512
rect 317748 45500 317754 45552
rect 288802 45432 288808 45484
rect 288860 45472 288866 45484
rect 289078 45472 289084 45484
rect 288860 45444 289084 45472
rect 288860 45432 288866 45444
rect 289078 45432 289084 45444
rect 289136 45432 289142 45484
rect 290108 45472 290136 45500
rect 290182 45472 290188 45484
rect 290108 45444 290188 45472
rect 290182 45432 290188 45444
rect 290240 45432 290246 45484
rect 291580 45472 291608 45500
rect 291654 45472 291660 45484
rect 291580 45444 291660 45472
rect 291654 45432 291660 45444
rect 291712 45432 291718 45484
rect 299750 42032 299756 42084
rect 299808 42072 299814 42084
rect 300118 42072 300124 42084
rect 299808 42044 300124 42072
rect 299808 42032 299814 42044
rect 300118 42032 300124 42044
rect 300176 42032 300182 42084
rect 421006 42032 421012 42084
rect 421064 42072 421070 42084
rect 421193 42075 421251 42081
rect 421193 42072 421205 42075
rect 421064 42044 421205 42072
rect 421064 42032 421070 42044
rect 421193 42041 421205 42044
rect 421239 42041 421251 42075
rect 421193 42035 421251 42041
rect 251450 41460 251456 41472
rect 251376 41432 251456 41460
rect 251376 41404 251404 41432
rect 251450 41420 251456 41432
rect 251508 41420 251514 41472
rect 284754 41460 284760 41472
rect 284680 41432 284760 41460
rect 284680 41404 284708 41432
rect 284754 41420 284760 41432
rect 284812 41420 284818 41472
rect 362218 41460 362224 41472
rect 362179 41432 362224 41460
rect 362218 41420 362224 41432
rect 362276 41420 362282 41472
rect 251358 41352 251364 41404
rect 251416 41352 251422 41404
rect 284662 41352 284668 41404
rect 284720 41352 284726 41404
rect 360286 41352 360292 41404
rect 360344 41392 360350 41404
rect 360470 41392 360476 41404
rect 360344 41364 360476 41392
rect 360344 41352 360350 41364
rect 360470 41352 360476 41364
rect 360528 41352 360534 41404
rect 388990 41352 388996 41404
rect 389048 41392 389054 41404
rect 389358 41392 389364 41404
rect 389048 41364 389364 41392
rect 389048 41352 389054 41364
rect 389358 41352 389364 41364
rect 389416 41352 389422 41404
rect 239122 41324 239128 41336
rect 239083 41296 239128 41324
rect 239122 41284 239128 41296
rect 239180 41284 239186 41336
rect 377122 41324 377128 41336
rect 377083 41296 377128 41324
rect 377122 41284 377128 41296
rect 377180 41284 377186 41336
rect 396074 40196 396080 40248
rect 396132 40236 396138 40248
rect 399018 40236 399024 40248
rect 396132 40208 399024 40236
rect 396132 40196 396138 40208
rect 399018 40196 399024 40208
rect 399076 40196 399082 40248
rect 437198 40196 437204 40248
rect 437256 40236 437262 40248
rect 437474 40236 437480 40248
rect 437256 40208 437480 40236
rect 437256 40196 437262 40208
rect 437474 40196 437480 40208
rect 437532 40196 437538 40248
rect 303798 40168 303804 40180
rect 303759 40140 303804 40168
rect 303798 40128 303804 40140
rect 303856 40128 303862 40180
rect 306374 40128 306380 40180
rect 306432 40168 306438 40180
rect 315942 40168 315948 40180
rect 306432 40140 315948 40168
rect 306432 40128 306438 40140
rect 315942 40128 315948 40140
rect 316000 40128 316006 40180
rect 417878 40128 417884 40180
rect 417936 40168 417942 40180
rect 418246 40168 418252 40180
rect 417936 40140 418252 40168
rect 417936 40128 417942 40140
rect 418246 40128 418252 40140
rect 418304 40128 418310 40180
rect 456518 40128 456524 40180
rect 456576 40168 456582 40180
rect 456886 40168 456892 40180
rect 456576 40140 456892 40168
rect 456576 40128 456582 40140
rect 456886 40128 456892 40140
rect 456944 40128 456950 40180
rect 232314 38700 232320 38752
rect 232372 38740 232378 38752
rect 232406 38740 232412 38752
rect 232372 38712 232412 38740
rect 232372 38700 232378 38712
rect 232406 38700 232412 38712
rect 232464 38700 232470 38752
rect 244366 38700 244372 38752
rect 244424 38700 244430 38752
rect 377030 38700 377036 38752
rect 377088 38740 377094 38752
rect 377125 38743 377183 38749
rect 377125 38740 377137 38743
rect 377088 38712 377137 38740
rect 377088 38700 377094 38712
rect 377125 38709 377137 38712
rect 377171 38709 377183 38743
rect 377125 38703 377183 38709
rect 244384 38672 244412 38700
rect 244458 38672 244464 38684
rect 244384 38644 244464 38672
rect 244458 38632 244464 38644
rect 244516 38632 244522 38684
rect 245562 38632 245568 38684
rect 245620 38672 245626 38684
rect 245930 38672 245936 38684
rect 245620 38644 245936 38672
rect 245620 38632 245626 38644
rect 245930 38632 245936 38644
rect 245988 38632 245994 38684
rect 270678 38632 270684 38684
rect 270736 38672 270742 38684
rect 270770 38672 270776 38684
rect 270736 38644 270776 38672
rect 270736 38632 270742 38644
rect 270770 38632 270776 38644
rect 270828 38632 270834 38684
rect 272150 38632 272156 38684
rect 272208 38672 272214 38684
rect 272242 38672 272248 38684
rect 272208 38644 272248 38672
rect 272208 38632 272214 38644
rect 272242 38632 272248 38644
rect 272300 38632 272306 38684
rect 273530 38672 273536 38684
rect 273491 38644 273536 38672
rect 273530 38632 273536 38644
rect 273588 38632 273594 38684
rect 323302 38632 323308 38684
rect 323360 38632 323366 38684
rect 296806 38604 296812 38616
rect 296767 38576 296812 38604
rect 296806 38564 296812 38576
rect 296864 38564 296870 38616
rect 323320 38536 323348 38632
rect 362218 38604 362224 38616
rect 362179 38576 362224 38604
rect 362218 38564 362224 38576
rect 362276 38564 362282 38616
rect 367002 38604 367008 38616
rect 366963 38576 367008 38604
rect 367002 38564 367008 38576
rect 367060 38564 367066 38616
rect 424502 38604 424508 38616
rect 424463 38576 424508 38604
rect 424502 38564 424508 38576
rect 424560 38564 424566 38616
rect 323394 38536 323400 38548
rect 323320 38508 323400 38536
rect 323394 38496 323400 38508
rect 323452 38496 323458 38548
rect 234985 37315 235043 37321
rect 234985 37281 234997 37315
rect 235031 37312 235043 37315
rect 235074 37312 235080 37324
rect 235031 37284 235080 37312
rect 235031 37281 235043 37284
rect 234985 37275 235043 37281
rect 235074 37272 235080 37284
rect 235132 37272 235138 37324
rect 236270 37312 236276 37324
rect 236231 37284 236276 37312
rect 236270 37272 236276 37284
rect 236328 37272 236334 37324
rect 239122 37312 239128 37324
rect 239083 37284 239128 37312
rect 239122 37272 239128 37284
rect 239180 37272 239186 37324
rect 325970 37272 325976 37324
rect 326028 37312 326034 37324
rect 326062 37312 326068 37324
rect 326028 37284 326068 37312
rect 326028 37272 326034 37284
rect 326062 37272 326068 37284
rect 326120 37272 326126 37324
rect 327258 37312 327264 37324
rect 327219 37284 327264 37312
rect 327258 37272 327264 37284
rect 327316 37272 327322 37324
rect 330110 37312 330116 37324
rect 330071 37284 330116 37312
rect 330110 37272 330116 37284
rect 330168 37272 330174 37324
rect 336918 37312 336924 37324
rect 336879 37284 336924 37312
rect 336918 37272 336924 37284
rect 336976 37272 336982 37324
rect 341242 37312 341248 37324
rect 341203 37284 341248 37312
rect 341242 37272 341248 37284
rect 341300 37272 341306 37324
rect 357526 37272 357532 37324
rect 357584 37312 357590 37324
rect 357710 37312 357716 37324
rect 357584 37284 357716 37312
rect 357584 37272 357590 37284
rect 357710 37272 357716 37284
rect 357768 37272 357774 37324
rect 358630 37312 358636 37324
rect 358591 37284 358636 37312
rect 358630 37272 358636 37284
rect 358688 37272 358694 37324
rect 359093 37315 359151 37321
rect 359093 37281 359105 37315
rect 359139 37312 359151 37315
rect 359182 37312 359188 37324
rect 359139 37284 359188 37312
rect 359139 37281 359151 37284
rect 359093 37275 359151 37281
rect 359182 37272 359188 37284
rect 359240 37272 359246 37324
rect 244369 37247 244427 37253
rect 244369 37213 244381 37247
rect 244415 37244 244427 37247
rect 244458 37244 244464 37256
rect 244415 37216 244464 37244
rect 244415 37213 244427 37216
rect 244369 37207 244427 37213
rect 244458 37204 244464 37216
rect 244516 37204 244522 37256
rect 245841 37247 245899 37253
rect 245841 37213 245853 37247
rect 245887 37244 245899 37247
rect 245930 37244 245936 37256
rect 245887 37216 245936 37244
rect 245887 37213 245899 37216
rect 245841 37207 245899 37213
rect 245930 37204 245936 37216
rect 245988 37204 245994 37256
rect 267826 37204 267832 37256
rect 267884 37244 267890 37256
rect 268010 37244 268016 37256
rect 267884 37216 268016 37244
rect 267884 37204 267890 37216
rect 268010 37204 268016 37216
rect 268068 37204 268074 37256
rect 337105 37247 337163 37253
rect 337105 37213 337117 37247
rect 337151 37244 337163 37247
rect 337194 37244 337200 37256
rect 337151 37216 337200 37244
rect 337151 37213 337163 37216
rect 337105 37207 337163 37213
rect 337194 37204 337200 37216
rect 337252 37204 337258 37256
rect 265250 35952 265256 35964
rect 265211 35924 265256 35952
rect 265250 35912 265256 35924
rect 265308 35912 265314 35964
rect 294138 35912 294144 35964
rect 294196 35952 294202 35964
rect 294230 35952 294236 35964
rect 294196 35924 294236 35952
rect 294196 35912 294202 35924
rect 294230 35912 294236 35924
rect 294288 35912 294294 35964
rect 301314 35952 301320 35964
rect 301275 35924 301320 35952
rect 301314 35912 301320 35924
rect 301372 35912 301378 35964
rect 307018 35952 307024 35964
rect 306979 35924 307024 35952
rect 307018 35912 307024 35924
rect 307076 35912 307082 35964
rect 3142 35844 3148 35896
rect 3200 35884 3206 35896
rect 6178 35884 6184 35896
rect 3200 35856 6184 35884
rect 3200 35844 3206 35856
rect 6178 35844 6184 35856
rect 6236 35844 6242 35896
rect 336734 33804 336740 33856
rect 336792 33844 336798 33856
rect 336918 33844 336924 33856
rect 336792 33816 336924 33844
rect 336792 33804 336798 33816
rect 336918 33804 336924 33816
rect 336976 33804 336982 33856
rect 303801 32419 303859 32425
rect 303801 32385 303813 32419
rect 303847 32416 303859 32419
rect 303890 32416 303896 32428
rect 303847 32388 303896 32416
rect 303847 32385 303859 32388
rect 303801 32379 303859 32385
rect 303890 32376 303896 32388
rect 303948 32376 303954 32428
rect 377122 31968 377128 32020
rect 377180 32008 377186 32020
rect 377306 32008 377312 32020
rect 377180 31980 377312 32008
rect 377180 31968 377186 31980
rect 377306 31968 377312 31980
rect 377364 31968 377370 32020
rect 265250 31764 265256 31816
rect 265308 31764 265314 31816
rect 317506 31764 317512 31816
rect 317564 31804 317570 31816
rect 317690 31804 317696 31816
rect 317564 31776 317696 31804
rect 317564 31764 317570 31776
rect 317690 31764 317696 31776
rect 317748 31764 317754 31816
rect 327258 31764 327264 31816
rect 327316 31764 327322 31816
rect 265268 31680 265296 31764
rect 265250 31628 265256 31680
rect 265308 31628 265314 31680
rect 327276 31612 327304 31764
rect 389358 31696 389364 31748
rect 389416 31736 389422 31748
rect 389542 31736 389548 31748
rect 389416 31708 389548 31736
rect 389416 31696 389422 31708
rect 389542 31696 389548 31708
rect 389600 31696 389606 31748
rect 266630 31560 266636 31612
rect 266688 31600 266694 31612
rect 266814 31600 266820 31612
rect 266688 31572 266820 31600
rect 266688 31560 266694 31572
rect 266814 31560 266820 31572
rect 266872 31560 266878 31612
rect 327258 31560 327264 31612
rect 327316 31560 327322 31612
rect 288805 29835 288863 29841
rect 288805 29801 288817 29835
rect 288851 29832 288863 29835
rect 289078 29832 289084 29844
rect 288851 29804 289084 29832
rect 288851 29801 288863 29804
rect 288805 29795 288863 29801
rect 289078 29792 289084 29804
rect 289136 29792 289142 29844
rect 267734 29180 267740 29232
rect 267792 29220 267798 29232
rect 277302 29220 277308 29232
rect 267792 29192 277308 29220
rect 267792 29180 267798 29192
rect 277302 29180 277308 29192
rect 277360 29180 277366 29232
rect 456518 29180 456524 29232
rect 456576 29220 456582 29232
rect 456978 29220 456984 29232
rect 456576 29192 456984 29220
rect 456576 29180 456582 29192
rect 456978 29180 456984 29192
rect 457036 29180 457042 29232
rect 238754 29112 238760 29164
rect 238812 29152 238818 29164
rect 256602 29152 256608 29164
rect 238812 29124 256608 29152
rect 238812 29112 238818 29124
rect 256602 29112 256608 29124
rect 256660 29112 256666 29164
rect 437198 29112 437204 29164
rect 437256 29152 437262 29164
rect 437474 29152 437480 29164
rect 437256 29124 437480 29152
rect 437256 29112 437262 29124
rect 437474 29112 437480 29124
rect 437532 29112 437538 29164
rect 286042 29084 286048 29096
rect 285968 29056 286048 29084
rect 285968 29028 285996 29056
rect 286042 29044 286048 29056
rect 286100 29044 286106 29096
rect 347774 29044 347780 29096
rect 347832 29084 347838 29096
rect 357342 29084 357348 29096
rect 347832 29056 357348 29084
rect 347832 29044 347838 29056
rect 357342 29044 357348 29056
rect 357400 29044 357406 29096
rect 359182 29044 359188 29096
rect 359240 29044 359246 29096
rect 367002 29084 367008 29096
rect 366963 29056 367008 29084
rect 367002 29044 367008 29056
rect 367060 29044 367066 29096
rect 492766 29044 492772 29096
rect 492824 29084 492830 29096
rect 502242 29084 502248 29096
rect 492824 29056 502248 29084
rect 492824 29044 492830 29056
rect 502242 29044 502248 29056
rect 502300 29044 502306 29096
rect 232222 28976 232228 29028
rect 232280 29016 232286 29028
rect 232406 29016 232412 29028
rect 232280 28988 232412 29016
rect 232280 28976 232286 28988
rect 232406 28976 232412 28988
rect 232464 28976 232470 29028
rect 284662 28976 284668 29028
rect 284720 29016 284726 29028
rect 284754 29016 284760 29028
rect 284720 28988 284760 29016
rect 284720 28976 284726 28988
rect 284754 28976 284760 28988
rect 284812 28976 284818 29028
rect 285950 28976 285956 29028
rect 286008 28976 286014 29028
rect 325970 28976 325976 29028
rect 326028 29016 326034 29028
rect 326062 29016 326068 29028
rect 326028 28988 326068 29016
rect 326028 28976 326034 28988
rect 326062 28976 326068 28988
rect 326120 28976 326126 29028
rect 358630 28976 358636 29028
rect 358688 29016 358694 29028
rect 358722 29016 358728 29028
rect 358688 28988 358728 29016
rect 358688 28976 358694 28988
rect 358722 28976 358728 28988
rect 358780 28976 358786 29028
rect 359200 28960 359228 29044
rect 424505 29019 424563 29025
rect 424505 28985 424517 29019
rect 424551 29016 424563 29019
rect 424594 29016 424600 29028
rect 424551 28988 424600 29016
rect 424551 28985 424563 28988
rect 424505 28979 424563 28985
rect 424594 28976 424600 28988
rect 424652 28976 424658 29028
rect 295518 28908 295524 28960
rect 295576 28948 295582 28960
rect 295610 28948 295616 28960
rect 295576 28920 295616 28948
rect 295576 28908 295582 28920
rect 295610 28908 295616 28920
rect 295668 28908 295674 28960
rect 323302 28908 323308 28960
rect 323360 28948 323366 28960
rect 323394 28948 323400 28960
rect 323360 28920 323400 28948
rect 323360 28908 323366 28920
rect 323394 28908 323400 28920
rect 323452 28908 323458 28960
rect 324590 28908 324596 28960
rect 324648 28948 324654 28960
rect 324682 28948 324688 28960
rect 324648 28920 324688 28948
rect 324648 28908 324654 28920
rect 324682 28908 324688 28920
rect 324740 28908 324746 28960
rect 359182 28908 359188 28960
rect 359240 28908 359246 28960
rect 367002 28948 367008 28960
rect 366963 28920 367008 28948
rect 367002 28908 367008 28920
rect 367060 28908 367066 28960
rect 389453 28951 389511 28957
rect 389453 28917 389465 28951
rect 389499 28948 389511 28951
rect 389542 28948 389548 28960
rect 389499 28920 389548 28948
rect 389499 28917 389511 28920
rect 389453 28911 389511 28917
rect 389542 28908 389548 28920
rect 389600 28908 389606 28960
rect 306374 28772 306380 28824
rect 306432 28812 306438 28824
rect 315942 28812 315948 28824
rect 306432 28784 315948 28812
rect 306432 28772 306438 28784
rect 315942 28772 315948 28784
rect 316000 28772 316006 28824
rect 244366 28064 244372 28076
rect 244327 28036 244372 28064
rect 244366 28024 244372 28036
rect 244424 28024 244430 28076
rect 268010 27724 268016 27736
rect 267936 27696 268016 27724
rect 245838 27656 245844 27668
rect 245799 27628 245844 27656
rect 245838 27616 245844 27628
rect 245896 27616 245902 27668
rect 267936 27600 267964 27696
rect 268010 27684 268016 27696
rect 268068 27684 268074 27736
rect 341242 27724 341248 27736
rect 341168 27696 341248 27724
rect 341168 27668 341196 27696
rect 341242 27684 341248 27696
rect 341300 27684 341306 27736
rect 337102 27656 337108 27668
rect 337063 27628 337108 27656
rect 337102 27616 337108 27628
rect 337160 27616 337166 27668
rect 341150 27616 341156 27668
rect 341208 27616 341214 27668
rect 421006 27616 421012 27668
rect 421064 27656 421070 27668
rect 421193 27659 421251 27665
rect 421193 27656 421205 27659
rect 421064 27628 421205 27656
rect 421064 27616 421070 27628
rect 421193 27625 421205 27628
rect 421239 27625 421251 27659
rect 421193 27619 421251 27625
rect 236270 27588 236276 27600
rect 236231 27560 236276 27588
rect 236270 27548 236276 27560
rect 236328 27548 236334 27600
rect 265250 27588 265256 27600
rect 265211 27560 265256 27588
rect 265250 27548 265256 27560
rect 265308 27548 265314 27600
rect 267918 27548 267924 27600
rect 267976 27548 267982 27600
rect 284573 27591 284631 27597
rect 284573 27557 284585 27591
rect 284619 27588 284631 27591
rect 284754 27588 284760 27600
rect 284619 27560 284760 27588
rect 284619 27557 284631 27560
rect 284573 27551 284631 27557
rect 284754 27548 284760 27560
rect 284812 27548 284818 27600
rect 285950 27588 285956 27600
rect 285911 27560 285956 27588
rect 285950 27548 285956 27560
rect 286008 27548 286014 27600
rect 299750 27548 299756 27600
rect 299808 27588 299814 27600
rect 299934 27588 299940 27600
rect 299808 27560 299940 27588
rect 299808 27548 299814 27560
rect 299934 27548 299940 27560
rect 299992 27548 299998 27600
rect 301130 27548 301136 27600
rect 301188 27588 301194 27600
rect 301222 27588 301228 27600
rect 301188 27560 301228 27588
rect 301188 27548 301194 27560
rect 301222 27548 301228 27560
rect 301280 27548 301286 27600
rect 306926 27548 306932 27600
rect 306984 27548 306990 27600
rect 358541 27591 358599 27597
rect 358541 27557 358553 27591
rect 358587 27588 358599 27591
rect 358722 27588 358728 27600
rect 358587 27560 358728 27588
rect 358587 27557 358599 27560
rect 358541 27551 358599 27557
rect 358722 27548 358728 27560
rect 358780 27548 358786 27600
rect 306834 27480 306840 27532
rect 306892 27520 306898 27532
rect 306944 27520 306972 27548
rect 306892 27492 306972 27520
rect 306892 27480 306898 27492
rect 244185 26231 244243 26237
rect 244185 26197 244197 26231
rect 244231 26228 244243 26231
rect 244366 26228 244372 26240
rect 244231 26200 244372 26228
rect 244231 26197 244243 26200
rect 244185 26191 244243 26197
rect 244366 26188 244372 26200
rect 244424 26188 244430 26240
rect 245838 26228 245844 26240
rect 245799 26200 245844 26228
rect 245838 26188 245844 26200
rect 245896 26188 245902 26240
rect 249978 26188 249984 26240
rect 250036 26228 250042 26240
rect 250162 26228 250168 26240
rect 250036 26200 250168 26228
rect 250036 26188 250042 26200
rect 250162 26188 250168 26200
rect 250220 26188 250226 26240
rect 267737 26231 267795 26237
rect 267737 26197 267749 26231
rect 267783 26228 267795 26231
rect 267918 26228 267924 26240
rect 267783 26200 267924 26228
rect 267783 26197 267795 26200
rect 267737 26191 267795 26197
rect 267918 26188 267924 26200
rect 267976 26188 267982 26240
rect 299750 26228 299756 26240
rect 299711 26200 299756 26228
rect 299750 26188 299756 26200
rect 299808 26188 299814 26240
rect 341150 26188 341156 26240
rect 341208 26228 341214 26240
rect 341245 26231 341303 26237
rect 341245 26228 341257 26231
rect 341208 26200 341257 26228
rect 341208 26188 341214 26200
rect 341245 26197 341257 26200
rect 341291 26197 341303 26231
rect 341245 26191 341303 26197
rect 421006 22720 421012 22772
rect 421064 22760 421070 22772
rect 421193 22763 421251 22769
rect 421193 22760 421205 22763
rect 421064 22732 421205 22760
rect 421064 22720 421070 22732
rect 421193 22729 421205 22732
rect 421239 22729 421251 22763
rect 421193 22723 421251 22729
rect 270494 22108 270500 22160
rect 270552 22148 270558 22160
rect 270770 22148 270776 22160
rect 270552 22120 270776 22148
rect 270552 22108 270558 22120
rect 270770 22108 270776 22120
rect 270828 22108 270834 22160
rect 377030 22108 377036 22160
rect 377088 22108 377094 22160
rect 424594 22148 424600 22160
rect 424520 22120 424600 22148
rect 377048 22012 377076 22108
rect 424520 22092 424548 22120
rect 424594 22108 424600 22120
rect 424652 22108 424658 22160
rect 424502 22040 424508 22092
rect 424560 22040 424566 22092
rect 377122 22012 377128 22024
rect 377048 21984 377128 22012
rect 377122 21972 377128 21984
rect 377180 21972 377186 22024
rect 232406 19320 232412 19372
rect 232464 19320 232470 19372
rect 302510 19320 302516 19372
rect 302568 19360 302574 19372
rect 302602 19360 302608 19372
rect 302568 19332 302608 19360
rect 302568 19320 302574 19332
rect 302602 19320 302608 19332
rect 302660 19320 302666 19372
rect 336734 19320 336740 19372
rect 336792 19360 336798 19372
rect 336918 19360 336924 19372
rect 336792 19332 336924 19360
rect 336792 19320 336798 19332
rect 336918 19320 336924 19332
rect 336976 19320 336982 19372
rect 367002 19360 367008 19372
rect 366963 19332 367008 19360
rect 367002 19320 367008 19332
rect 367060 19320 367066 19372
rect 389450 19360 389456 19372
rect 389411 19332 389456 19360
rect 389450 19320 389456 19332
rect 389508 19320 389514 19372
rect 232424 19224 232452 19320
rect 265250 19292 265256 19304
rect 265211 19264 265256 19292
rect 265250 19252 265256 19264
rect 265308 19252 265314 19304
rect 288802 19292 288808 19304
rect 288763 19264 288808 19292
rect 288802 19252 288808 19264
rect 288860 19252 288866 19304
rect 325970 19252 325976 19304
rect 326028 19252 326034 19304
rect 327258 19252 327264 19304
rect 327316 19252 327322 19304
rect 366910 19292 366916 19304
rect 366871 19264 366916 19292
rect 366910 19252 366916 19264
rect 366968 19252 366974 19304
rect 232498 19224 232504 19236
rect 232424 19196 232504 19224
rect 232498 19184 232504 19196
rect 232556 19184 232562 19236
rect 325988 19168 326016 19252
rect 327276 19168 327304 19252
rect 325970 19116 325976 19168
rect 326028 19116 326034 19168
rect 327258 19116 327264 19168
rect 327316 19116 327322 19168
rect 362221 18071 362279 18077
rect 362221 18037 362233 18071
rect 362267 18068 362279 18071
rect 362310 18068 362316 18080
rect 362267 18040 362316 18068
rect 362267 18037 362279 18040
rect 362221 18031 362279 18037
rect 362310 18028 362316 18040
rect 362368 18028 362374 18080
rect 236270 18000 236276 18012
rect 236231 17972 236276 18000
rect 236270 17960 236276 17972
rect 236328 17960 236334 18012
rect 270586 17960 270592 18012
rect 270644 17960 270650 18012
rect 271966 17960 271972 18012
rect 272024 17960 272030 18012
rect 284570 18000 284576 18012
rect 284531 17972 284576 18000
rect 284570 17960 284576 17972
rect 284628 17960 284634 18012
rect 285950 18000 285956 18012
rect 285911 17972 285956 18000
rect 285950 17960 285956 17972
rect 286008 17960 286014 18012
rect 294138 17960 294144 18012
rect 294196 18000 294202 18012
rect 294230 18000 294236 18012
rect 294196 17972 294236 18000
rect 294196 17960 294202 17972
rect 294230 17960 294236 17972
rect 294288 17960 294294 18012
rect 265250 17892 265256 17944
rect 265308 17932 265314 17944
rect 265434 17932 265440 17944
rect 265308 17904 265440 17932
rect 265308 17892 265314 17904
rect 265434 17892 265440 17904
rect 265492 17892 265498 17944
rect 270604 17876 270632 17960
rect 271984 17876 272012 17960
rect 273438 17932 273444 17944
rect 273399 17904 273444 17932
rect 273438 17892 273444 17904
rect 273496 17892 273502 17944
rect 376757 17935 376815 17941
rect 376757 17901 376769 17935
rect 376803 17932 376815 17935
rect 377122 17932 377128 17944
rect 376803 17904 377128 17932
rect 376803 17901 376815 17904
rect 376757 17895 376815 17901
rect 377122 17892 377128 17904
rect 377180 17892 377186 17944
rect 270586 17824 270592 17876
rect 270644 17824 270650 17876
rect 271966 17824 271972 17876
rect 272024 17824 272030 17876
rect 271874 17756 271880 17808
rect 271932 17796 271938 17808
rect 272334 17796 272340 17808
rect 271932 17768 272340 17796
rect 271932 17756 271938 17768
rect 272334 17756 272340 17768
rect 272392 17756 272398 17808
rect 395982 17144 395988 17196
rect 396040 17144 396046 17196
rect 306374 17008 306380 17060
rect 306432 17048 306438 17060
rect 315942 17048 315948 17060
rect 306432 17020 315948 17048
rect 306432 17008 306438 17020
rect 315942 17008 315948 17020
rect 316000 17008 316006 17060
rect 396000 16992 396028 17144
rect 395982 16940 395988 16992
rect 396040 16940 396046 16992
rect 347774 16872 347780 16924
rect 347832 16912 347838 16924
rect 352650 16912 352656 16924
rect 347832 16884 352656 16912
rect 347832 16872 347838 16884
rect 352650 16872 352656 16884
rect 352708 16872 352714 16924
rect 385126 16804 385132 16856
rect 385184 16844 385190 16856
rect 395890 16844 395896 16856
rect 385184 16816 395896 16844
rect 385184 16804 385190 16816
rect 395890 16804 395896 16816
rect 395948 16804 395954 16856
rect 417878 16804 417884 16856
rect 417936 16844 417942 16856
rect 418246 16844 418252 16856
rect 417936 16816 418252 16844
rect 417936 16804 417942 16816
rect 418246 16804 418252 16816
rect 418304 16804 418310 16856
rect 456518 16804 456524 16856
rect 456576 16844 456582 16856
rect 458818 16844 458824 16856
rect 456576 16816 458824 16844
rect 456576 16804 456582 16816
rect 458818 16804 458824 16816
rect 458876 16804 458882 16856
rect 289262 16736 289268 16788
rect 289320 16776 289326 16788
rect 289906 16776 289912 16788
rect 289320 16748 289912 16776
rect 289320 16736 289326 16748
rect 289906 16736 289912 16748
rect 289964 16736 289970 16788
rect 437198 16736 437204 16788
rect 437256 16776 437262 16788
rect 437474 16776 437480 16788
rect 437256 16748 437480 16776
rect 437256 16736 437262 16748
rect 437474 16736 437480 16748
rect 437532 16736 437538 16788
rect 310974 16708 310980 16720
rect 310808 16680 310980 16708
rect 310808 16652 310836 16680
rect 310974 16668 310980 16680
rect 311032 16668 311038 16720
rect 244182 16640 244188 16652
rect 244143 16612 244188 16640
rect 244182 16600 244188 16612
rect 244240 16600 244246 16652
rect 245841 16643 245899 16649
rect 245841 16609 245853 16643
rect 245887 16640 245899 16643
rect 246022 16640 246028 16652
rect 245887 16612 246028 16640
rect 245887 16609 245899 16612
rect 245841 16603 245899 16609
rect 246022 16600 246028 16612
rect 246080 16600 246086 16652
rect 299750 16640 299756 16652
rect 299711 16612 299756 16640
rect 299750 16600 299756 16612
rect 299808 16600 299814 16652
rect 310790 16600 310796 16652
rect 310848 16600 310854 16652
rect 298094 16532 298100 16584
rect 298152 16572 298158 16584
rect 298462 16572 298468 16584
rect 298152 16544 298468 16572
rect 298152 16532 298158 16544
rect 298462 16532 298468 16544
rect 298520 16532 298526 16584
rect 110322 15104 110328 15156
rect 110380 15144 110386 15156
rect 274726 15144 274732 15156
rect 110380 15116 274732 15144
rect 110380 15104 110386 15116
rect 274726 15104 274732 15116
rect 274784 15104 274790 15156
rect 107470 15036 107476 15088
rect 107528 15076 107534 15088
rect 273346 15076 273352 15088
rect 107528 15048 273352 15076
rect 107528 15036 107534 15048
rect 273346 15036 273352 15048
rect 273404 15036 273410 15088
rect 103422 14968 103428 15020
rect 103480 15008 103486 15020
rect 271966 15008 271972 15020
rect 103480 14980 271972 15008
rect 103480 14968 103486 14980
rect 271966 14968 271972 14980
rect 272024 14968 272030 15020
rect 99282 14900 99288 14952
rect 99340 14940 99346 14952
rect 270586 14940 270592 14952
rect 99340 14912 270592 14940
rect 99340 14900 99346 14912
rect 270586 14900 270592 14912
rect 270644 14900 270650 14952
rect 96522 14832 96528 14884
rect 96580 14872 96586 14884
rect 269206 14872 269212 14884
rect 96580 14844 269212 14872
rect 96580 14832 96586 14844
rect 269206 14832 269212 14844
rect 269264 14832 269270 14884
rect 92382 14764 92388 14816
rect 92440 14804 92446 14816
rect 266446 14804 266452 14816
rect 92440 14776 266452 14804
rect 92440 14764 92446 14776
rect 266446 14764 266452 14776
rect 266504 14764 266510 14816
rect 89622 14696 89628 14748
rect 89680 14736 89686 14748
rect 265066 14736 265072 14748
rect 89680 14708 265072 14736
rect 89680 14696 89686 14708
rect 265066 14696 265072 14708
rect 265124 14696 265130 14748
rect 85482 14628 85488 14680
rect 85540 14668 85546 14680
rect 263686 14668 263692 14680
rect 85540 14640 263692 14668
rect 85540 14628 85546 14640
rect 263686 14628 263692 14640
rect 263744 14628 263750 14680
rect 82722 14560 82728 14612
rect 82780 14600 82786 14612
rect 262582 14600 262588 14612
rect 82780 14572 262588 14600
rect 82780 14560 82786 14572
rect 262582 14560 262588 14572
rect 262640 14560 262646 14612
rect 78582 14492 78588 14544
rect 78640 14532 78646 14544
rect 260926 14532 260932 14544
rect 78640 14504 260932 14532
rect 78640 14492 78646 14504
rect 260926 14492 260932 14504
rect 260984 14492 260990 14544
rect 74442 14424 74448 14476
rect 74500 14464 74506 14476
rect 259638 14464 259644 14476
rect 74500 14436 259644 14464
rect 74500 14424 74506 14436
rect 259638 14424 259644 14436
rect 259696 14424 259702 14476
rect 114462 14356 114468 14408
rect 114520 14396 114526 14408
rect 276106 14396 276112 14408
rect 114520 14368 276112 14396
rect 114520 14356 114526 14368
rect 276106 14356 276112 14368
rect 276164 14356 276170 14408
rect 366818 14356 366824 14408
rect 366876 14396 366882 14408
rect 367002 14396 367008 14408
rect 366876 14368 367008 14396
rect 366876 14356 366882 14368
rect 367002 14356 367008 14368
rect 367060 14356 367066 14408
rect 117222 14288 117228 14340
rect 117280 14328 117286 14340
rect 277670 14328 277676 14340
rect 117280 14300 277676 14328
rect 117280 14288 117286 14300
rect 277670 14288 277676 14300
rect 277728 14288 277734 14340
rect 121362 14220 121368 14272
rect 121420 14260 121426 14272
rect 278774 14260 278780 14272
rect 121420 14232 278780 14260
rect 121420 14220 121426 14232
rect 278774 14220 278780 14232
rect 278832 14220 278838 14272
rect 125410 14152 125416 14204
rect 125468 14192 125474 14204
rect 280246 14192 280252 14204
rect 125468 14164 280252 14192
rect 125468 14152 125474 14164
rect 280246 14152 280252 14164
rect 280304 14152 280310 14204
rect 232130 14084 232136 14136
rect 232188 14124 232194 14136
rect 232498 14124 232504 14136
rect 232188 14096 232504 14124
rect 232188 14084 232194 14096
rect 232498 14084 232504 14096
rect 232556 14084 232562 14136
rect 183462 13744 183468 13796
rect 183520 13784 183526 13796
rect 303890 13784 303896 13796
rect 183520 13756 303896 13784
rect 183520 13744 183526 13756
rect 303890 13744 303896 13756
rect 303948 13744 303954 13796
rect 186222 13676 186228 13728
rect 186280 13716 186286 13728
rect 306558 13716 306564 13728
rect 186280 13688 306564 13716
rect 186280 13676 186286 13688
rect 306558 13676 306564 13688
rect 306616 13676 306622 13728
rect 179322 13608 179328 13660
rect 179380 13648 179386 13660
rect 302510 13648 302516 13660
rect 179380 13620 302516 13648
rect 179380 13608 179386 13620
rect 302510 13608 302516 13620
rect 302568 13608 302574 13660
rect 176562 13540 176568 13592
rect 176620 13580 176626 13592
rect 301130 13580 301136 13592
rect 176620 13552 301136 13580
rect 176620 13540 176626 13552
rect 301130 13540 301136 13552
rect 301188 13540 301194 13592
rect 172422 13472 172428 13524
rect 172480 13512 172486 13524
rect 299750 13512 299756 13524
rect 172480 13484 299756 13512
rect 172480 13472 172486 13484
rect 299750 13472 299756 13484
rect 299808 13472 299814 13524
rect 168282 13404 168288 13456
rect 168340 13444 168346 13456
rect 298278 13444 298284 13456
rect 168340 13416 298284 13444
rect 168340 13404 168346 13416
rect 298278 13404 298284 13416
rect 298336 13404 298342 13456
rect 165522 13336 165528 13388
rect 165580 13376 165586 13388
rect 296898 13376 296904 13388
rect 165580 13348 296904 13376
rect 165580 13336 165586 13348
rect 296898 13336 296904 13348
rect 296956 13336 296962 13388
rect 160002 13268 160008 13320
rect 160060 13308 160066 13320
rect 294230 13308 294236 13320
rect 160060 13280 294236 13308
rect 160060 13268 160066 13280
rect 294230 13268 294236 13280
rect 294288 13268 294294 13320
rect 155862 13200 155868 13252
rect 155920 13240 155926 13252
rect 292758 13240 292764 13252
rect 155920 13212 292764 13240
rect 155920 13200 155926 13212
rect 292758 13200 292764 13212
rect 292816 13200 292822 13252
rect 71682 13132 71688 13184
rect 71740 13172 71746 13184
rect 258166 13172 258172 13184
rect 71740 13144 258172 13172
rect 71740 13132 71746 13144
rect 258166 13132 258172 13144
rect 258224 13132 258230 13184
rect 31662 13064 31668 13116
rect 31720 13104 31726 13116
rect 241606 13104 241612 13116
rect 31720 13076 241612 13104
rect 31720 13064 31726 13076
rect 241606 13064 241612 13076
rect 241664 13064 241670 13116
rect 245838 13064 245844 13116
rect 245896 13104 245902 13116
rect 246022 13104 246028 13116
rect 245896 13076 246028 13104
rect 245896 13064 245902 13076
rect 246022 13064 246028 13076
rect 246080 13064 246086 13116
rect 190362 12996 190368 13048
rect 190420 13036 190426 13048
rect 307938 13036 307944 13048
rect 190420 13008 307944 13036
rect 190420 12996 190426 13008
rect 307938 12996 307944 13008
rect 307996 12996 308002 13048
rect 206922 12928 206928 12980
rect 206980 12968 206986 12980
rect 314838 12968 314844 12980
rect 206980 12940 314844 12968
rect 206980 12928 206986 12940
rect 314838 12928 314844 12940
rect 314896 12928 314902 12980
rect 211062 12860 211068 12912
rect 211120 12900 211126 12912
rect 316218 12900 316224 12912
rect 211120 12872 316224 12900
rect 211120 12860 211126 12872
rect 316218 12860 316224 12872
rect 316276 12860 316282 12912
rect 213822 12792 213828 12844
rect 213880 12832 213886 12844
rect 317598 12832 317604 12844
rect 213880 12804 317604 12832
rect 213880 12792 213886 12804
rect 317598 12792 317604 12804
rect 317656 12792 317662 12844
rect 217962 12724 217968 12776
rect 218020 12764 218026 12776
rect 318978 12764 318984 12776
rect 218020 12736 318984 12764
rect 218020 12724 218026 12736
rect 318978 12724 318984 12736
rect 319036 12724 319042 12776
rect 220722 12656 220728 12708
rect 220780 12696 220786 12708
rect 320266 12696 320272 12708
rect 220780 12668 320272 12696
rect 220780 12656 220786 12668
rect 320266 12656 320272 12668
rect 320324 12656 320330 12708
rect 224862 12588 224868 12640
rect 224920 12628 224926 12640
rect 321738 12628 321744 12640
rect 224920 12600 321744 12628
rect 224920 12588 224926 12600
rect 321738 12588 321744 12600
rect 321796 12588 321802 12640
rect 229002 12520 229008 12572
rect 229060 12560 229066 12572
rect 323118 12560 323124 12572
rect 229060 12532 323124 12560
rect 229060 12520 229066 12532
rect 323118 12520 323124 12532
rect 323176 12520 323182 12572
rect 295610 12492 295616 12504
rect 295571 12464 295616 12492
rect 295610 12452 295616 12464
rect 295668 12452 295674 12504
rect 173802 12384 173808 12436
rect 173860 12424 173866 12436
rect 300946 12424 300952 12436
rect 173860 12396 300952 12424
rect 173860 12384 173866 12396
rect 300946 12384 300952 12396
rect 301004 12384 301010 12436
rect 392118 12384 392124 12436
rect 392176 12424 392182 12436
rect 393038 12424 393044 12436
rect 392176 12396 393044 12424
rect 392176 12384 392182 12396
rect 393038 12384 393044 12396
rect 393096 12384 393102 12436
rect 426434 12384 426440 12436
rect 426492 12424 426498 12436
rect 427538 12424 427544 12436
rect 426492 12396 427544 12424
rect 426492 12384 426498 12396
rect 427538 12384 427544 12396
rect 427596 12384 427602 12436
rect 169662 12316 169668 12368
rect 169720 12356 169726 12368
rect 299566 12356 299572 12368
rect 169720 12328 299572 12356
rect 169720 12316 169726 12328
rect 299566 12316 299572 12328
rect 299624 12316 299630 12368
rect 166902 12248 166908 12300
rect 166960 12288 166966 12300
rect 298186 12288 298192 12300
rect 166960 12260 298192 12288
rect 166960 12248 166966 12260
rect 298186 12248 298192 12260
rect 298244 12248 298250 12300
rect 162762 12180 162768 12232
rect 162820 12220 162826 12232
rect 295613 12223 295671 12229
rect 295613 12220 295625 12223
rect 162820 12192 295625 12220
rect 162820 12180 162826 12192
rect 295613 12189 295625 12192
rect 295659 12189 295671 12223
rect 295613 12183 295671 12189
rect 151722 12112 151728 12164
rect 151780 12152 151786 12164
rect 291562 12152 291568 12164
rect 151780 12124 291568 12152
rect 151780 12112 151786 12124
rect 291562 12112 291568 12124
rect 291620 12112 291626 12164
rect 148962 12044 148968 12096
rect 149020 12084 149026 12096
rect 290274 12084 290280 12096
rect 149020 12056 290280 12084
rect 149020 12044 149026 12056
rect 290274 12044 290280 12056
rect 290332 12044 290338 12096
rect 144822 11976 144828 12028
rect 144880 12016 144886 12028
rect 288802 12016 288808 12028
rect 144880 11988 288808 12016
rect 144880 11976 144886 11988
rect 288802 11976 288808 11988
rect 288860 11976 288866 12028
rect 142062 11908 142068 11960
rect 142120 11948 142126 11960
rect 287330 11948 287336 11960
rect 142120 11920 287336 11948
rect 142120 11908 142126 11920
rect 287330 11908 287336 11920
rect 287388 11908 287394 11960
rect 128262 11840 128268 11892
rect 128320 11880 128326 11892
rect 281534 11880 281540 11892
rect 128320 11852 281540 11880
rect 128320 11840 128326 11852
rect 281534 11840 281540 11852
rect 281592 11840 281598 11892
rect 126882 11772 126888 11824
rect 126940 11812 126946 11824
rect 281626 11812 281632 11824
rect 126940 11784 281632 11812
rect 126940 11772 126946 11784
rect 281626 11772 281632 11784
rect 281684 11772 281690 11824
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 238938 11744 238944 11756
rect 23440 11716 238944 11744
rect 23440 11704 23446 11716
rect 238938 11704 238944 11716
rect 238996 11704 239002 11756
rect 176470 11636 176476 11688
rect 176528 11676 176534 11688
rect 302326 11676 302332 11688
rect 176528 11648 302332 11676
rect 176528 11636 176534 11648
rect 302326 11636 302332 11648
rect 302384 11636 302390 11688
rect 180702 11568 180708 11620
rect 180760 11608 180766 11620
rect 303706 11608 303712 11620
rect 180760 11580 303712 11608
rect 180760 11568 180766 11580
rect 303706 11568 303712 11580
rect 303764 11568 303770 11620
rect 184842 11500 184848 11552
rect 184900 11540 184906 11552
rect 305086 11540 305092 11552
rect 184900 11512 305092 11540
rect 184900 11500 184906 11512
rect 305086 11500 305092 11512
rect 305144 11500 305150 11552
rect 187602 11432 187608 11484
rect 187660 11472 187666 11484
rect 306466 11472 306472 11484
rect 187660 11444 306472 11472
rect 187660 11432 187666 11444
rect 306466 11432 306472 11444
rect 306524 11432 306530 11484
rect 191742 11364 191748 11416
rect 191800 11404 191806 11416
rect 308030 11404 308036 11416
rect 191800 11376 308036 11404
rect 191800 11364 191806 11376
rect 308030 11364 308036 11376
rect 308088 11364 308094 11416
rect 194502 11296 194508 11348
rect 194560 11336 194566 11348
rect 309410 11336 309416 11348
rect 194560 11308 309416 11336
rect 194560 11296 194566 11308
rect 309410 11296 309416 11308
rect 309468 11296 309474 11348
rect 198642 11228 198648 11280
rect 198700 11268 198706 11280
rect 307570 11268 307576 11280
rect 198700 11240 307576 11268
rect 198700 11228 198706 11240
rect 307570 11228 307576 11240
rect 307628 11228 307634 11280
rect 337102 11200 337108 11212
rect 337063 11172 337108 11200
rect 337102 11160 337108 11172
rect 337160 11160 337166 11212
rect 113082 10956 113088 11008
rect 113140 10996 113146 11008
rect 276014 10996 276020 11008
rect 113140 10968 276020 10996
rect 113140 10956 113146 10968
rect 276014 10956 276020 10968
rect 276072 10956 276078 11008
rect 108942 10888 108948 10940
rect 109000 10928 109006 10940
rect 273441 10931 273499 10937
rect 273441 10928 273453 10931
rect 109000 10900 273453 10928
rect 109000 10888 109006 10900
rect 273441 10897 273453 10900
rect 273487 10897 273499 10931
rect 273441 10891 273499 10897
rect 106182 10820 106188 10872
rect 106240 10860 106246 10872
rect 271874 10860 271880 10872
rect 106240 10832 271880 10860
rect 106240 10820 106246 10832
rect 271874 10820 271880 10832
rect 271932 10820 271938 10872
rect 102042 10752 102048 10804
rect 102100 10792 102106 10804
rect 270494 10792 270500 10804
rect 102100 10764 270500 10792
rect 102100 10752 102106 10764
rect 270494 10752 270500 10764
rect 270552 10752 270558 10804
rect 99190 10684 99196 10736
rect 99248 10724 99254 10736
rect 269298 10724 269304 10736
rect 99248 10696 269304 10724
rect 99248 10684 99254 10696
rect 269298 10684 269304 10696
rect 269356 10684 269362 10736
rect 95142 10616 95148 10668
rect 95200 10656 95206 10668
rect 267737 10659 267795 10665
rect 267737 10656 267749 10659
rect 95200 10628 267749 10656
rect 95200 10616 95206 10628
rect 267737 10625 267749 10628
rect 267783 10625 267795 10659
rect 267737 10619 267795 10625
rect 91002 10548 91008 10600
rect 91060 10588 91066 10600
rect 266722 10588 266728 10600
rect 91060 10560 266728 10588
rect 91060 10548 91066 10560
rect 266722 10548 266728 10560
rect 266780 10548 266786 10600
rect 64782 10480 64788 10532
rect 64840 10520 64846 10532
rect 255590 10520 255596 10532
rect 64840 10492 255596 10520
rect 64840 10480 64846 10492
rect 255590 10480 255596 10492
rect 255648 10480 255654 10532
rect 60642 10412 60648 10464
rect 60700 10452 60706 10464
rect 254026 10452 254032 10464
rect 60700 10424 254032 10452
rect 60700 10412 60706 10424
rect 254026 10412 254032 10424
rect 254084 10412 254090 10464
rect 56502 10344 56508 10396
rect 56560 10384 56566 10396
rect 252646 10384 252652 10396
rect 56560 10356 252652 10384
rect 56560 10344 56566 10356
rect 252646 10344 252652 10356
rect 252704 10344 252710 10396
rect 53742 10276 53748 10328
rect 53800 10316 53806 10328
rect 251266 10316 251272 10328
rect 53800 10288 251272 10316
rect 53800 10276 53806 10288
rect 251266 10276 251272 10288
rect 251324 10276 251330 10328
rect 117130 10208 117136 10260
rect 117188 10248 117194 10260
rect 277578 10248 277584 10260
rect 117188 10220 277584 10248
rect 117188 10208 117194 10220
rect 277578 10208 277584 10220
rect 277636 10208 277642 10260
rect 119982 10140 119988 10192
rect 120040 10180 120046 10192
rect 278958 10180 278964 10192
rect 120040 10152 278964 10180
rect 120040 10140 120046 10152
rect 278958 10140 278964 10152
rect 279016 10140 279022 10192
rect 124122 10072 124128 10124
rect 124180 10112 124186 10124
rect 280338 10112 280344 10124
rect 124180 10084 280344 10112
rect 124180 10072 124186 10084
rect 280338 10072 280344 10084
rect 280396 10072 280402 10124
rect 366910 10112 366916 10124
rect 366871 10084 366916 10112
rect 366910 10072 366916 10084
rect 366968 10072 366974 10124
rect 143442 10004 143448 10056
rect 143500 10044 143506 10056
rect 288526 10044 288532 10056
rect 143500 10016 288532 10044
rect 143500 10004 143506 10016
rect 288526 10004 288532 10016
rect 288584 10004 288590 10056
rect 147582 9936 147588 9988
rect 147640 9976 147646 9988
rect 289814 9976 289820 9988
rect 147640 9948 289820 9976
rect 147640 9936 147646 9948
rect 289814 9936 289820 9948
rect 289872 9936 289878 9988
rect 151630 9868 151636 9920
rect 151688 9908 151694 9920
rect 291286 9908 291292 9920
rect 151688 9880 291292 9908
rect 151688 9868 151694 9880
rect 291286 9868 291292 9880
rect 291344 9868 291350 9920
rect 154482 9800 154488 9852
rect 154540 9840 154546 9852
rect 292850 9840 292856 9852
rect 154540 9812 292856 9840
rect 154540 9800 154546 9812
rect 292850 9800 292856 9812
rect 292908 9800 292914 9852
rect 158622 9732 158628 9784
rect 158680 9772 158686 9784
rect 294046 9772 294052 9784
rect 158680 9744 294052 9772
rect 158680 9732 158686 9744
rect 294046 9732 294052 9744
rect 294104 9732 294110 9784
rect 161382 9664 161388 9716
rect 161440 9704 161446 9716
rect 295426 9704 295432 9716
rect 161440 9676 295432 9704
rect 161440 9664 161446 9676
rect 295426 9664 295432 9676
rect 295484 9664 295490 9716
rect 306650 9664 306656 9716
rect 306708 9704 306714 9716
rect 306926 9704 306932 9716
rect 306708 9676 306932 9704
rect 306708 9664 306714 9676
rect 306926 9664 306932 9676
rect 306984 9664 306990 9716
rect 341242 9704 341248 9716
rect 341203 9676 341248 9704
rect 341242 9664 341248 9676
rect 341300 9664 341306 9716
rect 358538 9704 358544 9716
rect 358499 9676 358544 9704
rect 358538 9664 358544 9676
rect 358596 9664 358602 9716
rect 421193 9707 421251 9713
rect 421193 9673 421205 9707
rect 421239 9704 421251 9707
rect 421466 9704 421472 9716
rect 421239 9676 421472 9704
rect 421239 9673 421251 9676
rect 421193 9667 421251 9673
rect 421466 9664 421472 9676
rect 421524 9664 421530 9716
rect 203886 9596 203892 9648
rect 203944 9636 203950 9648
rect 313366 9636 313372 9648
rect 203944 9608 313372 9636
rect 203944 9596 203950 9608
rect 313366 9596 313372 9608
rect 313424 9596 313430 9648
rect 330202 9636 330208 9648
rect 330163 9608 330208 9636
rect 330202 9596 330208 9608
rect 330260 9596 330266 9648
rect 336918 9636 336924 9648
rect 336879 9608 336924 9636
rect 336918 9596 336924 9608
rect 336976 9596 336982 9648
rect 389453 9639 389511 9645
rect 389453 9605 389465 9639
rect 389499 9636 389511 9639
rect 389542 9636 389548 9648
rect 389499 9608 389548 9636
rect 389499 9605 389511 9608
rect 389453 9599 389511 9605
rect 389542 9596 389548 9608
rect 389600 9596 389606 9648
rect 200390 9528 200396 9580
rect 200448 9568 200454 9580
rect 311986 9568 311992 9580
rect 200448 9540 311992 9568
rect 200448 9528 200454 9540
rect 311986 9528 311992 9540
rect 312044 9528 312050 9580
rect 196802 9460 196808 9512
rect 196860 9500 196866 9512
rect 310606 9500 310612 9512
rect 196860 9472 310612 9500
rect 196860 9460 196866 9472
rect 310606 9460 310612 9472
rect 310664 9460 310670 9512
rect 193214 9392 193220 9444
rect 193272 9432 193278 9444
rect 309226 9432 309232 9444
rect 193272 9404 309232 9432
rect 193272 9392 193278 9404
rect 309226 9392 309232 9404
rect 309284 9392 309290 9444
rect 139670 9324 139676 9376
rect 139728 9364 139734 9376
rect 287146 9364 287152 9376
rect 139728 9336 287152 9364
rect 139728 9324 139734 9336
rect 287146 9324 287152 9336
rect 287204 9324 287210 9376
rect 136082 9256 136088 9308
rect 136140 9296 136146 9308
rect 285858 9296 285864 9308
rect 136140 9268 285864 9296
rect 136140 9256 136146 9268
rect 285858 9256 285864 9268
rect 285916 9256 285922 9308
rect 49326 9188 49332 9240
rect 49384 9228 49390 9240
rect 249886 9228 249892 9240
rect 49384 9200 249892 9228
rect 49384 9188 49390 9200
rect 249886 9188 249892 9200
rect 249944 9188 249950 9240
rect 253842 9188 253848 9240
rect 253900 9228 253906 9240
rect 334158 9228 334164 9240
rect 253900 9200 334164 9228
rect 253900 9188 253906 9200
rect 334158 9188 334164 9200
rect 334216 9188 334222 9240
rect 44542 9120 44548 9172
rect 44600 9160 44606 9172
rect 247218 9160 247224 9172
rect 44600 9132 247224 9160
rect 44600 9120 44606 9132
rect 247218 9120 247224 9132
rect 247276 9120 247282 9172
rect 250346 9120 250352 9172
rect 250404 9160 250410 9172
rect 332778 9160 332784 9172
rect 250404 9132 332784 9160
rect 250404 9120 250410 9132
rect 332778 9120 332784 9132
rect 332836 9120 332842 9172
rect 27890 9052 27896 9104
rect 27948 9092 27954 9104
rect 233878 9092 233884 9104
rect 27948 9064 233884 9092
rect 27948 9052 27954 9064
rect 233878 9052 233884 9064
rect 233936 9052 233942 9104
rect 243170 9052 243176 9104
rect 243228 9092 243234 9104
rect 330018 9092 330024 9104
rect 243228 9064 330024 9092
rect 243228 9052 243234 9064
rect 330018 9052 330024 9064
rect 330076 9052 330082 9104
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 236178 9024 236184 9036
rect 18380 8996 236184 9024
rect 18380 8984 18386 8996
rect 236178 8984 236184 8996
rect 236236 8984 236242 9036
rect 239582 8984 239588 9036
rect 239640 9024 239646 9036
rect 328638 9024 328644 9036
rect 239640 8996 328644 9024
rect 239640 8984 239646 8996
rect 328638 8984 328644 8996
rect 328696 8984 328702 9036
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 234798 8956 234804 8968
rect 13688 8928 234804 8956
rect 13688 8916 13694 8928
rect 234798 8916 234804 8928
rect 234856 8916 234862 8968
rect 235994 8916 236000 8968
rect 236052 8956 236058 8968
rect 325970 8956 325976 8968
rect 236052 8928 325976 8956
rect 236052 8916 236058 8928
rect 325970 8916 325976 8928
rect 326028 8916 326034 8968
rect 207474 8848 207480 8900
rect 207532 8888 207538 8900
rect 314930 8888 314936 8900
rect 207532 8860 314936 8888
rect 207532 8848 207538 8860
rect 314930 8848 314936 8860
rect 314988 8848 314994 8900
rect 210970 8780 210976 8832
rect 211028 8820 211034 8832
rect 316126 8820 316132 8832
rect 211028 8792 316132 8820
rect 211028 8780 211034 8792
rect 316126 8780 316132 8792
rect 316184 8780 316190 8832
rect 214650 8712 214656 8764
rect 214708 8752 214714 8764
rect 317506 8752 317512 8764
rect 214708 8724 317512 8752
rect 214708 8712 214714 8724
rect 317506 8712 317512 8724
rect 317564 8712 317570 8764
rect 218146 8644 218152 8696
rect 218204 8684 218210 8696
rect 318886 8684 318892 8696
rect 218204 8656 318892 8684
rect 218204 8644 218210 8656
rect 318886 8644 318892 8656
rect 318944 8644 318950 8696
rect 221734 8576 221740 8628
rect 221792 8616 221798 8628
rect 320174 8616 320180 8628
rect 221792 8588 320180 8616
rect 221792 8576 221798 8588
rect 320174 8576 320180 8588
rect 320232 8576 320238 8628
rect 225322 8508 225328 8560
rect 225380 8548 225386 8560
rect 321646 8548 321652 8560
rect 225380 8520 321652 8548
rect 225380 8508 225386 8520
rect 321646 8508 321652 8520
rect 321704 8508 321710 8560
rect 228910 8440 228916 8492
rect 228968 8480 228974 8492
rect 323302 8480 323308 8492
rect 228968 8452 323308 8480
rect 228968 8440 228974 8452
rect 323302 8440 323308 8452
rect 323360 8440 323366 8492
rect 232498 8372 232504 8424
rect 232556 8412 232562 8424
rect 324590 8412 324596 8424
rect 232556 8384 324596 8412
rect 232556 8372 232562 8384
rect 324590 8372 324596 8384
rect 324648 8372 324654 8424
rect 234890 8304 234896 8356
rect 234948 8344 234954 8356
rect 235074 8344 235080 8356
rect 234948 8316 235080 8344
rect 234948 8304 234954 8316
rect 235074 8304 235080 8316
rect 235132 8304 235138 8356
rect 246758 8304 246764 8356
rect 246816 8344 246822 8356
rect 331398 8344 331404 8356
rect 246816 8316 331404 8344
rect 246816 8304 246822 8316
rect 331398 8304 331404 8316
rect 331456 8304 331462 8356
rect 362218 8344 362224 8356
rect 362179 8316 362224 8344
rect 362218 8304 362224 8316
rect 362276 8304 362282 8356
rect 376754 8344 376760 8356
rect 376715 8316 376760 8344
rect 376754 8304 376760 8316
rect 376812 8304 376818 8356
rect 468754 8304 468760 8356
rect 468812 8344 468818 8356
rect 469030 8344 469036 8356
rect 468812 8316 469036 8344
rect 468812 8304 468818 8316
rect 469030 8304 469036 8316
rect 469088 8304 469094 8356
rect 87322 8236 87328 8288
rect 87380 8276 87386 8288
rect 265158 8276 265164 8288
rect 87380 8248 265164 8276
rect 87380 8236 87386 8248
rect 265158 8236 265164 8248
rect 265216 8236 265222 8288
rect 270494 8236 270500 8288
rect 270552 8276 270558 8288
rect 340966 8276 340972 8288
rect 270552 8248 340972 8276
rect 270552 8236 270558 8248
rect 340966 8236 340972 8248
rect 341024 8236 341030 8288
rect 445478 8236 445484 8288
rect 445536 8276 445542 8288
rect 523862 8276 523868 8288
rect 445536 8248 523868 8276
rect 445536 8236 445542 8248
rect 523862 8236 523868 8248
rect 523920 8236 523926 8288
rect 83826 8168 83832 8220
rect 83884 8208 83890 8220
rect 263870 8208 263876 8220
rect 83884 8180 263876 8208
rect 83884 8168 83890 8180
rect 263870 8168 263876 8180
rect 263928 8168 263934 8220
rect 266998 8168 267004 8220
rect 267056 8208 267062 8220
rect 339586 8208 339592 8220
rect 267056 8180 339592 8208
rect 267056 8168 267062 8180
rect 339586 8168 339592 8180
rect 339644 8168 339650 8220
rect 446950 8168 446956 8220
rect 447008 8208 447014 8220
rect 527450 8208 527456 8220
rect 447008 8180 527456 8208
rect 447008 8168 447014 8180
rect 527450 8168 527456 8180
rect 527508 8168 527514 8220
rect 80238 8100 80244 8152
rect 80296 8140 80302 8152
rect 262398 8140 262404 8152
rect 80296 8112 262404 8140
rect 80296 8100 80302 8112
rect 262398 8100 262404 8112
rect 262456 8100 262462 8152
rect 263410 8100 263416 8152
rect 263468 8140 263474 8152
rect 338298 8140 338304 8152
rect 263468 8112 338304 8140
rect 263468 8100 263474 8112
rect 338298 8100 338304 8112
rect 338356 8100 338362 8152
rect 448238 8100 448244 8152
rect 448296 8140 448302 8152
rect 531038 8140 531044 8152
rect 448296 8112 531044 8140
rect 448296 8100 448302 8112
rect 531038 8100 531044 8112
rect 531096 8100 531102 8152
rect 40954 8032 40960 8084
rect 41012 8072 41018 8084
rect 245930 8072 245936 8084
rect 41012 8044 245936 8072
rect 41012 8032 41018 8044
rect 245930 8032 245936 8044
rect 245988 8032 245994 8084
rect 259822 8032 259828 8084
rect 259880 8072 259886 8084
rect 336921 8075 336979 8081
rect 336921 8072 336933 8075
rect 259880 8044 336933 8072
rect 259880 8032 259886 8044
rect 336921 8041 336933 8044
rect 336967 8041 336979 8075
rect 336921 8035 336979 8041
rect 450998 8032 451004 8084
rect 451056 8072 451062 8084
rect 534534 8072 534540 8084
rect 451056 8044 534540 8072
rect 451056 8032 451062 8044
rect 534534 8032 534540 8044
rect 534592 8032 534598 8084
rect 37366 7964 37372 8016
rect 37424 8004 37430 8016
rect 244182 8004 244188 8016
rect 37424 7976 244188 8004
rect 37424 7964 37430 7976
rect 244182 7964 244188 7976
rect 244240 7964 244246 8016
rect 256234 7964 256240 8016
rect 256292 8004 256298 8016
rect 334066 8004 334072 8016
rect 256292 7976 334072 8004
rect 256292 7964 256298 7976
rect 334066 7964 334072 7976
rect 334124 7964 334130 8016
rect 452470 7964 452476 8016
rect 452528 8004 452534 8016
rect 538122 8004 538128 8016
rect 452528 7976 538128 8004
rect 452528 7964 452534 7976
rect 538122 7964 538128 7976
rect 538180 7964 538186 8016
rect 33870 7896 33876 7948
rect 33928 7936 33934 7948
rect 242986 7936 242992 7948
rect 33928 7908 242992 7936
rect 33928 7896 33934 7908
rect 242986 7896 242992 7908
rect 243044 7896 243050 7948
rect 252646 7896 252652 7948
rect 252704 7936 252710 7948
rect 332686 7936 332692 7948
rect 252704 7908 332692 7936
rect 252704 7896 252710 7908
rect 332686 7896 332692 7908
rect 332744 7896 332750 7948
rect 453758 7896 453764 7948
rect 453816 7936 453822 7948
rect 541710 7936 541716 7948
rect 453816 7908 541716 7936
rect 453816 7896 453822 7908
rect 541710 7896 541716 7908
rect 541768 7896 541774 7948
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 241790 7868 241796 7880
rect 30340 7840 241796 7868
rect 30340 7828 30346 7840
rect 241790 7828 241796 7840
rect 241848 7828 241854 7880
rect 249150 7828 249156 7880
rect 249208 7868 249214 7880
rect 331306 7868 331312 7880
rect 249208 7840 331312 7868
rect 249208 7828 249214 7840
rect 331306 7828 331312 7840
rect 331364 7828 331370 7880
rect 455230 7828 455236 7880
rect 455288 7868 455294 7880
rect 545298 7868 545304 7880
rect 455288 7840 545304 7868
rect 455288 7828 455294 7840
rect 545298 7828 545304 7840
rect 545356 7828 545362 7880
rect 26694 7760 26700 7812
rect 26752 7800 26758 7812
rect 240410 7800 240416 7812
rect 26752 7772 240416 7800
rect 26752 7760 26758 7772
rect 240410 7760 240416 7772
rect 240468 7760 240474 7812
rect 245562 7760 245568 7812
rect 245620 7800 245626 7812
rect 330205 7803 330263 7809
rect 330205 7800 330217 7803
rect 245620 7772 330217 7800
rect 245620 7760 245626 7772
rect 330205 7769 330217 7772
rect 330251 7769 330263 7803
rect 330205 7763 330263 7769
rect 456610 7760 456616 7812
rect 456668 7800 456674 7812
rect 548886 7800 548892 7812
rect 456668 7772 548892 7800
rect 456668 7760 456674 7772
rect 548886 7760 548892 7772
rect 548944 7760 548950 7812
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 238846 7732 238852 7744
rect 21968 7704 238852 7732
rect 21968 7692 21974 7704
rect 238846 7692 238852 7704
rect 238904 7692 238910 7744
rect 241974 7692 241980 7744
rect 242032 7732 242038 7744
rect 328546 7732 328552 7744
rect 242032 7704 328552 7732
rect 242032 7692 242038 7704
rect 328546 7692 328552 7704
rect 328604 7692 328610 7744
rect 457990 7692 457996 7744
rect 458048 7732 458054 7744
rect 552382 7732 552388 7744
rect 458048 7704 552388 7732
rect 458048 7692 458054 7704
rect 552382 7692 552388 7704
rect 552440 7692 552446 7744
rect 8846 7624 8852 7676
rect 8904 7664 8910 7676
rect 227533 7667 227591 7673
rect 227533 7664 227545 7667
rect 8904 7636 227545 7664
rect 8904 7624 8910 7636
rect 227533 7633 227545 7636
rect 227579 7633 227591 7667
rect 230658 7664 230664 7676
rect 227533 7627 227591 7633
rect 227640 7636 230664 7664
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 227640 7596 227668 7636
rect 230658 7624 230664 7636
rect 230716 7624 230722 7676
rect 234798 7624 234804 7676
rect 234856 7664 234862 7676
rect 325786 7664 325792 7676
rect 234856 7636 325792 7664
rect 234856 7624 234862 7636
rect 325786 7624 325792 7636
rect 325844 7624 325850 7676
rect 459370 7624 459376 7676
rect 459428 7664 459434 7676
rect 555970 7664 555976 7676
rect 459428 7636 555976 7664
rect 459428 7624 459434 7636
rect 555970 7624 555976 7636
rect 556028 7624 556034 7676
rect 4120 7568 227668 7596
rect 4120 7556 4126 7568
rect 227714 7556 227720 7608
rect 227772 7596 227778 7608
rect 229002 7596 229008 7608
rect 227772 7568 229008 7596
rect 227772 7556 227778 7568
rect 229002 7556 229008 7568
rect 229060 7556 229066 7608
rect 231302 7556 231308 7608
rect 231360 7596 231366 7608
rect 324406 7596 324412 7608
rect 231360 7568 324412 7596
rect 231360 7556 231366 7568
rect 324406 7556 324412 7568
rect 324464 7556 324470 7608
rect 460750 7556 460756 7608
rect 460808 7596 460814 7608
rect 559558 7596 559564 7608
rect 460808 7568 559564 7596
rect 460808 7556 460814 7568
rect 559558 7556 559564 7568
rect 559616 7556 559622 7608
rect 134886 7488 134892 7540
rect 134944 7528 134950 7540
rect 284570 7528 284576 7540
rect 134944 7500 284576 7528
rect 134944 7488 134950 7500
rect 284570 7488 284576 7500
rect 284628 7488 284634 7540
rect 444190 7488 444196 7540
rect 444248 7528 444254 7540
rect 520274 7528 520280 7540
rect 444248 7500 520280 7528
rect 444248 7488 444254 7500
rect 520274 7488 520280 7500
rect 520332 7488 520338 7540
rect 138474 7420 138480 7472
rect 138532 7460 138538 7472
rect 285950 7460 285956 7472
rect 138532 7432 285956 7460
rect 138532 7420 138538 7432
rect 285950 7420 285956 7432
rect 286008 7420 286014 7472
rect 442810 7420 442816 7472
rect 442868 7460 442874 7472
rect 516778 7460 516784 7472
rect 442868 7432 516784 7460
rect 442868 7420 442874 7432
rect 516778 7420 516784 7432
rect 516836 7420 516842 7472
rect 141970 7352 141976 7404
rect 142028 7392 142034 7404
rect 287054 7392 287060 7404
rect 142028 7364 287060 7392
rect 142028 7352 142034 7364
rect 287054 7352 287060 7364
rect 287112 7352 287118 7404
rect 441430 7352 441436 7404
rect 441488 7392 441494 7404
rect 513190 7392 513196 7404
rect 441488 7364 513196 7392
rect 441488 7352 441494 7364
rect 513190 7352 513196 7364
rect 513248 7352 513254 7404
rect 145650 7284 145656 7336
rect 145708 7324 145714 7336
rect 288434 7324 288440 7336
rect 145708 7296 288440 7324
rect 145708 7284 145714 7296
rect 288434 7284 288440 7296
rect 288492 7284 288498 7336
rect 440050 7284 440056 7336
rect 440108 7324 440114 7336
rect 509602 7324 509608 7336
rect 440108 7296 509608 7324
rect 440108 7284 440114 7296
rect 509602 7284 509608 7296
rect 509660 7284 509666 7336
rect 149238 7216 149244 7268
rect 149296 7256 149302 7268
rect 291194 7256 291200 7268
rect 149296 7228 291200 7256
rect 149296 7216 149302 7228
rect 291194 7216 291200 7228
rect 291252 7216 291258 7268
rect 152734 7148 152740 7200
rect 152792 7188 152798 7200
rect 292574 7188 292580 7200
rect 152792 7160 292580 7188
rect 152792 7148 152798 7160
rect 292574 7148 292580 7160
rect 292632 7148 292638 7200
rect 156322 7080 156328 7132
rect 156380 7120 156386 7132
rect 293954 7120 293960 7132
rect 156380 7092 293960 7120
rect 156380 7080 156386 7092
rect 293954 7080 293960 7092
rect 294012 7080 294018 7132
rect 159910 7012 159916 7064
rect 159968 7052 159974 7064
rect 295334 7052 295340 7064
rect 159968 7024 295340 7052
rect 159968 7012 159974 7024
rect 295334 7012 295340 7024
rect 295392 7012 295398 7064
rect 227533 6987 227591 6993
rect 227533 6953 227545 6987
rect 227579 6984 227591 6987
rect 233418 6984 233424 6996
rect 227579 6956 233424 6984
rect 227579 6953 227591 6956
rect 227533 6947 227591 6953
rect 233418 6944 233424 6956
rect 233476 6944 233482 6996
rect 238386 6944 238392 6996
rect 238444 6984 238450 6996
rect 327258 6984 327264 6996
rect 238444 6956 327264 6984
rect 238444 6944 238450 6956
rect 327258 6944 327264 6956
rect 327316 6944 327322 6996
rect 516686 6876 516692 6928
rect 516744 6916 516750 6928
rect 516870 6916 516876 6928
rect 516744 6888 516876 6916
rect 516744 6876 516750 6888
rect 516870 6876 516876 6888
rect 516928 6876 516934 6928
rect 170582 6808 170588 6860
rect 170640 6848 170646 6860
rect 299474 6848 299480 6860
rect 170640 6820 299480 6848
rect 170640 6808 170646 6820
rect 299474 6808 299480 6820
rect 299532 6808 299538 6860
rect 433242 6808 433248 6860
rect 433300 6848 433306 6860
rect 491754 6848 491760 6860
rect 433300 6820 491760 6848
rect 433300 6808 433306 6820
rect 491754 6808 491760 6820
rect 491812 6808 491818 6860
rect 167086 6740 167092 6792
rect 167144 6780 167150 6792
rect 298370 6780 298376 6792
rect 167144 6752 298376 6780
rect 167144 6740 167150 6752
rect 298370 6740 298376 6752
rect 298428 6740 298434 6792
rect 431770 6740 431776 6792
rect 431828 6780 431834 6792
rect 490558 6780 490564 6792
rect 431828 6752 490564 6780
rect 431828 6740 431834 6752
rect 490558 6740 490564 6752
rect 490616 6740 490622 6792
rect 163498 6672 163504 6724
rect 163556 6712 163562 6724
rect 296714 6712 296720 6724
rect 163556 6684 296720 6712
rect 163556 6672 163562 6684
rect 296714 6672 296720 6684
rect 296772 6672 296778 6724
rect 297358 6672 297364 6724
rect 297416 6712 297422 6724
rect 336826 6712 336832 6724
rect 297416 6684 336832 6712
rect 297416 6672 297422 6684
rect 336826 6672 336832 6684
rect 336884 6672 336890 6724
rect 434622 6672 434628 6724
rect 434680 6712 434686 6724
rect 495342 6712 495348 6724
rect 434680 6684 495348 6712
rect 434680 6672 434686 6684
rect 495342 6672 495348 6684
rect 495400 6672 495406 6724
rect 131390 6604 131396 6656
rect 131448 6644 131454 6656
rect 283006 6644 283012 6656
rect 131448 6616 283012 6644
rect 131448 6604 131454 6616
rect 283006 6604 283012 6616
rect 283064 6604 283070 6656
rect 298094 6604 298100 6656
rect 298152 6644 298158 6656
rect 338390 6644 338396 6656
rect 298152 6616 338396 6644
rect 298152 6604 298158 6616
rect 338390 6604 338396 6616
rect 338448 6604 338454 6656
rect 433150 6604 433156 6656
rect 433208 6644 433214 6656
rect 494146 6644 494152 6656
rect 433208 6616 494152 6644
rect 433208 6604 433214 6616
rect 494146 6604 494152 6616
rect 494204 6604 494210 6656
rect 76650 6536 76656 6588
rect 76708 6576 76714 6588
rect 261018 6576 261024 6588
rect 76708 6548 261024 6576
rect 76708 6536 76714 6548
rect 261018 6536 261024 6548
rect 261076 6536 261082 6588
rect 295886 6536 295892 6588
rect 295944 6576 295950 6588
rect 335446 6576 335452 6588
rect 295944 6548 335452 6576
rect 295944 6536 295950 6548
rect 335446 6536 335452 6548
rect 335504 6536 335510 6588
rect 435910 6536 435916 6588
rect 435968 6576 435974 6588
rect 497734 6576 497740 6588
rect 435968 6548 497740 6576
rect 435968 6536 435974 6548
rect 497734 6536 497740 6548
rect 497792 6536 497798 6588
rect 73062 6468 73068 6520
rect 73120 6508 73126 6520
rect 259454 6508 259460 6520
rect 73120 6480 259460 6508
rect 73120 6468 73126 6480
rect 259454 6468 259460 6480
rect 259512 6468 259518 6520
rect 289814 6468 289820 6520
rect 289872 6508 289878 6520
rect 339678 6508 339684 6520
rect 289872 6480 339684 6508
rect 289872 6468 289878 6480
rect 339678 6468 339684 6480
rect 339736 6468 339742 6520
rect 436002 6468 436008 6520
rect 436060 6508 436066 6520
rect 498930 6508 498936 6520
rect 436060 6480 498936 6508
rect 436060 6468 436066 6480
rect 498930 6468 498936 6480
rect 498988 6468 498994 6520
rect 69474 6400 69480 6452
rect 69532 6440 69538 6452
rect 258258 6440 258264 6452
rect 69532 6412 258264 6440
rect 69532 6400 69538 6412
rect 258258 6400 258264 6412
rect 258316 6400 258322 6452
rect 288434 6400 288440 6452
rect 288492 6440 288498 6452
rect 341242 6440 341248 6452
rect 288492 6412 341248 6440
rect 288492 6400 288498 6412
rect 341242 6400 341248 6412
rect 341300 6400 341306 6452
rect 437290 6400 437296 6452
rect 437348 6440 437354 6452
rect 501230 6440 501236 6452
rect 437348 6412 501236 6440
rect 437348 6400 437354 6412
rect 501230 6400 501236 6412
rect 501288 6400 501294 6452
rect 65978 6332 65984 6384
rect 66036 6372 66042 6384
rect 256786 6372 256792 6384
rect 66036 6344 256792 6372
rect 66036 6332 66042 6344
rect 256786 6332 256792 6344
rect 256844 6332 256850 6384
rect 288526 6332 288532 6384
rect 288584 6372 288590 6384
rect 343634 6372 343640 6384
rect 288584 6344 343640 6372
rect 288584 6332 288590 6344
rect 343634 6332 343640 6344
rect 343692 6332 343698 6384
rect 437382 6332 437388 6384
rect 437440 6372 437446 6384
rect 502426 6372 502432 6384
rect 437440 6344 502432 6372
rect 437440 6332 437446 6344
rect 502426 6332 502432 6344
rect 502484 6332 502490 6384
rect 62390 6264 62396 6316
rect 62448 6304 62454 6316
rect 255498 6304 255504 6316
rect 62448 6276 255504 6304
rect 62448 6264 62454 6276
rect 255498 6264 255504 6276
rect 255556 6264 255562 6316
rect 294322 6264 294328 6316
rect 294380 6304 294386 6316
rect 350626 6304 350632 6316
rect 294380 6276 350632 6304
rect 294380 6264 294386 6276
rect 350626 6264 350632 6276
rect 350684 6264 350690 6316
rect 438762 6264 438768 6316
rect 438820 6304 438826 6316
rect 504818 6304 504824 6316
rect 438820 6276 504824 6304
rect 438820 6264 438826 6276
rect 504818 6264 504824 6276
rect 504876 6264 504882 6316
rect 58802 6196 58808 6248
rect 58860 6236 58866 6248
rect 253934 6236 253940 6248
rect 58860 6208 253940 6236
rect 58860 6196 58866 6208
rect 253934 6196 253940 6208
rect 253992 6196 253998 6248
rect 280062 6196 280068 6248
rect 280120 6236 280126 6248
rect 345198 6236 345204 6248
rect 280120 6208 345204 6236
rect 280120 6196 280126 6208
rect 345198 6196 345204 6208
rect 345256 6196 345262 6248
rect 438670 6196 438676 6248
rect 438728 6236 438734 6248
rect 506014 6236 506020 6248
rect 438728 6208 506020 6236
rect 438728 6196 438734 6208
rect 506014 6196 506020 6208
rect 506072 6196 506078 6248
rect 55214 6128 55220 6180
rect 55272 6168 55278 6180
rect 251358 6168 251364 6180
rect 55272 6140 251364 6168
rect 55272 6128 55278 6140
rect 251358 6128 251364 6140
rect 251416 6128 251422 6180
rect 274082 6128 274088 6180
rect 274140 6168 274146 6180
rect 342346 6168 342352 6180
rect 274140 6140 342352 6168
rect 274140 6128 274146 6140
rect 342346 6128 342352 6140
rect 342404 6128 342410 6180
rect 440142 6128 440148 6180
rect 440200 6168 440206 6180
rect 508406 6168 508412 6180
rect 440200 6140 508412 6168
rect 440200 6128 440206 6140
rect 508406 6128 508412 6140
rect 508464 6128 508470 6180
rect 174170 6060 174176 6112
rect 174228 6100 174234 6112
rect 300854 6100 300860 6112
rect 174228 6072 300860 6100
rect 174228 6060 174234 6072
rect 300854 6060 300860 6072
rect 300912 6060 300918 6112
rect 430390 6060 430396 6112
rect 430448 6100 430454 6112
rect 486970 6100 486976 6112
rect 430448 6072 486976 6100
rect 430448 6060 430454 6072
rect 486970 6060 486976 6072
rect 487028 6060 487034 6112
rect 177758 5992 177764 6044
rect 177816 6032 177822 6044
rect 302234 6032 302240 6044
rect 177816 6004 302240 6032
rect 177816 5992 177822 6004
rect 302234 5992 302240 6004
rect 302292 5992 302298 6044
rect 431862 5992 431868 6044
rect 431920 6032 431926 6044
rect 488166 6032 488172 6044
rect 431920 6004 488172 6032
rect 431920 5992 431926 6004
rect 488166 5992 488172 6004
rect 488224 5992 488230 6044
rect 181346 5924 181352 5976
rect 181404 5964 181410 5976
rect 303614 5964 303620 5976
rect 181404 5936 303620 5964
rect 181404 5924 181410 5936
rect 303614 5924 303620 5936
rect 303672 5924 303678 5976
rect 429102 5924 429108 5976
rect 429160 5964 429166 5976
rect 483474 5964 483480 5976
rect 429160 5936 483480 5964
rect 429160 5924 429166 5936
rect 483474 5924 483480 5936
rect 483532 5924 483538 5976
rect 184842 5856 184848 5908
rect 184900 5896 184906 5908
rect 304994 5896 305000 5908
rect 184900 5868 305000 5896
rect 184900 5856 184906 5868
rect 304994 5856 305000 5868
rect 305052 5856 305058 5908
rect 430482 5856 430488 5908
rect 430540 5896 430546 5908
rect 484578 5896 484584 5908
rect 430540 5868 484584 5896
rect 430540 5856 430546 5868
rect 484578 5856 484584 5868
rect 484636 5856 484642 5908
rect 188430 5788 188436 5840
rect 188488 5828 188494 5840
rect 306650 5828 306656 5840
rect 188488 5800 306656 5828
rect 188488 5788 188494 5800
rect 306650 5788 306656 5800
rect 306708 5788 306714 5840
rect 427722 5788 427728 5840
rect 427780 5828 427786 5840
rect 479886 5828 479892 5840
rect 427780 5800 479892 5828
rect 427780 5788 427786 5800
rect 479886 5788 479892 5800
rect 479944 5788 479950 5840
rect 192018 5720 192024 5772
rect 192076 5760 192082 5772
rect 307754 5760 307760 5772
rect 192076 5732 307760 5760
rect 192076 5720 192082 5732
rect 307754 5720 307760 5732
rect 307812 5720 307818 5772
rect 426342 5720 426348 5772
rect 426400 5760 426406 5772
rect 476298 5760 476304 5772
rect 426400 5732 476304 5760
rect 426400 5720 426406 5732
rect 476298 5720 476304 5732
rect 476356 5720 476362 5772
rect 195606 5652 195612 5704
rect 195664 5692 195670 5704
rect 309134 5692 309140 5704
rect 195664 5664 309140 5692
rect 195664 5652 195670 5664
rect 309134 5652 309140 5664
rect 309192 5652 309198 5704
rect 199194 5584 199200 5636
rect 199252 5624 199258 5636
rect 310514 5624 310520 5636
rect 199252 5596 310520 5624
rect 199252 5584 199258 5596
rect 310514 5584 310520 5596
rect 310572 5584 310578 5636
rect 470594 5584 470600 5636
rect 470652 5624 470658 5636
rect 471517 5627 471575 5633
rect 471517 5624 471529 5627
rect 470652 5596 471529 5624
rect 470652 5584 470658 5596
rect 471517 5593 471529 5596
rect 471563 5593 471575 5627
rect 471517 5587 471575 5593
rect 202690 5516 202696 5568
rect 202748 5556 202754 5568
rect 313274 5556 313280 5568
rect 202748 5528 313280 5556
rect 202748 5516 202754 5528
rect 313274 5516 313280 5528
rect 313332 5516 313338 5568
rect 468938 5516 468944 5568
rect 468996 5556 469002 5568
rect 471425 5559 471483 5565
rect 471425 5556 471437 5559
rect 468996 5528 471437 5556
rect 468996 5516 469002 5528
rect 471425 5525 471437 5528
rect 471471 5525 471483 5559
rect 471425 5519 471483 5525
rect 137278 5448 137284 5500
rect 137336 5488 137342 5500
rect 285674 5488 285680 5500
rect 137336 5460 285680 5488
rect 137336 5448 137342 5460
rect 285674 5448 285680 5460
rect 285732 5448 285738 5500
rect 297818 5448 297824 5500
rect 297876 5488 297882 5500
rect 352098 5488 352104 5500
rect 297876 5460 352104 5488
rect 297876 5448 297882 5460
rect 352098 5448 352104 5460
rect 352156 5448 352162 5500
rect 452562 5448 452568 5500
rect 452620 5488 452626 5500
rect 540514 5488 540520 5500
rect 452620 5460 540520 5488
rect 452620 5448 452626 5460
rect 540514 5448 540520 5460
rect 540572 5448 540578 5500
rect 133782 5380 133788 5432
rect 133840 5420 133846 5432
rect 284294 5420 284300 5432
rect 133840 5392 284300 5420
rect 133840 5380 133846 5392
rect 284294 5380 284300 5392
rect 284352 5380 284358 5432
rect 290734 5380 290740 5432
rect 290792 5420 290798 5432
rect 349338 5420 349344 5432
rect 290792 5392 349344 5420
rect 290792 5380 290798 5392
rect 349338 5380 349344 5392
rect 349396 5380 349402 5432
rect 408402 5380 408408 5432
rect 408460 5420 408466 5432
rect 433518 5420 433524 5432
rect 408460 5392 433524 5420
rect 408460 5380 408466 5392
rect 433518 5380 433524 5392
rect 433576 5380 433582 5432
rect 453850 5380 453856 5432
rect 453908 5420 453914 5432
rect 544102 5420 544108 5432
rect 453908 5392 544108 5420
rect 453908 5380 453914 5392
rect 544102 5380 544108 5392
rect 544160 5380 544166 5432
rect 130194 5312 130200 5364
rect 130252 5352 130258 5364
rect 283190 5352 283196 5364
rect 130252 5324 283196 5352
rect 130252 5312 130258 5324
rect 283190 5312 283196 5324
rect 283248 5312 283254 5364
rect 287146 5312 287152 5364
rect 287204 5352 287210 5364
rect 347958 5352 347964 5364
rect 287204 5324 347964 5352
rect 287204 5312 287210 5324
rect 347958 5312 347964 5324
rect 348016 5312 348022 5364
rect 412358 5312 412364 5364
rect 412416 5352 412422 5364
rect 440602 5352 440608 5364
rect 412416 5324 440608 5352
rect 412416 5312 412422 5324
rect 440602 5312 440608 5324
rect 440660 5312 440666 5364
rect 455322 5312 455328 5364
rect 455380 5352 455386 5364
rect 547690 5352 547696 5364
rect 455380 5324 547696 5352
rect 455380 5312 455386 5324
rect 547690 5312 547696 5324
rect 547748 5312 547754 5364
rect 67174 5244 67180 5296
rect 67232 5284 67238 5296
rect 256970 5284 256976 5296
rect 67232 5256 256976 5284
rect 67232 5244 67238 5256
rect 256970 5244 256976 5256
rect 257028 5244 257034 5296
rect 283650 5244 283656 5296
rect 283708 5284 283714 5296
rect 346578 5284 346584 5296
rect 283708 5256 346584 5284
rect 283708 5244 283714 5256
rect 346578 5244 346584 5256
rect 346636 5244 346642 5296
rect 413830 5244 413836 5296
rect 413888 5284 413894 5296
rect 444190 5284 444196 5296
rect 413888 5256 444196 5284
rect 413888 5244 413894 5256
rect 444190 5244 444196 5256
rect 444248 5244 444254 5296
rect 459462 5244 459468 5296
rect 459520 5284 459526 5296
rect 466089 5287 466147 5293
rect 459520 5256 466040 5284
rect 459520 5244 459526 5256
rect 48130 5176 48136 5228
rect 48188 5216 48194 5228
rect 248506 5216 248512 5228
rect 48188 5188 248512 5216
rect 48188 5176 48194 5188
rect 248506 5176 248512 5188
rect 248564 5176 248570 5228
rect 251450 5176 251456 5228
rect 251508 5216 251514 5228
rect 332594 5216 332600 5228
rect 251508 5188 332600 5216
rect 251508 5176 251514 5188
rect 332594 5176 332600 5188
rect 332652 5176 332658 5228
rect 415302 5176 415308 5228
rect 415360 5216 415366 5228
rect 447778 5216 447784 5228
rect 415360 5188 447784 5216
rect 415360 5176 415366 5188
rect 447778 5176 447784 5188
rect 447836 5176 447842 5228
rect 460842 5176 460848 5228
rect 460900 5216 460906 5228
rect 466012 5216 466040 5256
rect 466089 5253 466101 5287
rect 466135 5284 466147 5287
rect 551186 5284 551192 5296
rect 466135 5256 551192 5284
rect 466135 5253 466147 5256
rect 466089 5247 466147 5253
rect 551186 5244 551192 5256
rect 551244 5244 551250 5296
rect 554774 5216 554780 5228
rect 460900 5188 465948 5216
rect 466012 5188 554780 5216
rect 460900 5176 460906 5188
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 236086 5148 236092 5160
rect 17276 5120 236092 5148
rect 17276 5108 17282 5120
rect 236086 5108 236092 5120
rect 236144 5108 236150 5160
rect 247954 5108 247960 5160
rect 248012 5148 248018 5160
rect 331214 5148 331220 5160
rect 248012 5120 331220 5148
rect 248012 5108 248018 5120
rect 331214 5108 331220 5120
rect 331272 5108 331278 5160
rect 416498 5108 416504 5160
rect 416556 5148 416562 5160
rect 451274 5148 451280 5160
rect 416556 5120 451280 5148
rect 416556 5108 416562 5120
rect 451274 5108 451280 5120
rect 451332 5108 451338 5160
rect 461213 5151 461271 5157
rect 461213 5117 461225 5151
rect 461259 5148 461271 5151
rect 461259 5120 462268 5148
rect 461259 5117 461271 5120
rect 461213 5111 461271 5117
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 234706 5080 234712 5092
rect 12492 5052 234712 5080
rect 12492 5040 12498 5052
rect 234706 5040 234712 5052
rect 234764 5040 234770 5092
rect 244366 5040 244372 5092
rect 244424 5080 244430 5092
rect 321557 5083 321615 5089
rect 321557 5080 321569 5083
rect 244424 5052 321569 5080
rect 244424 5040 244430 5052
rect 321557 5049 321569 5052
rect 321603 5049 321615 5083
rect 321557 5043 321615 5049
rect 321646 5040 321652 5092
rect 321704 5080 321710 5092
rect 327074 5080 327080 5092
rect 321704 5052 327080 5080
rect 321704 5040 321710 5052
rect 327074 5040 327080 5052
rect 327132 5040 327138 5092
rect 327169 5083 327227 5089
rect 327169 5049 327181 5083
rect 327215 5080 327227 5083
rect 329834 5080 329840 5092
rect 327215 5052 329840 5080
rect 327215 5049 327227 5052
rect 327169 5043 327227 5049
rect 329834 5040 329840 5052
rect 329892 5040 329898 5092
rect 337102 5040 337108 5092
rect 337160 5080 337166 5092
rect 368566 5080 368572 5092
rect 337160 5052 368572 5080
rect 337160 5040 337166 5052
rect 368566 5040 368572 5052
rect 368624 5040 368630 5092
rect 376757 5083 376815 5089
rect 376757 5049 376769 5083
rect 376803 5080 376815 5083
rect 381538 5080 381544 5092
rect 376803 5052 381544 5080
rect 376803 5049 376815 5052
rect 376757 5043 376815 5049
rect 381538 5040 381544 5052
rect 381596 5040 381602 5092
rect 417970 5040 417976 5092
rect 418028 5080 418034 5092
rect 454862 5080 454868 5092
rect 418028 5052 454868 5080
rect 418028 5040 418034 5052
rect 454862 5040 454868 5052
rect 454920 5040 454926 5092
rect 458082 5040 458088 5092
rect 458140 5080 458146 5092
rect 458140 5052 462176 5080
rect 458140 5040 458146 5052
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 232130 5012 232136 5024
rect 7708 4984 232136 5012
rect 7708 4972 7714 4984
rect 232130 4972 232136 4984
rect 232188 4972 232194 5024
rect 240778 4972 240784 5024
rect 240836 5012 240842 5024
rect 328730 5012 328736 5024
rect 240836 4984 328736 5012
rect 240836 4972 240842 4984
rect 328730 4972 328736 4984
rect 328788 4972 328794 5024
rect 333606 4972 333612 5024
rect 333664 5012 333670 5024
rect 367186 5012 367192 5024
rect 333664 4984 367192 5012
rect 333664 4972 333670 4984
rect 367186 4972 367192 4984
rect 367244 4972 367250 5024
rect 419442 4972 419448 5024
rect 419500 5012 419506 5024
rect 458450 5012 458456 5024
rect 419500 4984 458456 5012
rect 419500 4972 419506 4984
rect 458450 4972 458456 4984
rect 458508 4972 458514 5024
rect 462038 5012 462044 5024
rect 459388 4984 462044 5012
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 224221 4947 224279 4953
rect 224221 4944 224233 4947
rect 2924 4916 224233 4944
rect 2924 4904 2930 4916
rect 224221 4913 224233 4916
rect 224267 4913 224279 4947
rect 229094 4944 229100 4956
rect 224221 4907 224279 4913
rect 224328 4916 229100 4944
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 224328 4876 224356 4916
rect 229094 4904 229100 4916
rect 229152 4904 229158 4956
rect 237190 4904 237196 4956
rect 237248 4944 237254 4956
rect 321646 4944 321652 4956
rect 237248 4916 321652 4944
rect 237248 4904 237254 4916
rect 321646 4904 321652 4916
rect 321704 4904 321710 4956
rect 321741 4947 321799 4953
rect 321741 4913 321753 4947
rect 321787 4944 321799 4947
rect 326985 4947 327043 4953
rect 326985 4944 326997 4947
rect 321787 4916 326997 4944
rect 321787 4913 321799 4916
rect 321741 4907 321799 4913
rect 326985 4913 326997 4916
rect 327031 4913 327043 4947
rect 326985 4907 327043 4913
rect 327074 4904 327080 4956
rect 327132 4944 327138 4956
rect 361666 4944 361672 4956
rect 327132 4916 361672 4944
rect 327132 4904 327138 4916
rect 361666 4904 361672 4916
rect 361724 4904 361730 4956
rect 376849 4947 376907 4953
rect 376849 4913 376861 4947
rect 376895 4944 376907 4947
rect 380158 4944 380164 4956
rect 376895 4916 380164 4944
rect 376895 4913 376907 4916
rect 376849 4907 376907 4913
rect 380158 4904 380164 4916
rect 380216 4904 380222 4956
rect 420730 4904 420736 4956
rect 420788 4944 420794 4956
rect 459388 4944 459416 4984
rect 462038 4972 462044 4984
rect 462096 4972 462102 5024
rect 420788 4916 459416 4944
rect 462148 4944 462176 5052
rect 462240 5012 462268 5120
rect 463510 5108 463516 5160
rect 463568 5148 463574 5160
rect 465920 5148 465948 5188
rect 554774 5176 554780 5188
rect 554832 5176 554838 5228
rect 558362 5148 558368 5160
rect 463568 5120 465856 5148
rect 465920 5120 558368 5148
rect 463568 5108 463574 5120
rect 464982 5040 464988 5092
rect 465040 5080 465046 5092
rect 465828 5080 465856 5120
rect 558362 5108 558368 5120
rect 558420 5108 558426 5160
rect 471333 5083 471391 5089
rect 465040 5052 465764 5080
rect 465828 5052 471284 5080
rect 465040 5040 465046 5052
rect 465626 5012 465632 5024
rect 462240 4984 465632 5012
rect 465626 4972 465632 4984
rect 465684 4972 465690 5024
rect 465736 5012 465764 5052
rect 471256 5012 471284 5052
rect 471333 5049 471345 5083
rect 471379 5080 471391 5083
rect 561950 5080 561956 5092
rect 471379 5052 561956 5080
rect 471379 5049 471391 5052
rect 471333 5043 471391 5049
rect 561950 5040 561956 5052
rect 562008 5040 562014 5092
rect 565538 5012 565544 5024
rect 465736 4984 471192 5012
rect 471256 4984 565544 5012
rect 466089 4947 466147 4953
rect 466089 4944 466101 4947
rect 462148 4916 466101 4944
rect 420788 4904 420794 4916
rect 466089 4913 466101 4916
rect 466135 4913 466147 4947
rect 466089 4907 466147 4913
rect 466178 4904 466184 4956
rect 466236 4944 466242 4956
rect 471164 4944 471192 4984
rect 565538 4972 565544 4984
rect 565596 4972 565602 5024
rect 569034 4944 569040 4956
rect 466236 4916 471100 4944
rect 471164 4916 569040 4944
rect 466236 4904 466242 4916
rect 624 4848 224356 4876
rect 624 4836 630 4848
rect 230106 4836 230112 4888
rect 230164 4876 230170 4888
rect 324314 4876 324320 4888
rect 230164 4848 324320 4876
rect 230164 4836 230170 4848
rect 324314 4836 324320 4848
rect 324372 4836 324378 4888
rect 326338 4836 326344 4888
rect 326396 4876 326402 4888
rect 360286 4876 360292 4888
rect 326396 4848 360292 4876
rect 326396 4836 326402 4848
rect 360286 4836 360292 4848
rect 360344 4836 360350 4888
rect 422202 4836 422208 4888
rect 422260 4876 422266 4888
rect 461213 4879 461271 4885
rect 461213 4876 461225 4879
rect 422260 4848 461225 4876
rect 422260 4836 422266 4848
rect 461213 4845 461225 4848
rect 461259 4845 461271 4879
rect 469122 4876 469128 4888
rect 461213 4839 461271 4845
rect 461596 4848 469128 4876
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 224129 4811 224187 4817
rect 224129 4808 224141 4811
rect 1728 4780 224141 4808
rect 1728 4768 1734 4780
rect 224129 4777 224141 4780
rect 224175 4777 224187 4811
rect 224129 4771 224187 4777
rect 224221 4811 224279 4817
rect 224221 4777 224233 4811
rect 224267 4808 224279 4811
rect 230750 4808 230756 4820
rect 224267 4780 230756 4808
rect 224267 4777 224279 4780
rect 224221 4771 224279 4777
rect 230750 4768 230756 4780
rect 230808 4768 230814 4820
rect 233694 4768 233700 4820
rect 233752 4808 233758 4820
rect 325694 4808 325700 4820
rect 233752 4780 325700 4808
rect 233752 4768 233758 4780
rect 325694 4768 325700 4780
rect 325752 4768 325758 4820
rect 328454 4768 328460 4820
rect 328512 4808 328518 4820
rect 363046 4808 363052 4820
rect 328512 4780 363052 4808
rect 328512 4768 328518 4780
rect 363046 4768 363052 4780
rect 363104 4768 363110 4820
rect 423582 4768 423588 4820
rect 423640 4808 423646 4820
rect 461596 4808 461624 4848
rect 469122 4836 469128 4848
rect 469180 4836 469186 4888
rect 471072 4876 471100 4916
rect 569034 4904 569040 4916
rect 569092 4904 569098 4956
rect 572622 4876 572628 4888
rect 471072 4848 572628 4876
rect 572622 4836 572628 4848
rect 572680 4836 572686 4888
rect 423640 4780 461624 4808
rect 423640 4768 423646 4780
rect 462130 4768 462136 4820
rect 462188 4808 462194 4820
rect 471333 4811 471391 4817
rect 471333 4808 471345 4811
rect 462188 4780 471345 4808
rect 462188 4768 462194 4780
rect 471333 4777 471345 4780
rect 471379 4777 471391 4811
rect 471333 4771 471391 4777
rect 471425 4811 471483 4817
rect 471425 4777 471437 4811
rect 471471 4808 471483 4811
rect 579798 4808 579804 4820
rect 471471 4780 579804 4808
rect 471471 4777 471483 4780
rect 471425 4771 471483 4777
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 212258 4700 212264 4752
rect 212316 4740 212322 4752
rect 316034 4740 316040 4752
rect 212316 4712 316040 4740
rect 212316 4700 212322 4712
rect 316034 4700 316040 4712
rect 316092 4700 316098 4752
rect 318702 4700 318708 4752
rect 318760 4740 318766 4752
rect 318760 4712 323256 4740
rect 318760 4700 318766 4712
rect 215846 4632 215852 4684
rect 215904 4672 215910 4684
rect 317414 4672 317420 4684
rect 215904 4644 317420 4672
rect 215904 4632 215910 4644
rect 317414 4632 317420 4644
rect 317472 4632 317478 4684
rect 323228 4672 323256 4712
rect 323302 4700 323308 4752
rect 323360 4740 323366 4752
rect 359182 4740 359188 4752
rect 323360 4712 359188 4740
rect 323360 4700 323366 4712
rect 359182 4700 359188 4712
rect 359240 4700 359246 4752
rect 451090 4700 451096 4752
rect 451148 4740 451154 4752
rect 536926 4740 536932 4752
rect 451148 4712 536932 4740
rect 451148 4700 451154 4712
rect 536926 4700 536932 4712
rect 536984 4700 536990 4752
rect 333974 4672 333980 4684
rect 323228 4644 333980 4672
rect 333974 4632 333980 4644
rect 334032 4632 334038 4684
rect 449802 4632 449808 4684
rect 449860 4672 449866 4684
rect 533430 4672 533436 4684
rect 449860 4644 533436 4672
rect 449860 4632 449866 4644
rect 533430 4632 533436 4644
rect 533488 4632 533494 4684
rect 219342 4564 219348 4616
rect 219400 4604 219406 4616
rect 318794 4604 318800 4616
rect 219400 4576 318800 4604
rect 219400 4564 219406 4576
rect 318794 4564 318800 4576
rect 318852 4564 318858 4616
rect 321370 4604 321376 4616
rect 318904 4576 321376 4604
rect 222930 4496 222936 4548
rect 222988 4536 222994 4548
rect 318904 4536 318932 4576
rect 321370 4564 321376 4576
rect 321428 4564 321434 4616
rect 322750 4564 322756 4616
rect 322808 4604 322814 4616
rect 337105 4607 337163 4613
rect 337105 4604 337117 4607
rect 322808 4576 337117 4604
rect 322808 4564 322814 4576
rect 337105 4573 337117 4576
rect 337151 4573 337163 4607
rect 337105 4567 337163 4573
rect 448330 4564 448336 4616
rect 448388 4604 448394 4616
rect 529842 4604 529848 4616
rect 448388 4576 529848 4604
rect 448388 4564 448394 4576
rect 529842 4564 529848 4576
rect 529900 4564 529906 4616
rect 222988 4508 318932 4536
rect 222988 4496 222994 4508
rect 320358 4496 320364 4548
rect 320416 4536 320422 4548
rect 335354 4536 335360 4548
rect 320416 4508 335360 4536
rect 320416 4496 320422 4508
rect 335354 4496 335360 4508
rect 335412 4496 335418 4548
rect 447042 4496 447048 4548
rect 447100 4536 447106 4548
rect 526254 4536 526260 4548
rect 447100 4508 526260 4536
rect 447100 4496 447106 4508
rect 526254 4496 526260 4508
rect 526312 4496 526318 4548
rect 226518 4428 226524 4480
rect 226576 4468 226582 4480
rect 322934 4468 322940 4480
rect 226576 4440 322940 4468
rect 226576 4428 226582 4440
rect 322934 4428 322940 4440
rect 322992 4428 322998 4480
rect 325142 4428 325148 4480
rect 325200 4468 325206 4480
rect 338114 4468 338120 4480
rect 325200 4440 338120 4468
rect 325200 4428 325206 4440
rect 338114 4428 338120 4440
rect 338172 4428 338178 4480
rect 445570 4428 445576 4480
rect 445628 4468 445634 4480
rect 522666 4468 522672 4480
rect 445628 4440 522672 4468
rect 445628 4428 445634 4440
rect 522666 4428 522672 4440
rect 522724 4428 522730 4480
rect 201494 4360 201500 4412
rect 201552 4400 201558 4412
rect 271138 4400 271144 4412
rect 201552 4372 271144 4400
rect 201552 4360 201558 4372
rect 271138 4360 271144 4372
rect 271196 4360 271202 4412
rect 301406 4360 301412 4412
rect 301464 4400 301470 4412
rect 353478 4400 353484 4412
rect 301464 4372 353484 4400
rect 301464 4360 301470 4372
rect 353478 4360 353484 4372
rect 353536 4360 353542 4412
rect 354861 4403 354919 4409
rect 354861 4369 354873 4403
rect 354907 4400 354919 4403
rect 356057 4403 356115 4409
rect 356057 4400 356069 4403
rect 354907 4372 356069 4400
rect 354907 4369 354919 4372
rect 354861 4363 354919 4369
rect 356057 4369 356069 4372
rect 356103 4369 356115 4403
rect 356057 4363 356115 4369
rect 444282 4360 444288 4412
rect 444340 4400 444346 4412
rect 519078 4400 519084 4412
rect 444340 4372 519084 4400
rect 444340 4360 444346 4372
rect 519078 4360 519084 4372
rect 519136 4360 519142 4412
rect 205082 4292 205088 4344
rect 205140 4332 205146 4344
rect 272518 4332 272524 4344
rect 205140 4304 272524 4332
rect 205140 4292 205146 4304
rect 272518 4292 272524 4304
rect 272576 4292 272582 4344
rect 304994 4292 305000 4344
rect 305052 4332 305058 4344
rect 354950 4332 354956 4344
rect 305052 4304 354956 4332
rect 305052 4292 305058 4304
rect 354950 4292 354956 4304
rect 355008 4292 355014 4344
rect 442902 4292 442908 4344
rect 442960 4332 442966 4344
rect 515582 4332 515588 4344
rect 442960 4304 515588 4332
rect 442960 4292 442966 4304
rect 515582 4292 515588 4304
rect 515640 4292 515646 4344
rect 224129 4267 224187 4273
rect 224129 4233 224141 4267
rect 224175 4264 224187 4267
rect 230566 4264 230572 4276
rect 224175 4236 230572 4264
rect 224175 4233 224187 4236
rect 224129 4227 224187 4233
rect 230566 4224 230572 4236
rect 230624 4224 230630 4276
rect 308582 4224 308588 4276
rect 308640 4264 308646 4276
rect 356146 4264 356152 4276
rect 308640 4236 356152 4264
rect 308640 4224 308646 4236
rect 356146 4224 356152 4236
rect 356204 4224 356210 4276
rect 441522 4224 441528 4276
rect 441580 4264 441586 4276
rect 511994 4264 512000 4276
rect 441580 4236 512000 4264
rect 441580 4224 441586 4236
rect 511994 4224 512000 4236
rect 512052 4224 512058 4276
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 140866 4156 140872 4208
rect 140924 4196 140930 4208
rect 142062 4196 142068 4208
rect 140924 4168 142068 4196
rect 140924 4156 140930 4168
rect 142062 4156 142068 4168
rect 142120 4156 142126 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 160002 4196 160008 4208
rect 158772 4168 160008 4196
rect 158772 4156 158778 4168
rect 160002 4156 160008 4168
rect 160060 4156 160066 4208
rect 175366 4156 175372 4208
rect 175424 4196 175430 4208
rect 176562 4196 176568 4208
rect 175424 4168 176568 4196
rect 175424 4156 175430 4168
rect 176562 4156 176568 4168
rect 176620 4156 176626 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 287609 4199 287667 4205
rect 284680 4168 285720 4196
rect 34974 4088 34980 4140
rect 35032 4128 35038 4140
rect 50338 4128 50344 4140
rect 35032 4100 50344 4128
rect 35032 4088 35038 4100
rect 50338 4088 50344 4100
rect 50396 4088 50402 4140
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 250438 4128 250444 4140
rect 57664 4100 250444 4128
rect 57664 4088 57670 4100
rect 250438 4088 250444 4100
rect 250496 4088 250502 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269022 4128 269028 4140
rect 268160 4100 269028 4128
rect 268160 4088 268166 4100
rect 269022 4088 269028 4100
rect 269080 4088 269086 4140
rect 278041 4131 278099 4137
rect 278041 4097 278053 4131
rect 278087 4128 278099 4131
rect 284680 4128 284708 4168
rect 278087 4100 284708 4128
rect 278087 4097 278099 4100
rect 278041 4091 278099 4097
rect 284754 4088 284760 4140
rect 284812 4128 284818 4140
rect 285582 4128 285588 4140
rect 284812 4100 285588 4128
rect 284812 4088 284818 4100
rect 285582 4088 285588 4100
rect 285640 4088 285646 4140
rect 285692 4128 285720 4168
rect 287609 4165 287621 4199
rect 287655 4196 287667 4199
rect 287655 4168 287928 4196
rect 287655 4165 287667 4168
rect 287609 4159 287667 4165
rect 287900 4128 287928 4168
rect 312170 4156 312176 4208
rect 312228 4196 312234 4208
rect 357710 4196 357716 4208
rect 312228 4168 357716 4196
rect 312228 4156 312234 4168
rect 357710 4156 357716 4168
rect 357768 4156 357774 4208
rect 424962 4156 424968 4208
rect 425020 4196 425026 4208
rect 472710 4196 472716 4208
rect 425020 4168 472716 4196
rect 425020 4156 425026 4168
rect 472710 4156 472716 4168
rect 472768 4156 472774 4208
rect 295886 4128 295892 4140
rect 285692 4100 287836 4128
rect 287900 4100 295892 4128
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 28258 4060 28264 4072
rect 20772 4032 28264 4060
rect 20772 4020 20778 4032
rect 28258 4020 28264 4032
rect 28316 4020 28322 4072
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 249058 4060 249064 4072
rect 50580 4032 249064 4060
rect 50580 4020 50586 4032
rect 249058 4020 249064 4032
rect 249116 4020 249122 4072
rect 264609 4063 264667 4069
rect 264609 4029 264621 4063
rect 264655 4060 264667 4063
rect 282917 4063 282975 4069
rect 282917 4060 282929 4063
rect 264655 4032 282929 4060
rect 264655 4029 264667 4032
rect 264609 4023 264667 4029
rect 282917 4029 282929 4032
rect 282963 4029 282975 4063
rect 287808 4060 287836 4100
rect 295886 4088 295892 4100
rect 295944 4088 295950 4140
rect 296714 4088 296720 4140
rect 296772 4128 296778 4140
rect 297910 4128 297916 4140
rect 296772 4100 297916 4128
rect 296772 4088 296778 4100
rect 297910 4088 297916 4100
rect 297968 4088 297974 4140
rect 300302 4088 300308 4140
rect 300360 4128 300366 4140
rect 332321 4131 332379 4137
rect 332321 4128 332333 4131
rect 300360 4100 332333 4128
rect 300360 4088 300366 4100
rect 332321 4097 332333 4100
rect 332367 4097 332379 4131
rect 332321 4091 332379 4097
rect 332410 4088 332416 4140
rect 332468 4128 332474 4140
rect 333238 4128 333244 4140
rect 332468 4100 333244 4128
rect 332468 4088 332474 4100
rect 333238 4088 333244 4100
rect 333296 4088 333302 4140
rect 334710 4088 334716 4140
rect 334768 4128 334774 4140
rect 335262 4128 335268 4140
rect 334768 4100 335268 4128
rect 334768 4088 334774 4100
rect 335262 4088 335268 4100
rect 335320 4088 335326 4140
rect 335357 4131 335415 4137
rect 335357 4097 335369 4131
rect 335403 4128 335415 4131
rect 338758 4128 338764 4140
rect 335403 4100 338764 4128
rect 335403 4097 335415 4100
rect 335357 4091 335415 4097
rect 338758 4088 338764 4100
rect 338816 4088 338822 4140
rect 339494 4088 339500 4140
rect 339552 4128 339558 4140
rect 340782 4128 340788 4140
rect 339552 4100 340788 4128
rect 339552 4088 339558 4100
rect 340782 4088 340788 4100
rect 340840 4088 340846 4140
rect 341245 4131 341303 4137
rect 341245 4097 341257 4131
rect 341291 4128 341303 4131
rect 345658 4128 345664 4140
rect 341291 4100 345664 4128
rect 341291 4097 341303 4100
rect 341245 4091 341303 4097
rect 345658 4088 345664 4100
rect 345716 4088 345722 4140
rect 347866 4088 347872 4140
rect 347924 4128 347930 4140
rect 349062 4128 349068 4140
rect 347924 4100 349068 4128
rect 347924 4088 347930 4100
rect 349062 4088 349068 4100
rect 349120 4088 349126 4140
rect 349157 4131 349215 4137
rect 349157 4097 349169 4131
rect 349203 4128 349215 4131
rect 351178 4128 351184 4140
rect 349203 4100 351184 4128
rect 349203 4097 349215 4100
rect 349157 4091 349215 4097
rect 351178 4088 351184 4100
rect 351236 4088 351242 4140
rect 351362 4088 351368 4140
rect 351420 4128 351426 4140
rect 351822 4128 351828 4140
rect 351420 4100 351828 4128
rect 351420 4088 351426 4100
rect 351822 4088 351828 4100
rect 351880 4088 351886 4140
rect 352009 4131 352067 4137
rect 352009 4097 352021 4131
rect 352055 4128 352067 4131
rect 354861 4131 354919 4137
rect 354861 4128 354873 4131
rect 352055 4100 354873 4128
rect 352055 4097 352067 4100
rect 352009 4091 352067 4097
rect 354861 4097 354873 4100
rect 354907 4097 354919 4131
rect 354861 4091 354919 4097
rect 354950 4088 354956 4140
rect 355008 4128 355014 4140
rect 355962 4128 355968 4140
rect 355008 4100 355968 4128
rect 355008 4088 355014 4100
rect 355962 4088 355968 4100
rect 356020 4088 356026 4140
rect 356057 4131 356115 4137
rect 356057 4097 356069 4131
rect 356103 4128 356115 4131
rect 358078 4128 358084 4140
rect 356103 4100 358084 4128
rect 356103 4097 356115 4100
rect 356057 4091 356115 4097
rect 358078 4088 358084 4100
rect 358136 4088 358142 4140
rect 362126 4088 362132 4140
rect 362184 4128 362190 4140
rect 362862 4128 362868 4140
rect 362184 4100 362868 4128
rect 362184 4088 362190 4100
rect 362862 4088 362868 4100
rect 362920 4088 362926 4140
rect 363322 4088 363328 4140
rect 363380 4128 363386 4140
rect 364242 4128 364248 4140
rect 363380 4100 364248 4128
rect 363380 4088 363386 4100
rect 364242 4088 364248 4100
rect 364300 4088 364306 4140
rect 365714 4088 365720 4140
rect 365772 4128 365778 4140
rect 366910 4128 366916 4140
rect 365772 4100 366916 4128
rect 365772 4088 365778 4100
rect 366910 4088 366916 4100
rect 366968 4088 366974 4140
rect 369210 4088 369216 4140
rect 369268 4128 369274 4140
rect 369762 4128 369768 4140
rect 369268 4100 369768 4128
rect 369268 4088 369274 4100
rect 369762 4088 369768 4100
rect 369820 4088 369826 4140
rect 370406 4088 370412 4140
rect 370464 4128 370470 4140
rect 371142 4128 371148 4140
rect 370464 4100 371148 4128
rect 370464 4088 370470 4100
rect 371142 4088 371148 4100
rect 371200 4088 371206 4140
rect 377582 4088 377588 4140
rect 377640 4128 377646 4140
rect 378042 4128 378048 4140
rect 377640 4100 378048 4128
rect 377640 4088 377646 4100
rect 378042 4088 378048 4100
rect 378100 4088 378106 4140
rect 378778 4088 378784 4140
rect 378836 4128 378842 4140
rect 385310 4128 385316 4140
rect 378836 4100 385316 4128
rect 378836 4088 378842 4100
rect 385310 4088 385316 4100
rect 385368 4088 385374 4140
rect 390554 4088 390560 4140
rect 390612 4128 390618 4140
rect 391842 4128 391848 4140
rect 390612 4100 391848 4128
rect 390612 4088 390618 4100
rect 391842 4088 391848 4100
rect 391900 4088 391906 4140
rect 393130 4088 393136 4140
rect 393188 4128 393194 4140
rect 395430 4128 395436 4140
rect 393188 4100 395436 4128
rect 393188 4088 393194 4100
rect 395430 4088 395436 4100
rect 395488 4088 395494 4140
rect 398098 4088 398104 4140
rect 398156 4128 398162 4140
rect 403710 4128 403716 4140
rect 398156 4100 403716 4128
rect 398156 4088 398162 4100
rect 403710 4088 403716 4100
rect 403768 4088 403774 4140
rect 414017 4131 414075 4137
rect 414017 4097 414029 4131
rect 414063 4128 414075 4131
rect 438210 4128 438216 4140
rect 414063 4100 438216 4128
rect 414063 4097 414075 4100
rect 414017 4091 414075 4097
rect 438210 4088 438216 4100
rect 438268 4088 438274 4140
rect 442258 4088 442264 4140
rect 442316 4128 442322 4140
rect 445481 4131 445539 4137
rect 445481 4128 445493 4131
rect 442316 4100 445493 4128
rect 442316 4088 442322 4100
rect 445481 4097 445493 4100
rect 445527 4097 445539 4131
rect 445481 4091 445539 4097
rect 445662 4088 445668 4140
rect 445720 4128 445726 4140
rect 521470 4128 521476 4140
rect 445720 4100 521476 4128
rect 445720 4088 445726 4100
rect 521470 4088 521476 4100
rect 521528 4088 521534 4140
rect 529198 4088 529204 4140
rect 529256 4128 529262 4140
rect 575014 4128 575020 4140
rect 529256 4100 575020 4128
rect 529256 4088 529262 4100
rect 575014 4088 575020 4100
rect 575072 4088 575078 4140
rect 298094 4060 298100 4072
rect 287808 4032 298100 4060
rect 282917 4023 282975 4029
rect 298094 4020 298100 4032
rect 298152 4020 298158 4072
rect 302602 4020 302608 4072
rect 302660 4060 302666 4072
rect 309778 4060 309784 4072
rect 302660 4032 309784 4060
rect 302660 4020 302666 4032
rect 309778 4020 309784 4032
rect 309836 4020 309842 4072
rect 313366 4020 313372 4072
rect 313424 4060 313430 4072
rect 352377 4063 352435 4069
rect 313424 4032 352328 4060
rect 313424 4020 313430 4032
rect 46934 3952 46940 4004
rect 46992 3992 46998 4004
rect 248690 3992 248696 4004
rect 46992 3964 248696 3992
rect 46992 3952 46998 3964
rect 248690 3952 248696 3964
rect 248748 3952 248754 4004
rect 257430 3952 257436 4004
rect 257488 3992 257494 4004
rect 287609 3995 287667 4001
rect 287609 3992 287621 3995
rect 257488 3964 287621 3992
rect 257488 3952 257494 3964
rect 287609 3961 287621 3964
rect 287655 3961 287667 3995
rect 287609 3955 287667 3961
rect 287701 3995 287759 4001
rect 287701 3961 287713 3995
rect 287747 3992 287759 3995
rect 297358 3992 297364 4004
rect 287747 3964 297364 3992
rect 287747 3961 287759 3964
rect 287701 3955 287759 3961
rect 297358 3952 297364 3964
rect 297416 3952 297422 4004
rect 314562 3952 314568 4004
rect 314620 3992 314626 4004
rect 352193 3995 352251 4001
rect 352193 3992 352205 3995
rect 314620 3964 352205 3992
rect 314620 3952 314626 3964
rect 352193 3961 352205 3964
rect 352239 3961 352251 3995
rect 352300 3992 352328 4032
rect 352377 4029 352389 4063
rect 352423 4060 352435 4063
rect 373994 4060 374000 4072
rect 352423 4032 374000 4060
rect 352423 4029 352435 4032
rect 352377 4023 352435 4029
rect 373994 4020 374000 4032
rect 374052 4020 374058 4072
rect 376754 4020 376760 4072
rect 376812 4020 376818 4072
rect 383562 4020 383568 4072
rect 383620 4060 383626 4072
rect 384298 4060 384304 4072
rect 383620 4032 384304 4060
rect 383620 4020 383626 4032
rect 384298 4020 384304 4032
rect 384356 4020 384362 4072
rect 393222 4020 393228 4072
rect 393280 4060 393286 4072
rect 396626 4060 396632 4072
rect 393280 4032 396632 4060
rect 393280 4020 393286 4032
rect 396626 4020 396632 4032
rect 396684 4020 396690 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 439406 4060 439412 4072
rect 411220 4032 439412 4060
rect 411220 4020 411226 4032
rect 439406 4020 439412 4032
rect 439464 4020 439470 4072
rect 439590 4020 439596 4072
rect 439648 4060 439654 4072
rect 446309 4063 446367 4069
rect 446309 4060 446321 4063
rect 439648 4032 446321 4060
rect 439648 4020 439654 4032
rect 446309 4029 446321 4032
rect 446355 4029 446367 4063
rect 446309 4023 446367 4029
rect 448422 4020 448428 4072
rect 448480 4060 448486 4072
rect 528646 4060 528652 4072
rect 448480 4032 528652 4060
rect 448480 4020 448486 4032
rect 528646 4020 528652 4032
rect 528704 4020 528710 4072
rect 530578 4020 530584 4072
rect 530636 4060 530642 4072
rect 582190 4060 582196 4072
rect 530636 4032 582196 4060
rect 530636 4020 530642 4032
rect 582190 4020 582196 4032
rect 582248 4020 582254 4072
rect 358814 3992 358820 4004
rect 352300 3964 358820 3992
rect 352193 3955 352251 3961
rect 358814 3952 358820 3964
rect 358872 3952 358878 4004
rect 359734 3952 359740 4004
rect 359792 3992 359798 4004
rect 376772 3992 376800 4020
rect 359792 3964 376800 3992
rect 359792 3952 359798 3964
rect 402882 3952 402888 4004
rect 402940 3992 402946 4004
rect 419166 3992 419172 4004
rect 402940 3964 419172 3992
rect 402940 3952 402946 3964
rect 419166 3952 419172 3964
rect 419224 3952 419230 4004
rect 420270 3952 420276 4004
rect 420328 3992 420334 4004
rect 423950 3992 423956 4004
rect 420328 3964 423956 3992
rect 420328 3952 420334 3964
rect 423950 3952 423956 3964
rect 424008 3952 424014 4004
rect 424594 3952 424600 4004
rect 424652 3992 424658 4004
rect 425146 3992 425152 4004
rect 424652 3964 425152 3992
rect 424652 3952 424658 3964
rect 425146 3952 425152 3964
rect 425204 3952 425210 4004
rect 425241 3995 425299 4001
rect 425241 3961 425253 3995
rect 425287 3992 425299 3995
rect 450170 3992 450176 4004
rect 425287 3964 450176 3992
rect 425287 3961 425299 3964
rect 425241 3955 425299 3961
rect 450170 3952 450176 3964
rect 450228 3952 450234 4004
rect 451182 3952 451188 4004
rect 451240 3992 451246 4004
rect 535730 3992 535736 4004
rect 451240 3964 535736 3992
rect 451240 3952 451246 3964
rect 535730 3952 535736 3964
rect 535788 3952 535794 4004
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 247678 3924 247684 3936
rect 45796 3896 247684 3924
rect 45796 3884 45802 3896
rect 247678 3884 247684 3896
rect 247736 3884 247742 3936
rect 282454 3884 282460 3936
rect 282512 3924 282518 3936
rect 320821 3927 320879 3933
rect 320821 3924 320833 3927
rect 282512 3896 320833 3924
rect 282512 3884 282518 3896
rect 320821 3893 320833 3896
rect 320867 3893 320879 3927
rect 320821 3887 320879 3893
rect 326341 3927 326399 3933
rect 326341 3893 326353 3927
rect 326387 3924 326399 3927
rect 332229 3927 332287 3933
rect 332229 3924 332241 3927
rect 326387 3896 332241 3924
rect 326387 3893 326399 3896
rect 326341 3887 326399 3893
rect 332229 3893 332241 3896
rect 332275 3893 332287 3927
rect 332229 3887 332287 3893
rect 332321 3927 332379 3933
rect 332321 3893 332333 3927
rect 332367 3924 332379 3927
rect 336185 3927 336243 3933
rect 332367 3896 336136 3924
rect 332367 3893 332379 3896
rect 332321 3887 332379 3893
rect 39758 3816 39764 3868
rect 39816 3856 39822 3868
rect 245746 3856 245752 3868
rect 39816 3828 245752 3856
rect 39816 3816 39822 3828
rect 245746 3816 245752 3828
rect 245804 3816 245810 3868
rect 264606 3816 264612 3868
rect 264664 3856 264670 3868
rect 278041 3859 278099 3865
rect 278041 3856 278053 3859
rect 264664 3828 278053 3856
rect 264664 3816 264670 3828
rect 278041 3825 278053 3828
rect 278087 3825 278099 3859
rect 288621 3859 288679 3865
rect 288621 3856 288633 3859
rect 278041 3819 278099 3825
rect 285876 3828 288633 3856
rect 19518 3748 19524 3800
rect 19576 3788 19582 3800
rect 32398 3788 32404 3800
rect 19576 3760 32404 3788
rect 19576 3748 19582 3760
rect 32398 3748 32404 3760
rect 32456 3748 32462 3800
rect 38562 3748 38568 3800
rect 38620 3788 38626 3800
rect 245654 3788 245660 3800
rect 38620 3760 245660 3788
rect 38620 3748 38626 3760
rect 245654 3748 245660 3760
rect 245712 3748 245718 3800
rect 278866 3748 278872 3800
rect 278924 3788 278930 3800
rect 285876 3788 285904 3828
rect 288621 3825 288633 3828
rect 288667 3825 288679 3859
rect 288621 3819 288679 3825
rect 289538 3816 289544 3868
rect 289596 3856 289602 3868
rect 336108 3856 336136 3896
rect 336185 3893 336197 3927
rect 336231 3924 336243 3927
rect 365806 3924 365812 3936
rect 336231 3896 365812 3924
rect 336231 3893 336243 3896
rect 336185 3887 336243 3893
rect 365806 3884 365812 3896
rect 365864 3884 365870 3936
rect 371602 3884 371608 3936
rect 371660 3924 371666 3936
rect 376757 3927 376815 3933
rect 376757 3924 376769 3927
rect 371660 3896 376769 3924
rect 371660 3884 371666 3896
rect 376757 3893 376769 3896
rect 376803 3893 376815 3927
rect 376757 3887 376815 3893
rect 412450 3884 412456 3936
rect 412508 3924 412514 3936
rect 441614 3924 441620 3936
rect 412508 3896 441620 3924
rect 412508 3884 412514 3896
rect 441614 3884 441620 3896
rect 441672 3884 441678 3936
rect 441709 3927 441767 3933
rect 441709 3893 441721 3927
rect 441755 3924 441767 3927
rect 453666 3924 453672 3936
rect 441755 3896 453672 3924
rect 441755 3893 441767 3896
rect 441709 3887 441767 3893
rect 453666 3884 453672 3896
rect 453724 3884 453730 3936
rect 453942 3884 453948 3936
rect 454000 3924 454006 3936
rect 542906 3924 542912 3936
rect 454000 3896 542912 3924
rect 454000 3884 454006 3896
rect 542906 3884 542912 3896
rect 542964 3884 542970 3936
rect 342898 3856 342904 3868
rect 289596 3828 336044 3856
rect 336108 3828 342904 3856
rect 289596 3816 289602 3828
rect 278924 3760 285904 3788
rect 278924 3748 278930 3760
rect 285950 3748 285956 3800
rect 286008 3788 286014 3800
rect 332137 3791 332195 3797
rect 332137 3788 332149 3791
rect 286008 3760 332149 3788
rect 286008 3748 286014 3760
rect 332137 3757 332149 3760
rect 332183 3757 332195 3791
rect 332137 3751 332195 3757
rect 332229 3791 332287 3797
rect 332229 3757 332241 3791
rect 332275 3788 332287 3791
rect 335814 3788 335820 3800
rect 332275 3760 335820 3788
rect 332275 3757 332287 3760
rect 332229 3751 332287 3757
rect 335814 3748 335820 3760
rect 335872 3748 335878 3800
rect 336016 3788 336044 3828
rect 342898 3816 342904 3828
rect 342956 3816 342962 3868
rect 343082 3816 343088 3868
rect 343140 3856 343146 3868
rect 369118 3856 369124 3868
rect 343140 3828 369124 3856
rect 343140 3816 343146 3828
rect 369118 3816 369124 3828
rect 369176 3816 369182 3868
rect 372798 3816 372804 3868
rect 372856 3856 372862 3868
rect 373902 3856 373908 3868
rect 372856 3828 373908 3856
rect 372856 3816 372862 3828
rect 373902 3816 373908 3828
rect 373960 3816 373966 3868
rect 413922 3816 413928 3868
rect 413980 3856 413986 3868
rect 445386 3856 445392 3868
rect 413980 3828 445392 3856
rect 413980 3816 413986 3828
rect 445386 3816 445392 3828
rect 445444 3816 445450 3868
rect 445481 3859 445539 3865
rect 445481 3825 445493 3859
rect 445527 3856 445539 3859
rect 451921 3859 451979 3865
rect 451921 3856 451933 3859
rect 445527 3828 451933 3856
rect 445527 3825 445539 3828
rect 445481 3819 445539 3825
rect 451921 3825 451933 3828
rect 451967 3825 451979 3859
rect 451921 3819 451979 3825
rect 466365 3859 466423 3865
rect 466365 3825 466377 3859
rect 466411 3856 466423 3859
rect 550082 3856 550088 3868
rect 466411 3828 550088 3856
rect 466411 3825 466423 3828
rect 466365 3819 466423 3825
rect 550082 3816 550088 3828
rect 550140 3816 550146 3868
rect 341518 3788 341524 3800
rect 336016 3760 341524 3788
rect 341518 3748 341524 3760
rect 341576 3748 341582 3800
rect 341886 3748 341892 3800
rect 341944 3788 341950 3800
rect 370130 3788 370136 3800
rect 341944 3760 370136 3788
rect 341944 3748 341950 3760
rect 370130 3748 370136 3760
rect 370188 3748 370194 3800
rect 373994 3748 374000 3800
rect 374052 3788 374058 3800
rect 375282 3788 375288 3800
rect 374052 3760 375288 3788
rect 374052 3748 374058 3760
rect 375282 3748 375288 3760
rect 375340 3748 375346 3800
rect 399478 3748 399484 3800
rect 399536 3788 399542 3800
rect 408494 3788 408500 3800
rect 399536 3760 408500 3788
rect 399536 3748 399542 3760
rect 408494 3748 408500 3760
rect 408552 3748 408558 3800
rect 411070 3748 411076 3800
rect 411128 3788 411134 3800
rect 414017 3791 414075 3797
rect 414017 3788 414029 3791
rect 411128 3760 414029 3788
rect 411128 3748 411134 3760
rect 414017 3757 414029 3760
rect 414063 3757 414075 3791
rect 442994 3788 443000 3800
rect 414017 3751 414075 3757
rect 417436 3760 443000 3788
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 243078 3720 243084 3732
rect 32732 3692 243084 3720
rect 32732 3680 32738 3692
rect 243078 3680 243084 3692
rect 243136 3680 243142 3732
rect 282917 3723 282975 3729
rect 282917 3689 282929 3723
rect 282963 3720 282975 3723
rect 287701 3723 287759 3729
rect 287701 3720 287713 3723
rect 282963 3692 287713 3720
rect 282963 3689 282975 3692
rect 282917 3683 282975 3689
rect 287701 3689 287713 3692
rect 287747 3689 287759 3723
rect 287701 3683 287759 3689
rect 292485 3723 292543 3729
rect 292485 3689 292497 3723
rect 292531 3720 292543 3723
rect 326341 3723 326399 3729
rect 326341 3720 326353 3723
rect 292531 3692 326353 3720
rect 292531 3689 292543 3692
rect 292485 3683 292543 3689
rect 326341 3689 326353 3692
rect 326387 3689 326399 3723
rect 326341 3683 326399 3689
rect 326430 3680 326436 3732
rect 326488 3720 326494 3732
rect 328454 3720 328460 3732
rect 326488 3692 328460 3720
rect 326488 3680 326494 3692
rect 328454 3680 328460 3692
rect 328512 3680 328518 3732
rect 331214 3680 331220 3732
rect 331272 3720 331278 3732
rect 336185 3723 336243 3729
rect 336185 3720 336197 3723
rect 331272 3692 336197 3720
rect 331272 3680 331278 3692
rect 336185 3689 336197 3692
rect 336231 3689 336243 3723
rect 336185 3683 336243 3689
rect 338298 3680 338304 3732
rect 338356 3720 338362 3732
rect 368658 3720 368664 3732
rect 338356 3692 368664 3720
rect 338356 3680 338362 3692
rect 368658 3680 368664 3692
rect 368716 3680 368722 3732
rect 375190 3680 375196 3732
rect 375248 3720 375254 3732
rect 383838 3720 383844 3732
rect 375248 3692 383844 3720
rect 375248 3680 375254 3692
rect 383838 3680 383844 3692
rect 383896 3680 383902 3732
rect 400122 3680 400128 3732
rect 400180 3720 400186 3732
rect 412082 3720 412088 3732
rect 400180 3692 412088 3720
rect 400180 3680 400186 3692
rect 412082 3680 412088 3692
rect 412140 3680 412146 3732
rect 412542 3680 412548 3732
rect 412600 3720 412606 3732
rect 417436 3720 417464 3760
rect 442994 3748 443000 3760
rect 443052 3748 443058 3800
rect 443089 3791 443147 3797
rect 443089 3757 443101 3791
rect 443135 3788 443147 3791
rect 446677 3791 446735 3797
rect 446677 3788 446689 3791
rect 443135 3760 446689 3788
rect 443135 3757 443147 3760
rect 443089 3751 443147 3757
rect 446677 3757 446689 3760
rect 446723 3757 446735 3791
rect 452470 3788 452476 3800
rect 446677 3751 446735 3757
rect 446784 3760 452476 3788
rect 422849 3723 422907 3729
rect 422849 3720 422861 3723
rect 412600 3692 417464 3720
rect 417528 3692 422861 3720
rect 412600 3680 412606 3692
rect 24302 3612 24308 3664
rect 24360 3652 24366 3664
rect 239030 3652 239036 3664
rect 24360 3624 239036 3652
rect 24360 3612 24366 3624
rect 239030 3612 239036 3624
rect 239088 3612 239094 3664
rect 262214 3612 262220 3664
rect 262272 3652 262278 3664
rect 320637 3655 320695 3661
rect 320637 3652 320649 3655
rect 262272 3624 320649 3652
rect 262272 3612 262278 3624
rect 320637 3621 320649 3624
rect 320683 3621 320695 3655
rect 325142 3652 325148 3664
rect 320637 3615 320695 3621
rect 320744 3624 325148 3652
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 19978 3584 19984 3596
rect 11296 3556 19984 3584
rect 11296 3544 11302 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 240318 3584 240324 3596
rect 25556 3556 240324 3584
rect 25556 3544 25562 3556
rect 240318 3544 240324 3556
rect 240376 3544 240382 3596
rect 265802 3544 265808 3596
rect 265860 3584 265866 3596
rect 320744 3584 320772 3624
rect 325142 3612 325148 3624
rect 325200 3612 325206 3664
rect 325234 3612 325240 3664
rect 325292 3652 325298 3664
rect 352101 3655 352159 3661
rect 352101 3652 352113 3655
rect 325292 3624 352113 3652
rect 325292 3612 325298 3624
rect 352101 3621 352113 3624
rect 352147 3621 352159 3655
rect 352101 3615 352159 3621
rect 352193 3655 352251 3661
rect 352193 3621 352205 3655
rect 352239 3652 352251 3655
rect 355045 3655 355103 3661
rect 355045 3652 355057 3655
rect 352239 3624 355057 3652
rect 352239 3621 352251 3624
rect 352193 3615 352251 3621
rect 355045 3621 355057 3624
rect 355091 3621 355103 3655
rect 355413 3655 355471 3661
rect 355413 3652 355425 3655
rect 355045 3615 355103 3621
rect 355152 3624 355425 3652
rect 265860 3556 320772 3584
rect 320821 3587 320879 3593
rect 265860 3544 265866 3556
rect 320821 3553 320833 3587
rect 320867 3584 320879 3587
rect 322753 3587 322811 3593
rect 322753 3584 322765 3587
rect 320867 3556 322765 3584
rect 320867 3553 320879 3556
rect 320821 3547 320879 3553
rect 322753 3553 322765 3556
rect 322799 3553 322811 3587
rect 322753 3547 322811 3553
rect 322842 3544 322848 3596
rect 322900 3584 322906 3596
rect 327074 3584 327080 3596
rect 322900 3556 327080 3584
rect 322900 3544 322906 3556
rect 327074 3544 327080 3556
rect 327132 3544 327138 3596
rect 332137 3587 332195 3593
rect 332137 3553 332149 3587
rect 332183 3584 332195 3587
rect 335357 3587 335415 3593
rect 335357 3584 335369 3587
rect 332183 3556 335369 3584
rect 332183 3553 332195 3556
rect 332137 3547 332195 3553
rect 335357 3553 335369 3556
rect 335403 3553 335415 3587
rect 335357 3547 335415 3553
rect 335909 3587 335967 3593
rect 335909 3553 335921 3587
rect 335955 3584 335967 3587
rect 355152 3584 355180 3624
rect 355413 3621 355425 3624
rect 355459 3621 355471 3655
rect 355413 3615 355471 3621
rect 355505 3655 355563 3661
rect 355505 3621 355517 3655
rect 355551 3652 355563 3655
rect 358906 3652 358912 3664
rect 355551 3624 358912 3652
rect 355551 3621 355563 3624
rect 355505 3615 355563 3621
rect 358906 3612 358912 3624
rect 358964 3612 358970 3664
rect 360930 3612 360936 3664
rect 360988 3652 360994 3664
rect 377398 3652 377404 3664
rect 360988 3624 377404 3652
rect 360988 3612 360994 3624
rect 377398 3612 377404 3624
rect 377456 3612 377462 3664
rect 400030 3612 400036 3664
rect 400088 3652 400094 3664
rect 413186 3652 413192 3664
rect 400088 3624 413192 3652
rect 400088 3612 400094 3624
rect 413186 3612 413192 3624
rect 413244 3612 413250 3664
rect 416682 3612 416688 3664
rect 416740 3652 416746 3664
rect 417528 3652 417556 3692
rect 422849 3689 422861 3692
rect 422895 3689 422907 3723
rect 422849 3683 422907 3689
rect 431865 3723 431923 3729
rect 431865 3689 431877 3723
rect 431911 3720 431923 3723
rect 441617 3723 441675 3729
rect 441617 3720 441629 3723
rect 431911 3692 441629 3720
rect 431911 3689 431923 3692
rect 431865 3683 431923 3689
rect 441617 3689 441629 3692
rect 441663 3689 441675 3723
rect 441617 3683 441675 3689
rect 416740 3624 417556 3652
rect 416740 3612 416746 3624
rect 421558 3612 421564 3664
rect 421616 3652 421622 3664
rect 425241 3655 425299 3661
rect 425241 3652 425253 3655
rect 421616 3624 425253 3652
rect 421616 3612 421622 3624
rect 425241 3621 425253 3624
rect 425287 3621 425299 3655
rect 425241 3615 425299 3621
rect 427078 3612 427084 3664
rect 427136 3652 427142 3664
rect 431126 3652 431132 3664
rect 427136 3624 431132 3652
rect 427136 3612 427142 3624
rect 431126 3612 431132 3624
rect 431184 3612 431190 3664
rect 431221 3655 431279 3661
rect 431221 3621 431233 3655
rect 431267 3652 431279 3655
rect 441709 3655 441767 3661
rect 441709 3652 441721 3655
rect 431267 3624 441721 3652
rect 431267 3621 431279 3624
rect 431221 3615 431279 3621
rect 441709 3621 441721 3624
rect 441755 3621 441767 3655
rect 441709 3615 441767 3621
rect 442350 3612 442356 3664
rect 442408 3652 442414 3664
rect 443089 3655 443147 3661
rect 443089 3652 443101 3655
rect 442408 3624 443101 3652
rect 442408 3612 442414 3624
rect 443089 3621 443101 3624
rect 443135 3621 443147 3655
rect 443089 3615 443147 3621
rect 443638 3612 443644 3664
rect 443696 3652 443702 3664
rect 446493 3655 446551 3661
rect 446493 3652 446505 3655
rect 443696 3624 446505 3652
rect 443696 3612 443702 3624
rect 446493 3621 446505 3624
rect 446539 3621 446551 3655
rect 446493 3615 446551 3621
rect 446582 3612 446588 3664
rect 446640 3652 446646 3664
rect 446784 3652 446812 3760
rect 452470 3748 452476 3760
rect 452528 3748 452534 3800
rect 456702 3748 456708 3800
rect 456760 3788 456766 3800
rect 460106 3788 460112 3800
rect 456760 3760 460112 3788
rect 456760 3748 456766 3760
rect 460106 3748 460112 3760
rect 460164 3748 460170 3800
rect 460290 3748 460296 3800
rect 460348 3788 460354 3800
rect 463234 3788 463240 3800
rect 460348 3760 463240 3788
rect 460348 3748 460354 3760
rect 463234 3748 463240 3760
rect 463292 3748 463298 3800
rect 557166 3788 557172 3800
rect 463344 3760 557172 3788
rect 456797 3723 456855 3729
rect 456797 3689 456809 3723
rect 456843 3720 456855 3723
rect 456843 3692 457392 3720
rect 456843 3689 456855 3692
rect 456797 3683 456855 3689
rect 446640 3624 446812 3652
rect 446640 3612 446646 3624
rect 449158 3612 449164 3664
rect 449216 3652 449222 3664
rect 457165 3655 457223 3661
rect 457165 3652 457177 3655
rect 449216 3624 457177 3652
rect 449216 3612 449222 3624
rect 457165 3621 457177 3624
rect 457211 3621 457223 3655
rect 457165 3615 457223 3621
rect 361850 3584 361856 3596
rect 335955 3556 355180 3584
rect 355244 3556 361856 3584
rect 335955 3553 335967 3556
rect 335909 3547 335967 3553
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 236270 3516 236276 3528
rect 16080 3488 236276 3516
rect 16080 3476 16086 3488
rect 236270 3476 236276 3488
rect 236328 3476 236334 3528
rect 258626 3476 258632 3528
rect 258684 3516 258690 3528
rect 320358 3516 320364 3528
rect 258684 3488 320364 3516
rect 258684 3476 258690 3488
rect 320358 3476 320364 3488
rect 320416 3476 320422 3528
rect 320450 3476 320456 3528
rect 320508 3516 320514 3528
rect 321186 3516 321192 3528
rect 320508 3488 321192 3516
rect 320508 3476 320514 3488
rect 321186 3476 321192 3488
rect 321244 3476 321250 3528
rect 321646 3476 321652 3528
rect 321704 3516 321710 3528
rect 355244 3516 355272 3556
rect 361850 3544 361856 3556
rect 361908 3544 361914 3596
rect 402238 3544 402244 3596
rect 402296 3584 402302 3596
rect 415670 3584 415676 3596
rect 402296 3556 415676 3584
rect 402296 3544 402302 3556
rect 415670 3544 415676 3556
rect 415728 3544 415734 3596
rect 418062 3544 418068 3596
rect 418120 3584 418126 3596
rect 457254 3584 457260 3596
rect 418120 3556 457260 3584
rect 418120 3544 418126 3556
rect 457254 3544 457260 3556
rect 457312 3544 457318 3596
rect 457364 3584 457392 3692
rect 460198 3680 460204 3732
rect 460256 3720 460262 3732
rect 460256 3692 461716 3720
rect 460256 3680 460262 3692
rect 461688 3652 461716 3692
rect 463344 3652 463372 3760
rect 557166 3748 557172 3760
rect 557224 3748 557230 3800
rect 564342 3720 564348 3732
rect 461688 3624 463372 3652
rect 463436 3692 564348 3720
rect 457364 3556 460980 3584
rect 363138 3516 363144 3528
rect 321704 3488 355272 3516
rect 355336 3488 363144 3516
rect 321704 3476 321710 3488
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 234982 3448 234988 3460
rect 14884 3420 234988 3448
rect 14884 3408 14890 3420
rect 234982 3408 234988 3420
rect 235040 3408 235046 3460
rect 255038 3408 255044 3460
rect 255096 3448 255102 3460
rect 318702 3448 318708 3460
rect 255096 3420 318708 3448
rect 255096 3408 255102 3420
rect 318702 3408 318708 3420
rect 318760 3408 318766 3460
rect 320637 3451 320695 3457
rect 320637 3417 320649 3451
rect 320683 3448 320695 3451
rect 322750 3448 322756 3460
rect 320683 3420 322756 3448
rect 320683 3417 320695 3420
rect 320637 3411 320695 3417
rect 322750 3408 322756 3420
rect 322808 3408 322814 3460
rect 324038 3408 324044 3460
rect 324096 3448 324102 3460
rect 355336 3448 355364 3488
rect 363138 3476 363144 3488
rect 363196 3476 363202 3528
rect 376757 3519 376815 3525
rect 376757 3516 376769 3519
rect 370240 3488 376769 3516
rect 324096 3420 355364 3448
rect 355413 3451 355471 3457
rect 324096 3408 324102 3420
rect 355413 3417 355425 3451
rect 355459 3448 355471 3451
rect 363598 3448 363604 3460
rect 355459 3420 363604 3448
rect 355459 3417 355471 3420
rect 355413 3411 355471 3417
rect 363598 3408 363604 3420
rect 363656 3408 363662 3460
rect 368014 3408 368020 3460
rect 368072 3448 368078 3460
rect 370240 3448 370268 3488
rect 376757 3485 376769 3488
rect 376803 3485 376815 3519
rect 376757 3479 376815 3485
rect 379974 3476 379980 3528
rect 380032 3516 380038 3528
rect 380802 3516 380808 3528
rect 380032 3488 380808 3516
rect 380032 3476 380038 3488
rect 380802 3476 380808 3488
rect 380860 3476 380866 3528
rect 381170 3476 381176 3528
rect 381228 3516 381234 3528
rect 382182 3516 382188 3528
rect 381228 3488 382188 3516
rect 381228 3476 381234 3488
rect 382182 3476 382188 3488
rect 382240 3476 382246 3528
rect 388254 3476 388260 3528
rect 388312 3516 388318 3528
rect 389082 3516 389088 3528
rect 388312 3488 389088 3516
rect 388312 3476 388318 3488
rect 389082 3476 389088 3488
rect 389140 3476 389146 3528
rect 395982 3476 395988 3528
rect 396040 3516 396046 3528
rect 401318 3516 401324 3528
rect 396040 3488 401324 3516
rect 396040 3476 396046 3488
rect 401318 3476 401324 3488
rect 401376 3476 401382 3528
rect 402790 3476 402796 3528
rect 402848 3516 402854 3528
rect 413189 3519 413247 3525
rect 413189 3516 413201 3519
rect 402848 3488 413201 3516
rect 402848 3476 402854 3488
rect 413189 3485 413201 3488
rect 413235 3485 413247 3519
rect 413189 3479 413247 3485
rect 413278 3476 413284 3528
rect 413336 3516 413342 3528
rect 414474 3516 414480 3528
rect 413336 3488 414480 3516
rect 413336 3476 413342 3488
rect 414474 3476 414480 3488
rect 414532 3476 414538 3528
rect 420822 3476 420828 3528
rect 420880 3516 420886 3528
rect 460842 3516 460848 3528
rect 420880 3488 460848 3516
rect 420880 3476 420886 3488
rect 460842 3476 460848 3488
rect 460900 3476 460906 3528
rect 460952 3516 460980 3556
rect 462222 3544 462228 3596
rect 462280 3584 462286 3596
rect 463436 3584 463464 3692
rect 564342 3680 564348 3692
rect 564400 3680 564406 3732
rect 463602 3612 463608 3664
rect 463660 3652 463666 3664
rect 566734 3652 566740 3664
rect 463660 3624 566740 3652
rect 463660 3612 463666 3624
rect 566734 3612 566740 3624
rect 566792 3612 566798 3664
rect 462280 3556 463464 3584
rect 462280 3544 462286 3556
rect 463510 3544 463516 3596
rect 463568 3584 463574 3596
rect 466089 3587 466147 3593
rect 466089 3584 466101 3587
rect 463568 3556 466101 3584
rect 463568 3544 463574 3556
rect 466089 3553 466101 3556
rect 466135 3553 466147 3587
rect 466089 3547 466147 3553
rect 466362 3544 466368 3596
rect 466420 3584 466426 3596
rect 571426 3584 571432 3596
rect 466420 3556 571432 3584
rect 466420 3544 466426 3556
rect 571426 3544 571432 3556
rect 571484 3544 571490 3596
rect 466181 3519 466239 3525
rect 466181 3516 466193 3519
rect 460952 3488 466193 3516
rect 466181 3485 466193 3488
rect 466227 3485 466239 3519
rect 466181 3479 466239 3485
rect 466270 3476 466276 3528
rect 466328 3516 466334 3528
rect 573818 3516 573824 3528
rect 466328 3488 573824 3516
rect 466328 3476 466334 3488
rect 573818 3476 573824 3488
rect 573876 3476 573882 3528
rect 368072 3420 370268 3448
rect 370317 3451 370375 3457
rect 368072 3408 368078 3420
rect 370317 3417 370329 3451
rect 370363 3448 370375 3451
rect 379698 3448 379704 3460
rect 370363 3420 379704 3448
rect 370363 3417 370375 3420
rect 370317 3411 370375 3417
rect 379698 3408 379704 3420
rect 379756 3408 379762 3460
rect 382366 3408 382372 3460
rect 382424 3448 382430 3460
rect 386598 3448 386604 3460
rect 382424 3420 386604 3448
rect 382424 3408 382430 3420
rect 386598 3408 386604 3420
rect 386656 3408 386662 3460
rect 395890 3408 395896 3460
rect 395948 3448 395954 3460
rect 402514 3448 402520 3460
rect 395948 3420 402520 3448
rect 395948 3408 395954 3420
rect 402514 3408 402520 3420
rect 402572 3408 402578 3460
rect 403618 3408 403624 3460
rect 403676 3448 403682 3460
rect 407298 3448 407304 3460
rect 403676 3420 407304 3448
rect 403676 3408 403682 3420
rect 407298 3408 407304 3420
rect 407356 3408 407362 3460
rect 422754 3448 422760 3460
rect 407408 3420 422760 3448
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 35158 3380 35164 3392
rect 29144 3352 35164 3380
rect 29144 3340 29150 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 39298 3380 39304 3392
rect 36228 3352 39304 3380
rect 36228 3340 36234 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 45465 3383 45523 3389
rect 45465 3349 45477 3383
rect 45511 3380 45523 3383
rect 45511 3352 58296 3380
rect 45511 3349 45523 3352
rect 45465 3343 45523 3349
rect 10042 3272 10048 3324
rect 10100 3312 10106 3324
rect 13078 3312 13084 3324
rect 10100 3284 13084 3312
rect 10100 3272 10106 3284
rect 13078 3272 13084 3284
rect 13136 3272 13142 3324
rect 42150 3272 42156 3324
rect 42208 3312 42214 3324
rect 57238 3312 57244 3324
rect 42208 3284 57244 3312
rect 42208 3272 42214 3284
rect 57238 3272 57244 3284
rect 57296 3272 57302 3324
rect 58268 3312 58296 3352
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 251818 3380 251824 3392
rect 71792 3352 251824 3380
rect 61378 3312 61384 3324
rect 58268 3284 61384 3312
rect 61378 3272 61384 3284
rect 61436 3272 61442 3324
rect 52822 3204 52828 3256
rect 52880 3244 52886 3256
rect 53742 3244 53748 3256
rect 52880 3216 53748 3244
rect 52880 3204 52886 3216
rect 53742 3204 53748 3216
rect 53800 3204 53806 3256
rect 54018 3204 54024 3256
rect 54076 3244 54082 3256
rect 54076 3216 59676 3244
rect 54076 3204 54082 3216
rect 43346 3136 43352 3188
rect 43404 3176 43410 3188
rect 45465 3179 45523 3185
rect 45465 3176 45477 3179
rect 43404 3148 45477 3176
rect 43404 3136 43410 3148
rect 45465 3145 45477 3148
rect 45511 3145 45523 3179
rect 45465 3139 45523 3145
rect 59648 3108 59676 3216
rect 64782 3204 64788 3256
rect 64840 3244 64846 3256
rect 71792 3244 71820 3352
rect 251818 3340 251824 3352
rect 251876 3340 251882 3392
rect 282825 3383 282883 3389
rect 282825 3349 282837 3383
rect 282871 3380 282883 3383
rect 289814 3380 289820 3392
rect 282871 3352 289820 3380
rect 282871 3349 282883 3352
rect 282825 3343 282883 3349
rect 289814 3340 289820 3352
rect 289872 3340 289878 3392
rect 299106 3340 299112 3392
rect 299164 3380 299170 3392
rect 302878 3380 302884 3392
rect 299164 3352 302884 3380
rect 299164 3340 299170 3352
rect 302878 3340 302884 3352
rect 302936 3340 302942 3392
rect 310974 3340 310980 3392
rect 311032 3380 311038 3392
rect 341429 3383 341487 3389
rect 341429 3380 341441 3383
rect 311032 3352 341441 3380
rect 311032 3340 311038 3352
rect 341429 3349 341441 3352
rect 341475 3349 341487 3383
rect 341429 3343 341487 3349
rect 341518 3340 341524 3392
rect 341576 3380 341582 3392
rect 345661 3383 345719 3389
rect 341576 3352 344416 3380
rect 341576 3340 341582 3352
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 253198 3312 253204 3324
rect 71924 3284 253204 3312
rect 71924 3272 71930 3284
rect 253198 3272 253204 3284
rect 253256 3272 253262 3324
rect 288434 3312 288440 3324
rect 276400 3284 288440 3312
rect 64840 3216 71820 3244
rect 71884 3216 74580 3244
rect 64840 3204 64846 3216
rect 61194 3136 61200 3188
rect 61252 3176 61258 3188
rect 61252 3148 67956 3176
rect 61252 3136 61258 3148
rect 66898 3108 66904 3120
rect 59648 3080 66904 3108
rect 66898 3068 66904 3080
rect 66956 3068 66962 3120
rect 67928 3108 67956 3148
rect 68278 3136 68284 3188
rect 68336 3176 68342 3188
rect 71884 3176 71912 3216
rect 68336 3148 71912 3176
rect 68336 3136 68342 3148
rect 71038 3108 71044 3120
rect 67928 3080 71044 3108
rect 71038 3068 71044 3080
rect 71096 3068 71102 3120
rect 74552 3040 74580 3216
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 84838 3244 84844 3256
rect 82832 3216 84844 3244
rect 75454 3136 75460 3188
rect 75512 3176 75518 3188
rect 79318 3176 79324 3188
rect 75512 3148 79324 3176
rect 75512 3136 75518 3148
rect 79318 3136 79324 3148
rect 79376 3136 79382 3188
rect 82630 3136 82636 3188
rect 82688 3176 82694 3188
rect 82832 3176 82860 3216
rect 84838 3204 84844 3216
rect 84896 3204 84902 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 88518 3204 88524 3256
rect 88576 3244 88582 3256
rect 89622 3244 89628 3256
rect 88576 3216 89628 3244
rect 88576 3204 88582 3216
rect 89622 3204 89628 3216
rect 89680 3204 89686 3256
rect 254578 3244 254584 3256
rect 89732 3216 254584 3244
rect 82688 3148 82860 3176
rect 82909 3179 82967 3185
rect 82688 3136 82694 3148
rect 82909 3145 82921 3179
rect 82955 3176 82967 3179
rect 89732 3176 89760 3216
rect 254578 3204 254584 3216
rect 254636 3204 254642 3256
rect 269298 3204 269304 3256
rect 269356 3244 269362 3256
rect 273257 3247 273315 3253
rect 273257 3244 273269 3247
rect 269356 3216 273269 3244
rect 269356 3204 269362 3216
rect 273257 3213 273269 3216
rect 273303 3213 273315 3247
rect 273257 3207 273315 3213
rect 255958 3176 255964 3188
rect 82955 3148 89760 3176
rect 94424 3148 255964 3176
rect 82955 3145 82967 3148
rect 82909 3139 82967 3145
rect 89714 3068 89720 3120
rect 89772 3108 89778 3120
rect 94424 3108 94452 3148
rect 255958 3136 255964 3148
rect 256016 3136 256022 3188
rect 272886 3136 272892 3188
rect 272944 3176 272950 3188
rect 276400 3176 276428 3284
rect 288434 3272 288440 3284
rect 288492 3272 288498 3324
rect 288621 3315 288679 3321
rect 288621 3281 288633 3315
rect 288667 3312 288679 3315
rect 292485 3315 292543 3321
rect 292485 3312 292497 3315
rect 288667 3284 292497 3312
rect 288667 3281 288679 3284
rect 288621 3275 288679 3281
rect 292485 3281 292497 3284
rect 292531 3281 292543 3315
rect 292485 3275 292543 3281
rect 303798 3272 303804 3324
rect 303856 3312 303862 3324
rect 344278 3312 344284 3324
rect 303856 3284 344284 3312
rect 303856 3272 303862 3284
rect 344278 3272 344284 3284
rect 344336 3272 344342 3324
rect 344388 3312 344416 3352
rect 345661 3349 345673 3383
rect 345707 3380 345719 3383
rect 352929 3383 352987 3389
rect 352929 3380 352941 3383
rect 345707 3352 352941 3380
rect 345707 3349 345719 3352
rect 345661 3343 345719 3349
rect 352929 3349 352941 3352
rect 352975 3349 352987 3383
rect 352929 3343 352987 3349
rect 353754 3340 353760 3392
rect 353812 3380 353818 3392
rect 375650 3380 375656 3392
rect 353812 3352 375656 3380
rect 353812 3340 353818 3352
rect 375650 3340 375656 3352
rect 375708 3340 375714 3392
rect 404262 3340 404268 3392
rect 404320 3380 404326 3392
rect 407408 3380 407436 3420
rect 422754 3408 422760 3420
rect 422812 3408 422818 3460
rect 424318 3408 424324 3460
rect 424376 3448 424382 3460
rect 467926 3448 467932 3460
rect 424376 3420 467932 3448
rect 424376 3408 424382 3420
rect 467926 3408 467932 3420
rect 467984 3408 467990 3460
rect 469030 3408 469036 3460
rect 469088 3448 469094 3460
rect 578602 3448 578608 3460
rect 469088 3420 578608 3448
rect 469088 3408 469094 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 404320 3352 407436 3380
rect 404320 3340 404326 3352
rect 409782 3340 409788 3392
rect 409840 3380 409846 3392
rect 433889 3383 433947 3389
rect 433889 3380 433901 3383
rect 409840 3352 433901 3380
rect 409840 3340 409846 3352
rect 433889 3349 433901 3352
rect 433935 3349 433947 3383
rect 433889 3343 433947 3349
rect 433978 3340 433984 3392
rect 434036 3380 434042 3392
rect 435818 3380 435824 3392
rect 434036 3352 435824 3380
rect 434036 3340 434042 3352
rect 435818 3340 435824 3352
rect 435876 3340 435882 3392
rect 438118 3340 438124 3392
rect 438176 3380 438182 3392
rect 446401 3383 446459 3389
rect 446401 3380 446413 3383
rect 438176 3352 446413 3380
rect 438176 3340 438182 3352
rect 446401 3349 446413 3352
rect 446447 3349 446459 3383
rect 446401 3343 446459 3349
rect 446493 3383 446551 3389
rect 446493 3349 446505 3383
rect 446539 3380 446551 3383
rect 446539 3352 510108 3380
rect 446539 3349 446551 3352
rect 446493 3343 446551 3349
rect 348418 3312 348424 3324
rect 344388 3284 348424 3312
rect 348418 3272 348424 3284
rect 348476 3272 348482 3324
rect 349062 3272 349068 3324
rect 349120 3312 349126 3324
rect 364981 3315 365039 3321
rect 364981 3312 364993 3315
rect 349120 3284 364993 3312
rect 349120 3272 349126 3284
rect 364981 3281 364993 3284
rect 365027 3281 365039 3315
rect 364981 3275 365039 3281
rect 365530 3272 365536 3324
rect 365588 3312 365594 3324
rect 369857 3315 369915 3321
rect 369857 3312 369869 3315
rect 365588 3284 369869 3312
rect 365588 3272 365594 3284
rect 369857 3281 369869 3284
rect 369903 3281 369915 3315
rect 369857 3275 369915 3281
rect 394510 3272 394516 3324
rect 394568 3312 394574 3324
rect 399018 3312 399024 3324
rect 394568 3284 399024 3312
rect 394568 3272 394574 3284
rect 399018 3272 399024 3284
rect 399076 3272 399082 3324
rect 404998 3272 405004 3324
rect 405056 3312 405062 3324
rect 416866 3312 416872 3324
rect 405056 3284 416872 3312
rect 405056 3272 405062 3284
rect 416866 3272 416872 3284
rect 416924 3272 416930 3324
rect 420178 3272 420184 3324
rect 420236 3312 420242 3324
rect 446582 3312 446588 3324
rect 420236 3284 446588 3312
rect 420236 3272 420242 3284
rect 446582 3272 446588 3284
rect 446640 3272 446646 3324
rect 446677 3315 446735 3321
rect 446677 3281 446689 3315
rect 446723 3312 446735 3315
rect 503622 3312 503628 3324
rect 446723 3284 503628 3312
rect 446723 3281 446735 3284
rect 446677 3275 446735 3281
rect 503622 3272 503628 3284
rect 503680 3272 503686 3324
rect 510080 3312 510108 3352
rect 514018 3340 514024 3392
rect 514076 3380 514082 3392
rect 517882 3380 517888 3392
rect 514076 3352 517888 3380
rect 514076 3340 514082 3352
rect 517882 3340 517888 3352
rect 517940 3340 517946 3392
rect 525058 3380 525064 3392
rect 517992 3352 525064 3380
rect 514386 3312 514392 3324
rect 510080 3284 514392 3312
rect 514386 3272 514392 3284
rect 514444 3272 514450 3324
rect 516870 3272 516876 3324
rect 516928 3312 516934 3324
rect 517992 3312 518020 3352
rect 525058 3340 525064 3352
rect 525116 3340 525122 3392
rect 527818 3340 527824 3392
rect 527876 3380 527882 3392
rect 567838 3380 567844 3392
rect 527876 3352 567844 3380
rect 527876 3340 527882 3352
rect 567838 3340 567844 3352
rect 567896 3340 567902 3392
rect 577406 3312 577412 3324
rect 516928 3284 518020 3312
rect 518084 3284 577412 3312
rect 516928 3272 516934 3284
rect 276474 3204 276480 3256
rect 276532 3244 276538 3256
rect 288526 3244 288532 3256
rect 276532 3216 288532 3244
rect 276532 3204 276538 3216
rect 288526 3204 288532 3216
rect 288584 3204 288590 3256
rect 291930 3204 291936 3256
rect 291988 3244 291994 3256
rect 316678 3244 316684 3256
rect 291988 3216 316684 3244
rect 291988 3204 291994 3216
rect 316678 3204 316684 3216
rect 316736 3204 316742 3256
rect 318058 3204 318064 3256
rect 318116 3244 318122 3256
rect 345569 3247 345627 3253
rect 345569 3244 345581 3247
rect 318116 3216 345581 3244
rect 318116 3204 318122 3216
rect 345569 3213 345581 3216
rect 345615 3213 345627 3247
rect 345569 3207 345627 3213
rect 345750 3204 345756 3256
rect 345808 3244 345814 3256
rect 349157 3247 349215 3253
rect 349157 3244 349169 3247
rect 345808 3216 349169 3244
rect 345808 3204 345814 3216
rect 349157 3213 349169 3216
rect 349203 3213 349215 3247
rect 349157 3207 349215 3213
rect 350258 3204 350264 3256
rect 350316 3244 350322 3256
rect 352377 3247 352435 3253
rect 352377 3244 352389 3247
rect 350316 3216 352389 3244
rect 350316 3204 350322 3216
rect 352377 3213 352389 3216
rect 352423 3213 352435 3247
rect 352377 3207 352435 3213
rect 352929 3247 352987 3253
rect 352929 3213 352941 3247
rect 352975 3244 352987 3247
rect 355318 3244 355324 3256
rect 352975 3216 355324 3244
rect 352975 3213 352987 3216
rect 352929 3207 352987 3213
rect 355318 3204 355324 3216
rect 355376 3204 355382 3256
rect 357342 3204 357348 3256
rect 357400 3244 357406 3256
rect 376018 3244 376024 3256
rect 357400 3216 376024 3244
rect 357400 3204 357406 3216
rect 376018 3204 376024 3216
rect 376076 3204 376082 3256
rect 394602 3204 394608 3256
rect 394660 3244 394666 3256
rect 400214 3244 400220 3256
rect 394660 3216 400220 3244
rect 394660 3204 394666 3216
rect 400214 3204 400220 3216
rect 400272 3204 400278 3256
rect 409138 3204 409144 3256
rect 409196 3244 409202 3256
rect 432322 3244 432328 3256
rect 409196 3216 432328 3244
rect 409196 3204 409202 3216
rect 432322 3204 432328 3216
rect 432380 3204 432386 3256
rect 433889 3247 433947 3253
rect 433889 3213 433901 3247
rect 433935 3244 433947 3247
rect 437014 3244 437020 3256
rect 433935 3216 437020 3244
rect 433935 3213 433947 3216
rect 433889 3207 433947 3213
rect 437014 3204 437020 3216
rect 437072 3204 437078 3256
rect 441617 3247 441675 3253
rect 441617 3213 441629 3247
rect 441663 3244 441675 3247
rect 446214 3244 446220 3256
rect 441663 3216 446220 3244
rect 441663 3213 441675 3216
rect 441617 3207 441675 3213
rect 446214 3204 446220 3216
rect 446272 3204 446278 3256
rect 446309 3247 446367 3253
rect 446309 3213 446321 3247
rect 446355 3244 446367 3247
rect 496538 3244 496544 3256
rect 446355 3216 496544 3244
rect 446355 3213 446367 3216
rect 446309 3207 446367 3213
rect 496538 3204 496544 3216
rect 496596 3204 496602 3256
rect 512638 3204 512644 3256
rect 512696 3244 512702 3256
rect 518084 3244 518112 3284
rect 577406 3272 577412 3284
rect 577464 3272 577470 3324
rect 512696 3216 518112 3244
rect 518161 3247 518219 3253
rect 512696 3204 512702 3216
rect 518161 3213 518173 3247
rect 518207 3244 518219 3247
rect 570230 3244 570236 3256
rect 518207 3216 570236 3244
rect 518207 3213 518219 3216
rect 518161 3207 518219 3213
rect 570230 3204 570236 3216
rect 570288 3204 570294 3256
rect 272944 3148 276428 3176
rect 272944 3136 272950 3148
rect 277670 3136 277676 3188
rect 277728 3176 277734 3188
rect 290458 3176 290464 3188
rect 277728 3148 290464 3176
rect 277728 3136 277734 3148
rect 290458 3136 290464 3148
rect 290516 3136 290522 3188
rect 309778 3136 309784 3188
rect 309836 3176 309842 3188
rect 335998 3176 336004 3188
rect 309836 3148 336004 3176
rect 309836 3136 309842 3148
rect 335998 3136 336004 3148
rect 336056 3136 336062 3188
rect 336093 3179 336151 3185
rect 336093 3145 336105 3179
rect 336139 3176 336151 3179
rect 340601 3179 340659 3185
rect 340601 3176 340613 3179
rect 336139 3148 340613 3176
rect 336139 3145 336151 3148
rect 336093 3139 336151 3145
rect 340601 3145 340613 3148
rect 340647 3145 340659 3179
rect 340601 3139 340659 3145
rect 340690 3136 340696 3188
rect 340748 3176 340754 3188
rect 345661 3179 345719 3185
rect 345661 3176 345673 3179
rect 340748 3148 345673 3176
rect 340748 3136 340754 3148
rect 345661 3145 345673 3148
rect 345707 3145 345719 3179
rect 345661 3139 345719 3145
rect 346670 3136 346676 3188
rect 346728 3176 346734 3188
rect 370498 3176 370504 3188
rect 346728 3148 370504 3176
rect 346728 3136 346734 3148
rect 370498 3136 370504 3148
rect 370556 3136 370562 3188
rect 407022 3136 407028 3188
rect 407080 3176 407086 3188
rect 429930 3176 429936 3188
rect 407080 3148 429936 3176
rect 407080 3136 407086 3148
rect 429930 3136 429936 3148
rect 429988 3136 429994 3188
rect 431218 3136 431224 3188
rect 431276 3176 431282 3188
rect 431276 3148 477632 3176
rect 431276 3136 431282 3148
rect 89772 3080 94452 3108
rect 89772 3068 89778 3080
rect 94498 3068 94504 3120
rect 94556 3108 94562 3120
rect 95142 3108 95148 3120
rect 94556 3080 95148 3108
rect 94556 3068 94562 3080
rect 95142 3068 95148 3080
rect 95200 3068 95206 3120
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 98086 3068 98092 3120
rect 98144 3108 98150 3120
rect 99190 3108 99196 3120
rect 98144 3080 99196 3108
rect 98144 3068 98150 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 101582 3068 101588 3120
rect 101640 3108 101646 3120
rect 102042 3108 102048 3120
rect 101640 3080 102048 3108
rect 101640 3068 101646 3080
rect 102042 3068 102048 3080
rect 102100 3068 102106 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 105170 3068 105176 3120
rect 105228 3108 105234 3120
rect 106182 3108 106188 3120
rect 105228 3080 106188 3108
rect 105228 3068 105234 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107470 3108 107476 3120
rect 106424 3080 107476 3108
rect 106424 3068 106430 3080
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 257338 3108 257344 3120
rect 108316 3080 257344 3108
rect 77938 3040 77944 3052
rect 74552 3012 77944 3040
rect 77938 3000 77944 3012
rect 77996 3000 78002 3052
rect 93302 3000 93308 3052
rect 93360 3040 93366 3052
rect 102594 3040 102600 3052
rect 93360 3012 102600 3040
rect 93360 3000 93366 3012
rect 102594 3000 102600 3012
rect 102652 3000 102658 3052
rect 79042 2932 79048 2984
rect 79100 2972 79106 2984
rect 82909 2975 82967 2981
rect 82909 2972 82921 2975
rect 79100 2944 82921 2972
rect 79100 2932 79106 2944
rect 82909 2941 82921 2944
rect 82955 2941 82967 2975
rect 82909 2935 82967 2941
rect 86126 2932 86132 2984
rect 86184 2972 86190 2984
rect 93857 2975 93915 2981
rect 93857 2972 93869 2975
rect 86184 2944 93869 2972
rect 86184 2932 86190 2944
rect 93857 2941 93869 2944
rect 93903 2941 93915 2975
rect 93857 2935 93915 2941
rect 96890 2932 96896 2984
rect 96948 2972 96954 2984
rect 108316 2972 108344 3080
rect 257338 3068 257344 3080
rect 257396 3068 257402 3120
rect 295518 3068 295524 3120
rect 295576 3108 295582 3120
rect 319438 3108 319444 3120
rect 295576 3080 319444 3108
rect 295576 3068 295582 3080
rect 319438 3068 319444 3080
rect 319496 3068 319502 3120
rect 322753 3111 322811 3117
rect 322753 3077 322765 3111
rect 322799 3108 322811 3111
rect 327718 3108 327724 3120
rect 322799 3080 327724 3108
rect 322799 3077 322811 3080
rect 322753 3071 322811 3077
rect 327718 3068 327724 3080
rect 327776 3068 327782 3120
rect 328822 3068 328828 3120
rect 328880 3108 328886 3120
rect 355505 3111 355563 3117
rect 355505 3108 355517 3111
rect 328880 3080 355517 3108
rect 328880 3068 328886 3080
rect 355505 3077 355517 3080
rect 355551 3077 355563 3111
rect 355505 3071 355563 3077
rect 355597 3111 355655 3117
rect 355597 3077 355609 3111
rect 355643 3108 355655 3111
rect 359458 3108 359464 3120
rect 355643 3080 359464 3108
rect 355643 3077 355655 3080
rect 355597 3071 355655 3077
rect 359458 3068 359464 3080
rect 359516 3068 359522 3120
rect 364981 3111 365039 3117
rect 364981 3077 364993 3111
rect 365027 3108 365039 3111
rect 372982 3108 372988 3120
rect 365027 3080 372988 3108
rect 365027 3077 365039 3080
rect 364981 3071 365039 3077
rect 372982 3068 372988 3080
rect 373040 3068 373046 3120
rect 405642 3068 405648 3120
rect 405700 3108 405706 3120
rect 426342 3108 426348 3120
rect 405700 3080 426348 3108
rect 405700 3068 405706 3080
rect 426342 3068 426348 3080
rect 426400 3068 426406 3120
rect 428458 3068 428464 3120
rect 428516 3108 428522 3120
rect 475102 3108 475108 3120
rect 428516 3080 475108 3108
rect 428516 3068 428522 3080
rect 475102 3068 475108 3080
rect 475160 3068 475166 3120
rect 475378 3068 475384 3120
rect 475436 3108 475442 3120
rect 477494 3108 477500 3120
rect 475436 3080 477500 3108
rect 475436 3068 475442 3080
rect 477494 3068 477500 3080
rect 477552 3068 477558 3120
rect 477604 3108 477632 3148
rect 505738 3136 505744 3188
rect 505796 3176 505802 3188
rect 563146 3176 563152 3188
rect 505796 3148 563152 3176
rect 505796 3136 505802 3148
rect 563146 3136 563152 3148
rect 563204 3136 563210 3188
rect 482278 3108 482284 3120
rect 477604 3080 482284 3108
rect 482278 3068 482284 3080
rect 482336 3068 482342 3120
rect 524966 3068 524972 3120
rect 525024 3108 525030 3120
rect 560754 3108 560760 3120
rect 525024 3080 560760 3108
rect 525024 3068 525030 3080
rect 560754 3068 560760 3080
rect 560812 3068 560818 3120
rect 258718 3040 258724 3052
rect 96948 2944 108344 2972
rect 108408 3012 258724 3040
rect 96948 2932 96954 2944
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 108408 2904 108436 3012
rect 258718 3000 258724 3012
rect 258776 3000 258782 3052
rect 273257 3043 273315 3049
rect 273257 3009 273269 3043
rect 273303 3040 273315 3043
rect 282825 3043 282883 3049
rect 282825 3040 282837 3043
rect 273303 3012 282837 3040
rect 273303 3009 273315 3012
rect 273257 3003 273315 3009
rect 282825 3009 282837 3012
rect 282871 3009 282883 3043
rect 282825 3003 282883 3009
rect 293126 3000 293132 3052
rect 293184 3040 293190 3052
rect 312538 3040 312544 3052
rect 293184 3012 312544 3040
rect 293184 3000 293190 3012
rect 312538 3000 312544 3012
rect 312596 3000 312602 3052
rect 315758 3000 315764 3052
rect 315816 3040 315822 3052
rect 323302 3040 323308 3052
rect 315816 3012 323308 3040
rect 315816 3000 315822 3012
rect 323302 3000 323308 3012
rect 323360 3000 323366 3052
rect 327626 3000 327632 3052
rect 327684 3040 327690 3052
rect 335909 3043 335967 3049
rect 335909 3040 335921 3043
rect 327684 3012 335921 3040
rect 327684 3000 327690 3012
rect 335909 3009 335921 3012
rect 335955 3009 335967 3043
rect 335909 3003 335967 3009
rect 336182 3000 336188 3052
rect 336240 3040 336246 3052
rect 360289 3043 360347 3049
rect 360289 3040 360301 3043
rect 336240 3012 360301 3040
rect 336240 3000 336246 3012
rect 360289 3009 360301 3012
rect 360335 3009 360347 3043
rect 360289 3003 360347 3009
rect 360396 3012 364472 3040
rect 112346 2932 112352 2984
rect 112404 2972 112410 2984
rect 113082 2972 113088 2984
rect 112404 2944 113088 2972
rect 112404 2932 112410 2944
rect 113082 2932 113088 2944
rect 113140 2932 113146 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 115934 2932 115940 2984
rect 115992 2972 115998 2984
rect 116946 2972 116952 2984
rect 115992 2944 116952 2972
rect 115992 2932 115998 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 119430 2932 119436 2984
rect 119488 2972 119494 2984
rect 119982 2972 119988 2984
rect 119488 2944 119988 2972
rect 119488 2932 119494 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 258810 2972 258816 2984
rect 121472 2944 258816 2972
rect 104032 2876 108436 2904
rect 104032 2864 104038 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 121472 2904 121500 2944
rect 258810 2932 258816 2944
rect 258868 2932 258874 2984
rect 316954 2932 316960 2984
rect 317012 2972 317018 2984
rect 335541 2975 335599 2981
rect 335541 2972 335553 2975
rect 317012 2944 335553 2972
rect 317012 2932 317018 2944
rect 335541 2941 335553 2944
rect 335587 2941 335599 2975
rect 335541 2935 335599 2941
rect 335998 2932 336004 2984
rect 336056 2972 336062 2984
rect 341337 2975 341395 2981
rect 341337 2972 341349 2975
rect 336056 2944 341349 2972
rect 336056 2932 336062 2944
rect 341337 2941 341349 2944
rect 341383 2941 341395 2975
rect 341337 2935 341395 2941
rect 341429 2975 341487 2981
rect 341429 2941 341441 2975
rect 341475 2972 341487 2975
rect 352466 2972 352472 2984
rect 341475 2944 352472 2972
rect 341475 2941 341487 2944
rect 341429 2935 341487 2941
rect 352466 2932 352472 2944
rect 352524 2932 352530 2984
rect 352558 2932 352564 2984
rect 352616 2972 352622 2984
rect 360396 2972 360424 3012
rect 352616 2944 360424 2972
rect 360473 2975 360531 2981
rect 352616 2932 352622 2944
rect 360473 2941 360485 2975
rect 360519 2972 360531 2975
rect 364444 2972 364472 3012
rect 364518 3000 364524 3052
rect 364576 3040 364582 3052
rect 365530 3040 365536 3052
rect 364576 3012 365536 3040
rect 364576 3000 364582 3012
rect 365530 3000 365536 3012
rect 365588 3000 365594 3052
rect 376386 3000 376392 3052
rect 376444 3040 376450 3052
rect 381630 3040 381636 3052
rect 376444 3012 381636 3040
rect 376444 3000 376450 3012
rect 381630 3000 381636 3012
rect 381688 3000 381694 3052
rect 406378 3000 406384 3052
rect 406436 3040 406442 3052
rect 410886 3040 410892 3052
rect 406436 3012 410892 3040
rect 406436 3000 406442 3012
rect 410886 3000 410892 3012
rect 410944 3000 410950 3052
rect 413189 3043 413247 3049
rect 413189 3009 413201 3043
rect 413235 3040 413247 3043
rect 420362 3040 420368 3052
rect 413235 3012 420368 3040
rect 413235 3009 413247 3012
rect 413189 3003 413247 3009
rect 420362 3000 420368 3012
rect 420420 3000 420426 3052
rect 422941 3043 422999 3049
rect 422941 3009 422953 3043
rect 422987 3040 422999 3043
rect 431221 3043 431279 3049
rect 431221 3040 431233 3043
rect 422987 3012 431233 3040
rect 422987 3009 422999 3012
rect 422941 3003 422999 3009
rect 431221 3009 431233 3012
rect 431267 3009 431279 3043
rect 431221 3003 431279 3009
rect 431310 3000 431316 3052
rect 431368 3040 431374 3052
rect 459646 3040 459652 3052
rect 431368 3012 459652 3040
rect 431368 3000 431374 3012
rect 459646 3000 459652 3012
rect 459704 3000 459710 3052
rect 461581 3043 461639 3049
rect 461581 3009 461593 3043
rect 461627 3040 461639 3043
rect 489362 3040 489368 3052
rect 461627 3012 489368 3040
rect 461627 3009 461639 3012
rect 461581 3003 461639 3009
rect 489362 3000 489368 3012
rect 489420 3000 489426 3052
rect 509878 3000 509884 3052
rect 509936 3040 509942 3052
rect 518161 3043 518219 3049
rect 518161 3040 518173 3043
rect 509936 3012 518173 3040
rect 509936 3000 509942 3012
rect 518161 3009 518173 3012
rect 518207 3009 518219 3043
rect 518161 3003 518219 3009
rect 523678 3000 523684 3052
rect 523736 3040 523742 3052
rect 553578 3040 553584 3052
rect 523736 3012 553584 3040
rect 523736 3000 523742 3012
rect 553578 3000 553584 3012
rect 553636 3000 553642 3052
rect 374086 2972 374092 2984
rect 360519 2944 362356 2972
rect 364444 2944 374092 2972
rect 360519 2941 360531 2944
rect 360473 2935 360531 2941
rect 260098 2904 260104 2916
rect 111208 2876 121500 2904
rect 121564 2876 260104 2904
rect 111208 2864 111214 2876
rect 93857 2839 93915 2845
rect 93857 2805 93869 2839
rect 93903 2836 93915 2839
rect 95878 2836 95884 2848
rect 93903 2808 95884 2836
rect 93903 2805 93915 2808
rect 93857 2799 93915 2805
rect 95878 2796 95884 2808
rect 95936 2796 95942 2848
rect 114738 2796 114744 2848
rect 114796 2836 114802 2848
rect 121564 2836 121592 2876
rect 260098 2864 260104 2876
rect 260156 2864 260162 2916
rect 275278 2864 275284 2916
rect 275336 2904 275342 2916
rect 275922 2904 275928 2916
rect 275336 2876 275928 2904
rect 275336 2864 275342 2876
rect 275922 2864 275928 2876
rect 275980 2864 275986 2916
rect 319254 2864 319260 2916
rect 319312 2904 319318 2916
rect 326338 2904 326344 2916
rect 319312 2876 326344 2904
rect 319312 2864 319318 2876
rect 326338 2864 326344 2876
rect 326396 2864 326402 2916
rect 335906 2864 335912 2916
rect 335964 2904 335970 2916
rect 336182 2904 336188 2916
rect 335964 2876 336188 2904
rect 335964 2864 335970 2876
rect 336182 2864 336188 2876
rect 336240 2864 336246 2916
rect 340785 2907 340843 2913
rect 340785 2873 340797 2907
rect 340831 2904 340843 2907
rect 340966 2904 340972 2916
rect 340831 2876 340972 2904
rect 340831 2873 340843 2876
rect 340785 2867 340843 2873
rect 340966 2864 340972 2876
rect 341024 2864 341030 2916
rect 344278 2864 344284 2916
rect 344336 2904 344342 2916
rect 352009 2907 352067 2913
rect 352009 2904 352021 2907
rect 344336 2876 352021 2904
rect 344336 2864 344342 2876
rect 352009 2873 352021 2876
rect 352055 2873 352067 2907
rect 352009 2867 352067 2873
rect 352101 2907 352159 2913
rect 352101 2873 352113 2907
rect 352147 2904 352159 2907
rect 355597 2907 355655 2913
rect 355597 2904 355609 2907
rect 352147 2876 355609 2904
rect 352147 2873 352159 2876
rect 352101 2867 352159 2873
rect 355597 2873 355609 2876
rect 355643 2873 355655 2907
rect 356698 2904 356704 2916
rect 355597 2867 355655 2873
rect 355704 2876 356704 2904
rect 114796 2808 121592 2836
rect 114796 2796 114802 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 261478 2836 261484 2848
rect 121880 2808 261484 2836
rect 121880 2796 121886 2808
rect 261478 2796 261484 2808
rect 261536 2796 261542 2848
rect 330018 2796 330024 2848
rect 330076 2836 330082 2848
rect 335449 2839 335507 2845
rect 335449 2836 335461 2839
rect 330076 2808 335461 2836
rect 330076 2796 330082 2808
rect 335449 2805 335461 2808
rect 335495 2805 335507 2839
rect 335449 2799 335507 2805
rect 335541 2839 335599 2845
rect 335541 2805 335553 2839
rect 335587 2836 335599 2839
rect 341245 2839 341303 2845
rect 341245 2836 341257 2839
rect 335587 2808 341257 2836
rect 335587 2805 335599 2808
rect 335541 2799 335599 2805
rect 341245 2805 341257 2808
rect 341291 2805 341303 2839
rect 341245 2799 341303 2805
rect 341337 2839 341395 2845
rect 341337 2805 341349 2839
rect 341383 2836 341395 2839
rect 344370 2836 344376 2848
rect 341383 2808 344376 2836
rect 341383 2805 341395 2808
rect 341337 2799 341395 2805
rect 344370 2796 344376 2808
rect 344428 2796 344434 2848
rect 345569 2839 345627 2845
rect 345569 2805 345581 2839
rect 345615 2836 345627 2839
rect 355704 2836 355732 2876
rect 356698 2864 356704 2876
rect 356756 2864 356762 2916
rect 362328 2904 362356 2944
rect 374086 2932 374092 2944
rect 374144 2932 374150 2984
rect 398190 2932 398196 2984
rect 398248 2972 398254 2984
rect 404906 2972 404912 2984
rect 398248 2944 404912 2972
rect 398248 2932 398254 2944
rect 404906 2932 404912 2944
rect 404964 2932 404970 2984
rect 417418 2932 417424 2984
rect 417476 2972 417482 2984
rect 428734 2972 428740 2984
rect 417476 2944 428740 2972
rect 417476 2932 417482 2944
rect 428734 2932 428740 2944
rect 428792 2932 428798 2984
rect 429838 2932 429844 2984
rect 429896 2972 429902 2984
rect 448974 2972 448980 2984
rect 429896 2944 448980 2972
rect 429896 2932 429902 2944
rect 448974 2932 448980 2944
rect 449032 2932 449038 2984
rect 451829 2975 451887 2981
rect 451829 2972 451841 2975
rect 451292 2944 451841 2972
rect 367278 2904 367284 2916
rect 362328 2876 367284 2904
rect 367278 2864 367284 2876
rect 367336 2864 367342 2916
rect 385862 2864 385868 2916
rect 385920 2904 385926 2916
rect 387058 2904 387064 2916
rect 385920 2876 387064 2904
rect 385920 2864 385926 2876
rect 387058 2864 387064 2876
rect 387116 2864 387122 2916
rect 416590 2864 416596 2916
rect 416648 2904 416654 2916
rect 422941 2907 422999 2913
rect 422941 2904 422953 2907
rect 416648 2876 422953 2904
rect 416648 2864 416654 2876
rect 422941 2873 422953 2876
rect 422987 2873 422999 2907
rect 451185 2907 451243 2913
rect 451185 2904 451197 2907
rect 422941 2867 422999 2873
rect 446324 2876 451197 2904
rect 345615 2808 355732 2836
rect 345615 2805 345627 2808
rect 345569 2799 345627 2805
rect 356146 2796 356152 2848
rect 356204 2836 356210 2848
rect 356790 2836 356796 2848
rect 356204 2808 356796 2836
rect 356204 2796 356210 2808
rect 356790 2796 356796 2808
rect 356848 2796 356854 2848
rect 357066 2796 357072 2848
rect 357124 2836 357130 2848
rect 375834 2836 375840 2848
rect 357124 2808 375840 2836
rect 357124 2796 357130 2808
rect 375834 2796 375840 2808
rect 375892 2796 375898 2848
rect 388438 2836 388444 2848
rect 387076 2808 388444 2836
rect 387076 2780 387104 2808
rect 388438 2796 388444 2808
rect 388496 2796 388502 2848
rect 422849 2839 422907 2845
rect 422849 2805 422861 2839
rect 422895 2836 422907 2839
rect 431865 2839 431923 2845
rect 431865 2836 431877 2839
rect 422895 2808 431877 2836
rect 422895 2805 422907 2808
rect 422849 2799 422907 2805
rect 431865 2805 431877 2808
rect 431911 2805 431923 2839
rect 431865 2799 431923 2805
rect 439498 2796 439504 2848
rect 439556 2836 439562 2848
rect 446324 2836 446352 2876
rect 451185 2873 451197 2876
rect 451231 2873 451243 2907
rect 451185 2867 451243 2873
rect 439556 2808 446352 2836
rect 446401 2839 446459 2845
rect 439556 2796 439562 2808
rect 446401 2805 446413 2839
rect 446447 2836 446459 2839
rect 451292 2836 451320 2944
rect 451829 2941 451841 2944
rect 451875 2941 451887 2975
rect 451829 2935 451887 2941
rect 451921 2975 451979 2981
rect 451921 2941 451933 2975
rect 451967 2972 451979 2975
rect 481082 2972 481088 2984
rect 451967 2944 481088 2972
rect 451967 2941 451979 2944
rect 451921 2935 451979 2941
rect 481082 2932 481088 2944
rect 481140 2932 481146 2984
rect 521010 2932 521016 2984
rect 521068 2972 521074 2984
rect 546494 2972 546500 2984
rect 521068 2944 546500 2972
rect 521068 2932 521074 2944
rect 546494 2932 546500 2944
rect 546552 2932 546558 2984
rect 451369 2907 451427 2913
rect 451369 2873 451381 2907
rect 451415 2904 451427 2907
rect 456797 2907 456855 2913
rect 456797 2904 456809 2907
rect 451415 2876 456809 2904
rect 451415 2873 451427 2876
rect 451369 2867 451427 2873
rect 456797 2873 456809 2876
rect 456843 2873 456855 2907
rect 456797 2867 456855 2873
rect 457165 2907 457223 2913
rect 457165 2873 457177 2907
rect 457211 2904 457223 2907
rect 461581 2907 461639 2913
rect 461581 2904 461593 2907
rect 457211 2876 461593 2904
rect 457211 2873 457223 2876
rect 457165 2867 457223 2873
rect 461581 2873 461593 2876
rect 461627 2873 461639 2907
rect 461581 2867 461639 2873
rect 466365 2907 466423 2913
rect 466365 2873 466377 2907
rect 466411 2904 466423 2907
rect 473906 2904 473912 2916
rect 466411 2876 473912 2904
rect 466411 2873 466423 2876
rect 466365 2867 466423 2873
rect 473906 2864 473912 2876
rect 473964 2864 473970 2916
rect 520918 2864 520924 2916
rect 520976 2904 520982 2916
rect 539318 2904 539324 2916
rect 520976 2876 539324 2904
rect 520976 2864 520982 2876
rect 539318 2864 539324 2876
rect 539376 2864 539382 2916
rect 446447 2808 451320 2836
rect 451829 2839 451887 2845
rect 446447 2805 446459 2808
rect 446401 2799 446459 2805
rect 451829 2805 451841 2839
rect 451875 2836 451887 2839
rect 466822 2836 466828 2848
rect 451875 2808 466828 2836
rect 451875 2805 451887 2808
rect 451829 2799 451887 2805
rect 466822 2796 466828 2808
rect 466880 2796 466886 2848
rect 518158 2796 518164 2848
rect 518216 2836 518222 2848
rect 532234 2836 532240 2848
rect 518216 2808 532240 2836
rect 518216 2796 518222 2808
rect 532234 2796 532240 2808
rect 532292 2796 532298 2848
rect 355505 2771 355563 2777
rect 355505 2737 355517 2771
rect 355551 2768 355563 2771
rect 362218 2768 362224 2780
rect 355551 2740 362224 2768
rect 355551 2737 355563 2740
rect 355505 2731 355563 2737
rect 362218 2728 362224 2740
rect 362276 2728 362282 2780
rect 387058 2728 387064 2780
rect 387116 2728 387122 2780
rect 261018 1096 261024 1148
rect 261076 1136 261082 1148
rect 264609 1139 264667 1145
rect 264609 1136 264621 1139
rect 261076 1108 264621 1136
rect 261076 1096 261082 1108
rect 264609 1105 264621 1108
rect 264655 1105 264667 1139
rect 264609 1099 264667 1105
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 164694 552 164700 604
rect 164752 592 164758 604
rect 165522 592 165528 604
rect 164752 564 165528 592
rect 164752 552 164758 564
rect 165522 552 165528 564
rect 165580 552 165586 604
rect 165890 552 165896 604
rect 165948 592 165954 604
rect 166902 592 166908 604
rect 165948 564 166908 592
rect 165948 552 165954 564
rect 166902 552 166908 564
rect 166960 552 166966 604
rect 169386 552 169392 604
rect 169444 592 169450 604
rect 169662 592 169668 604
rect 169444 564 169668 592
rect 169444 552 169450 564
rect 169662 552 169668 564
rect 169720 552 169726 604
rect 182542 552 182548 604
rect 182600 592 182606 604
rect 183462 592 183468 604
rect 182600 564 183468 592
rect 182600 552 182606 564
rect 183462 552 183468 564
rect 183520 552 183526 604
rect 183738 552 183744 604
rect 183796 592 183802 604
rect 184750 592 184756 604
rect 183796 564 184756 592
rect 183796 552 183802 564
rect 184750 552 184756 564
rect 184808 552 184814 604
rect 187234 552 187240 604
rect 187292 592 187298 604
rect 187602 592 187608 604
rect 187292 564 187608 592
rect 187292 552 187298 564
rect 187602 552 187608 564
rect 187660 552 187666 604
rect 189626 552 189632 604
rect 189684 592 189690 604
rect 190362 592 190368 604
rect 189684 564 190368 592
rect 189684 552 189690 564
rect 190362 552 190368 564
rect 190420 552 190426 604
rect 281258 552 281264 604
rect 281316 592 281322 604
rect 281442 592 281448 604
rect 281316 564 281448 592
rect 281316 552 281322 564
rect 281442 552 281448 564
rect 281500 552 281506 604
rect 389450 592 389456 604
rect 389411 564 389456 592
rect 389450 552 389456 564
rect 389508 552 389514 604
rect 393590 552 393596 604
rect 393648 592 393654 604
rect 394234 592 394240 604
rect 393648 564 394240 592
rect 393648 552 393654 564
rect 394234 552 394240 564
rect 394292 552 394298 604
rect 397454 552 397460 604
rect 397512 592 397518 604
rect 397822 592 397828 604
rect 397512 564 397828 592
rect 397512 552 397518 564
rect 397822 552 397828 564
rect 397880 552 397886 604
rect 405918 552 405924 604
rect 405976 592 405982 604
rect 406102 592 406108 604
rect 405976 564 406108 592
rect 405976 552 405982 564
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 463694 552 463700 604
rect 463752 592 463758 604
rect 464430 592 464436 604
rect 463752 564 464436 592
rect 463752 552 463758 564
rect 464430 552 464436 564
rect 464488 552 464494 604
rect 469214 552 469220 604
rect 469272 592 469278 604
rect 470318 592 470324 604
rect 469272 564 470324 592
rect 469272 552 469278 564
rect 470318 552 470324 564
rect 470376 552 470382 604
rect 471514 592 471520 604
rect 471475 564 471520 592
rect 471514 552 471520 564
rect 471572 552 471578 604
<< via1 >>
rect 202788 700952 202840 701004
rect 358820 700952 358872 701004
rect 170312 700884 170364 700936
rect 362960 700884 363012 700936
rect 328368 700816 328420 700868
rect 527180 700816 527232 700868
rect 329748 700748 329800 700800
rect 543464 700748 543516 700800
rect 154120 700680 154172 700732
rect 367100 700680 367152 700732
rect 137836 700612 137888 700664
rect 364340 700612 364392 700664
rect 105452 700544 105504 700596
rect 368480 700544 368532 700596
rect 89168 700476 89220 700528
rect 374000 700476 374052 700528
rect 72976 700408 73028 700460
rect 371240 700408 371292 700460
rect 40500 700340 40552 700392
rect 375380 700340 375432 700392
rect 24308 700272 24360 700324
rect 379520 700272 379572 700324
rect 218980 700204 219032 700256
rect 360200 700204 360252 700256
rect 336648 700136 336700 700188
rect 478512 700136 478564 700188
rect 335268 700068 335320 700120
rect 462320 700068 462372 700120
rect 235172 700000 235224 700052
rect 356060 700000 356112 700052
rect 267648 699932 267700 699984
rect 351920 699932 351972 699984
rect 283840 699864 283892 699916
rect 354680 699864 354732 699916
rect 343548 699796 343600 699848
rect 413652 699796 413704 699848
rect 340788 699728 340840 699780
rect 397460 699728 397512 699780
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 332508 699660 332560 699712
rect 346400 699660 346452 699712
rect 347780 699660 347832 699712
rect 348792 699660 348844 699712
rect 321468 696940 321520 696992
rect 580172 696940 580224 696992
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 364616 687760 364668 687812
rect 365168 687760 365220 687812
rect 324228 685856 324280 685908
rect 580172 685856 580224 685908
rect 364616 685788 364668 685840
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 382280 681708 382332 681760
rect 364524 676243 364576 676252
rect 364524 676209 364533 676243
rect 364533 676209 364567 676243
rect 364567 676209 364576 676243
rect 364524 676200 364576 676209
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 320088 673480 320140 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 386420 667904 386472 667956
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 383660 652740 383712 652792
rect 315948 650020 316000 650072
rect 580172 650020 580224 650072
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 317328 638936 317380 638988
rect 580172 638936 580224 638988
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 313188 626560 313240 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 387800 623772 387852 623824
rect 364616 618196 364668 618248
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3424 609968 3476 610020
rect 391940 609968 391992 610020
rect 364524 608651 364576 608660
rect 364524 608617 364533 608651
rect 364533 608617 364567 608651
rect 364567 608617 364576 608651
rect 364524 608608 364576 608617
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 309048 603100 309100 603152
rect 580172 603100 580224 603152
rect 429568 601672 429620 601724
rect 559288 601672 559340 601724
rect 364616 598927 364668 598936
rect 364616 598893 364625 598927
rect 364625 598893 364659 598927
rect 364659 598893 364668 598927
rect 364616 598884 364668 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 390560 594804 390612 594856
rect 311808 592016 311860 592068
rect 580172 592016 580224 592068
rect 364708 589296 364760 589348
rect 429660 589296 429712 589348
rect 559380 589296 559432 589348
rect 344468 584672 344520 584724
rect 364708 584672 364760 584724
rect 300768 584604 300820 584656
rect 350816 584604 350868 584656
rect 338212 584536 338264 584588
rect 429660 584536 429712 584588
rect 331864 584468 331916 584520
rect 494244 584468 494296 584520
rect 325516 584400 325568 584452
rect 559380 584400 559432 584452
rect 304540 583652 304592 583704
rect 471336 583652 471388 583704
rect 298192 583584 298244 583636
rect 471244 583584 471296 583636
rect 256056 583516 256108 583568
rect 580632 583516 580684 583568
rect 251824 583448 251876 583500
rect 580540 583448 580592 583500
rect 245568 583380 245620 583432
rect 580356 583380 580408 583432
rect 4712 583312 4764 583364
rect 399208 583312 399260 583364
rect 5448 583244 5500 583296
rect 405556 583244 405608 583296
rect 10324 583176 10376 583228
rect 411904 583176 411956 583228
rect 6276 583108 6328 583160
rect 409788 583108 409840 583160
rect 3148 583040 3200 583092
rect 407672 583040 407724 583092
rect 13084 582972 13136 583024
rect 418160 582972 418212 583024
rect 14464 582904 14516 582956
rect 424508 582904 424560 582956
rect 3240 582836 3292 582888
rect 414020 582836 414072 582888
rect 5356 582768 5408 582820
rect 422392 582768 422444 582820
rect 15844 582700 15896 582752
rect 437112 582700 437164 582752
rect 4068 582632 4120 582684
rect 430856 582632 430908 582684
rect 5264 582564 5316 582616
rect 432972 582564 433024 582616
rect 3884 582496 3936 582548
rect 434996 582496 435048 582548
rect 5172 582428 5224 582480
rect 445576 582428 445628 582480
rect 3700 582360 3752 582412
rect 443460 582360 443512 582412
rect 302424 581476 302476 581528
rect 469588 581476 469640 581528
rect 296076 581408 296128 581460
rect 469680 581408 469732 581460
rect 289728 581340 289780 581392
rect 469772 581340 469824 581392
rect 287612 581272 287664 581324
rect 470508 581272 470560 581324
rect 283472 581204 283524 581256
rect 470416 581204 470468 581256
rect 281356 581136 281408 581188
rect 470232 581136 470284 581188
rect 275008 581068 275060 581120
rect 470140 581068 470192 581120
rect 264520 581000 264572 581052
rect 580080 581000 580132 581052
rect 268660 580320 268712 580372
rect 469956 580320 470008 580372
rect 262404 580252 262456 580304
rect 469864 580252 469916 580304
rect 306564 580184 306616 580236
rect 580172 580184 580224 580236
rect 6644 580116 6696 580168
rect 395068 580116 395120 580168
rect 6552 580048 6604 580100
rect 397092 580048 397144 580100
rect 6460 579980 6512 580032
rect 400956 579980 401008 580032
rect 6368 579912 6420 579964
rect 403164 579912 403216 579964
rect 3792 579844 3844 579896
rect 438860 579844 438912 579896
rect 4988 579776 5040 579828
rect 451556 579776 451608 579828
rect 4896 579708 4948 579760
rect 458272 579708 458324 579760
rect 6184 579640 6236 579692
rect 464252 579640 464304 579692
rect 271144 579368 271196 579420
rect 247960 579343 248012 579352
rect 247960 579309 247969 579343
rect 247969 579309 248003 579343
rect 248003 579309 248012 579343
rect 247960 579300 248012 579309
rect 254216 579343 254268 579352
rect 254216 579309 254225 579343
rect 254225 579309 254259 579343
rect 254259 579309 254268 579343
rect 254216 579300 254268 579309
rect 258448 579300 258500 579352
rect 260656 579300 260708 579352
rect 266912 579300 266964 579352
rect 273168 579300 273220 579352
rect 277308 579300 277360 579352
rect 279608 579300 279660 579352
rect 285772 579300 285824 579352
rect 292120 579343 292172 579352
rect 292120 579309 292129 579343
rect 292129 579309 292163 579343
rect 292163 579309 292172 579343
rect 292120 579300 292172 579309
rect 415676 579343 415728 579352
rect 415676 579309 415685 579343
rect 415685 579309 415719 579343
rect 415719 579309 415728 579343
rect 415676 579300 415728 579309
rect 428372 579343 428424 579352
rect 428372 579309 428381 579343
rect 428381 579309 428415 579343
rect 428415 579309 428424 579343
rect 428372 579300 428424 579309
rect 441068 579343 441120 579352
rect 441068 579309 441077 579343
rect 441077 579309 441111 579343
rect 441111 579309 441120 579343
rect 441068 579300 441120 579309
rect 453580 579343 453632 579352
rect 453580 579309 453589 579343
rect 453589 579309 453623 579343
rect 453623 579309 453632 579343
rect 453580 579300 453632 579309
rect 455788 579343 455840 579352
rect 455788 579309 455797 579343
rect 455797 579309 455831 579343
rect 455831 579309 455840 579343
rect 455788 579300 455840 579309
rect 470324 579232 470376 579284
rect 470048 579164 470100 579216
rect 579804 579096 579856 579148
rect 579988 579028 580040 579080
rect 579896 578960 579948 579012
rect 580080 578892 580132 578944
rect 580908 578824 580960 578876
rect 580724 578756 580776 578808
rect 580816 578688 580868 578740
rect 580448 578620 580500 578672
rect 580264 578552 580316 578604
rect 3332 578484 3384 578536
rect 3976 578416 4028 578468
rect 3608 578348 3660 578400
rect 3424 578280 3476 578332
rect 3516 578212 3568 578264
rect 3056 567332 3108 567384
rect 6644 567332 6696 567384
rect 469588 557472 469640 557524
rect 579712 557472 579764 557524
rect 2780 553052 2832 553104
rect 4712 553052 4764 553104
rect 471336 546388 471388 546440
rect 579712 546388 579764 546440
rect 3056 538636 3108 538688
rect 6552 538636 6604 538688
rect 469680 510552 469732 510604
rect 579712 510552 579764 510604
rect 3056 510212 3108 510264
rect 6460 510212 6512 510264
rect 471244 499468 471296 499520
rect 579712 499468 579764 499520
rect 2780 496680 2832 496732
rect 5448 496680 5500 496732
rect 2964 481108 3016 481160
rect 6368 481108 6420 481160
rect 469772 463632 469824 463684
rect 579712 463632 579764 463684
rect 470508 440172 470560 440224
rect 579804 440172 579856 440224
rect 3148 438812 3200 438864
rect 10324 438812 10376 438864
rect 3148 424056 3200 424108
rect 6276 424056 6328 424108
rect 470416 416712 470468 416764
rect 579804 416712 579856 416764
rect 470324 405628 470376 405680
rect 579804 405628 579856 405680
rect 470232 393252 470284 393304
rect 579804 393252 579856 393304
rect 3240 380808 3292 380860
rect 13084 380808 13136 380860
rect 470140 346332 470192 346384
rect 579988 346332 580040 346384
rect 244648 338648 244700 338700
rect 348516 338648 348568 338700
rect 316132 338104 316184 338156
rect 316316 338104 316368 338156
rect 318800 338104 318852 338156
rect 319812 338104 319864 338156
rect 337384 338104 337436 338156
rect 337752 338104 337804 338156
rect 340328 338104 340380 338156
rect 340696 338104 340748 338156
rect 372068 338104 372120 338156
rect 460848 338104 460900 338156
rect 71044 338036 71096 338088
rect 254952 338036 255004 338088
rect 314660 338036 314712 338088
rect 315396 338036 315448 338088
rect 354404 338036 354456 338088
rect 358084 338036 358136 338088
rect 371516 338036 371568 338088
rect 406292 338036 406344 338088
rect 417424 338036 417476 338088
rect 419080 338036 419132 338088
rect 431408 338036 431460 338088
rect 435732 338036 435784 338088
rect 499580 338036 499632 338088
rect 66904 337968 66956 338020
rect 252008 337968 252060 338020
rect 306196 337968 306248 338020
rect 355876 337968 355928 338020
rect 364248 337968 364300 338020
rect 379336 337968 379388 338020
rect 61384 337900 61436 337952
rect 247592 337900 247644 337952
rect 303160 337900 303212 337952
rect 352932 337900 352984 337952
rect 355324 337900 355376 337952
rect 370044 337900 370096 337952
rect 371148 337900 371200 337952
rect 382280 337968 382332 338020
rect 397460 337968 397512 338020
rect 403624 337968 403676 338020
rect 414664 337968 414716 338020
rect 429752 337968 429804 338020
rect 437204 337968 437256 338020
rect 442356 337968 442408 338020
rect 446036 337968 446088 338020
rect 454776 337968 454828 338020
rect 461676 337968 461728 338020
rect 525064 337968 525116 338020
rect 400404 337900 400456 337952
rect 413284 337900 413336 337952
rect 413652 337900 413704 337952
rect 420184 337900 420236 337952
rect 420552 337900 420604 337952
rect 57244 337832 57296 337884
rect 247132 337832 247184 337884
rect 290464 337832 290516 337884
rect 347044 337832 347096 337884
rect 348424 337832 348476 337884
rect 365628 337832 365680 337884
rect 50344 337764 50396 337816
rect 244188 337764 244240 337816
rect 259644 337764 259696 337816
rect 260104 337764 260156 337816
rect 288256 337764 288308 337816
rect 351920 337764 351972 337816
rect 362868 337764 362920 337816
rect 378876 337832 378928 337884
rect 388444 337832 388496 337884
rect 389180 337832 389232 337884
rect 404820 337832 404872 337884
rect 39304 337696 39356 337748
rect 57980 337696 58032 337748
rect 67548 337696 67600 337748
rect 77300 337696 77352 337748
rect 86868 337696 86920 337748
rect 95240 337696 95292 337748
rect 104808 337696 104860 337748
rect 114560 337696 114612 337748
rect 124128 337696 124180 337748
rect 133880 337696 133932 337748
rect 143448 337696 143500 337748
rect 153200 337696 153252 337748
rect 162768 337696 162820 337748
rect 172520 337696 172572 337748
rect 182088 337696 182140 337748
rect 191840 337696 191892 337748
rect 201408 337696 201460 337748
rect 211160 337696 211212 337748
rect 220728 337696 220780 337748
rect 32404 337628 32456 337680
rect 230664 337628 230716 337680
rect 231124 337628 231176 337680
rect 254584 337696 254636 337748
rect 262312 337696 262364 337748
rect 307760 337696 307812 337748
rect 317328 337696 317380 337748
rect 356704 337696 356756 337748
rect 360752 337696 360804 337748
rect 377404 337764 377456 337816
rect 404360 337764 404412 337816
rect 416136 337764 416188 337816
rect 416688 337764 416740 337816
rect 417608 337832 417660 337884
rect 455604 337900 455656 337952
rect 458732 337900 458784 337952
rect 459376 337900 459428 337952
rect 467104 337900 467156 337952
rect 467748 337900 467800 337952
rect 468024 337900 468076 337952
rect 469128 337900 469180 337952
rect 527824 337900 527876 337952
rect 420276 337764 420328 337816
rect 422024 337764 422076 337816
rect 438124 337764 438176 337816
rect 438676 337764 438728 337816
rect 255964 337628 256016 337680
rect 260104 337628 260156 337680
rect 277032 337628 277084 337680
rect 285588 337628 285640 337680
rect 336096 337628 336148 337680
rect 344560 337628 344612 337680
rect 349988 337628 350040 337680
rect 35164 337560 35216 337612
rect 241704 337560 241756 337612
rect 261392 337560 261444 337612
rect 279976 337560 280028 337612
rect 281448 337560 281500 337612
rect 345572 337560 345624 337612
rect 345756 337560 345808 337612
rect 350172 337560 350224 337612
rect 28264 337492 28316 337544
rect 220820 337492 220872 337544
rect 221004 337492 221056 337544
rect 237840 337492 237892 337544
rect 253204 337492 253256 337544
rect 259368 337492 259420 337544
rect 19984 337424 20036 337476
rect 234344 337424 234396 337476
rect 238300 337424 238352 337476
rect 258816 337424 258868 337476
rect 275560 337492 275612 337544
rect 275928 337492 275980 337544
rect 13084 337356 13136 337408
rect 220820 337356 220872 337408
rect 221004 337356 221056 337408
rect 233516 337356 233568 337408
rect 233884 337356 233936 337408
rect 241244 337356 241296 337408
rect 250444 337356 250496 337408
rect 253480 337356 253532 337408
rect 257344 337356 257396 337408
rect 269672 337424 269724 337476
rect 271788 337424 271840 337476
rect 341616 337492 341668 337544
rect 342720 337492 342772 337544
rect 344284 337492 344336 337544
rect 354864 337628 354916 337680
rect 358728 337628 358780 337680
rect 375932 337696 375984 337748
rect 380164 337696 380216 337748
rect 381360 337696 381412 337748
rect 381544 337696 381596 337748
rect 382832 337696 382884 337748
rect 384948 337696 385000 337748
rect 388168 337696 388220 337748
rect 399484 337696 399536 337748
rect 400128 337696 400180 337748
rect 402428 337696 402480 337748
rect 402888 337696 402940 337748
rect 403348 337696 403400 337748
rect 380808 337628 380860 337680
rect 384304 337628 384356 337680
rect 387708 337628 387760 337680
rect 398932 337628 398984 337680
rect 406384 337628 406436 337680
rect 410248 337696 410300 337748
rect 411076 337696 411128 337748
rect 414204 337696 414256 337748
rect 415308 337696 415360 337748
rect 415584 337696 415636 337748
rect 416504 337696 416556 337748
rect 417056 337696 417108 337748
rect 417976 337696 418028 337748
rect 425428 337696 425480 337748
rect 428464 337696 428516 337748
rect 429384 337696 429436 337748
rect 430488 337696 430540 337748
rect 411260 337628 411312 337680
rect 412364 337628 412416 337680
rect 351184 337560 351236 337612
rect 367008 337560 367060 337612
rect 351828 337492 351880 337544
rect 266728 337356 266780 337408
rect 269028 337356 269080 337408
rect 344100 337424 344152 337476
rect 347504 337424 347556 337476
rect 349068 337424 349120 337476
rect 373908 337492 373960 337544
rect 383292 337560 383344 337612
rect 398012 337560 398064 337612
rect 399484 337560 399536 337612
rect 407304 337560 407356 337612
rect 427084 337628 427136 337680
rect 432328 337696 432380 337748
rect 433248 337696 433300 337748
rect 433708 337696 433760 337748
rect 434628 337696 434680 337748
rect 435180 337696 435232 337748
rect 436008 337696 436060 337748
rect 436652 337696 436704 337748
rect 437388 337696 437440 337748
rect 437664 337696 437716 337748
rect 438768 337696 438820 337748
rect 439136 337696 439188 337748
rect 440148 337696 440200 337748
rect 440608 337764 440660 337816
rect 441528 337764 441580 337816
rect 441620 337764 441672 337816
rect 443644 337764 443696 337816
rect 444564 337764 444616 337816
rect 445668 337764 445720 337816
rect 448980 337764 449032 337816
rect 424692 337560 424744 337612
rect 426440 337560 426492 337612
rect 430856 337628 430908 337680
rect 431868 337628 431920 337680
rect 434720 337628 434772 337680
rect 435916 337628 435968 337680
rect 436192 337628 436244 337680
rect 437296 337628 437348 337680
rect 428372 337560 428424 337612
rect 431224 337560 431276 337612
rect 431316 337560 431368 337612
rect 375288 337492 375340 337544
rect 383752 337492 383804 337544
rect 405832 337492 405884 337544
rect 79324 337288 79376 337340
rect 260840 337288 260892 337340
rect 132500 337220 132552 337272
rect 142068 337220 142120 337272
rect 151820 337220 151872 337272
rect 161388 337220 161440 337272
rect 171140 337220 171192 337272
rect 180708 337220 180760 337272
rect 190460 337220 190512 337272
rect 200028 337220 200080 337272
rect 209780 337220 209832 337272
rect 219348 337220 219400 337272
rect 221004 337263 221056 337272
rect 221004 337229 221013 337263
rect 221013 337229 221047 337263
rect 221047 337229 221056 337263
rect 221004 337220 221056 337229
rect 234620 337220 234672 337272
rect 257896 337220 257948 337272
rect 258724 337220 258776 337272
rect 272616 337288 272668 337340
rect 272800 337288 272852 337340
rect 271328 337220 271380 337272
rect 84844 337152 84896 337204
rect 263784 337152 263836 337204
rect 297916 337152 297968 337204
rect 77944 336948 77996 337000
rect 100668 337084 100720 337136
rect 271144 337084 271196 337136
rect 309784 337288 309836 337340
rect 316040 337288 316092 337340
rect 316868 337288 316920 337340
rect 317420 337288 317472 337340
rect 318340 337288 318392 337340
rect 318892 337288 318944 337340
rect 319260 337288 319312 337340
rect 320180 337288 320232 337340
rect 320732 337288 320784 337340
rect 361764 337288 361816 337340
rect 312544 337220 312596 337272
rect 341800 337220 341852 337272
rect 348976 337220 349028 337272
rect 359464 337220 359516 337272
rect 363696 337220 363748 337272
rect 374460 337424 374512 337476
rect 381820 337424 381872 337476
rect 387064 337424 387116 337476
rect 388720 337424 388772 337476
rect 397000 337424 397052 337476
rect 405924 337424 405976 337476
rect 421196 337424 421248 337476
rect 369768 337356 369820 337408
rect 382188 337356 382240 337408
rect 386696 337356 386748 337408
rect 400956 337356 401008 337408
rect 402244 337356 402296 337408
rect 407764 337356 407816 337408
rect 409144 337356 409196 337408
rect 427912 337492 427964 337544
rect 442080 337628 442132 337680
rect 442908 337628 442960 337680
rect 443552 337628 443604 337680
rect 444288 337628 444340 337680
rect 445024 337628 445076 337680
rect 445576 337628 445628 337680
rect 446496 337628 446548 337680
rect 447048 337628 447100 337680
rect 448244 337628 448296 337680
rect 448428 337628 448480 337680
rect 449900 337628 449952 337680
rect 451004 337628 451056 337680
rect 452844 337764 452896 337816
rect 453764 337764 453816 337816
rect 454316 337764 454368 337816
rect 455236 337764 455288 337816
rect 455788 337764 455840 337816
rect 456616 337764 456668 337816
rect 457720 337764 457772 337816
rect 523684 337832 523736 337884
rect 521016 337764 521068 337816
rect 506480 337696 506532 337748
rect 518164 337628 518216 337680
rect 440240 337492 440292 337544
rect 442264 337560 442316 337612
rect 449164 337560 449216 337612
rect 450452 337560 450504 337612
rect 451188 337560 451240 337612
rect 451372 337560 451424 337612
rect 452476 337560 452528 337612
rect 453304 337560 453356 337612
rect 453948 337560 454000 337612
rect 433984 337424 434036 337476
rect 434260 337424 434312 337476
rect 439596 337424 439648 337476
rect 447508 337492 447560 337544
rect 448428 337492 448480 337544
rect 456800 337492 456852 337544
rect 458088 337492 458140 337544
rect 520924 337560 520976 337612
rect 516784 337492 516836 337544
rect 443092 337424 443144 337476
rect 514024 337424 514076 337476
rect 426440 337356 426492 337408
rect 429844 337356 429896 337408
rect 509240 337356 509292 337408
rect 366916 337288 366968 337340
rect 380348 337288 380400 337340
rect 398472 337288 398524 337340
rect 408776 337288 408828 337340
rect 409236 337288 409288 337340
rect 372988 337220 373040 337272
rect 421012 337288 421064 337340
rect 423496 337220 423548 337272
rect 460296 337220 460348 337272
rect 463884 337288 463936 337340
rect 465080 337288 465132 337340
rect 466368 337288 466420 337340
rect 470600 337288 470652 337340
rect 470692 337288 470744 337340
rect 529204 337288 529256 337340
rect 463608 337220 463660 337272
rect 469496 337220 469548 337272
rect 530584 337220 530636 337272
rect 314200 337152 314252 337204
rect 321468 337152 321520 337204
rect 312728 337084 312780 337136
rect 316684 337084 316736 337136
rect 342904 337152 342956 337204
rect 355968 337152 356020 337204
rect 401876 337152 401928 337204
rect 416964 337152 417016 337204
rect 423956 337152 424008 337204
rect 432788 337152 432840 337204
rect 492680 337152 492732 337204
rect 509240 337152 509292 337204
rect 510620 337152 510672 337204
rect 335268 337084 335320 337136
rect 95884 337016 95936 337068
rect 265256 337016 265308 337068
rect 366640 337084 366692 337136
rect 369124 337084 369176 337136
rect 371056 337084 371108 337136
rect 415124 337084 415176 337136
rect 421564 337084 421616 337136
rect 367652 337016 367704 337068
rect 393596 337016 393648 337068
rect 397460 337016 397512 337068
rect 107568 336948 107620 337000
rect 274088 336948 274140 337000
rect 319444 336948 319496 337000
rect 102784 336880 102836 336932
rect 268200 336880 268252 336932
rect 333244 336880 333296 336932
rect 338764 336880 338816 336932
rect 118608 336812 118660 336864
rect 278504 336812 278556 336864
rect 327724 336812 327776 336864
rect 340788 336880 340840 336932
rect 125508 336744 125560 336796
rect 281172 336744 281224 336796
rect 340236 336744 340288 336796
rect 249064 336676 249116 336728
rect 250536 336676 250588 336728
rect 251824 336676 251876 336728
rect 256424 336676 256476 336728
rect 262864 336676 262916 336728
rect 263048 336676 263100 336728
rect 284392 336719 284444 336728
rect 284392 336685 284401 336719
rect 284401 336685 284435 336719
rect 284435 336685 284444 336719
rect 284392 336676 284444 336685
rect 288992 336676 289044 336728
rect 327632 336676 327684 336728
rect 337384 336719 337436 336728
rect 337384 336685 337393 336719
rect 337393 336685 337427 336719
rect 337427 336685 337436 336719
rect 337384 336676 337436 336685
rect 340328 336676 340380 336728
rect 343088 336744 343140 336796
rect 344376 336812 344428 336864
rect 345572 336744 345624 336796
rect 353392 336948 353444 337000
rect 369584 336948 369636 337000
rect 378048 336948 378100 337000
rect 385224 336948 385276 337000
rect 412732 336948 412784 337000
rect 413836 336948 413888 337000
rect 345940 336880 345992 336932
rect 360292 336880 360344 336932
rect 380808 336880 380860 336932
rect 386236 336880 386288 336932
rect 392124 336880 392176 336932
rect 393596 336880 393648 336932
rect 401416 336880 401468 336932
rect 405004 336880 405056 336932
rect 409052 336880 409104 336932
rect 433524 337084 433576 337136
rect 485780 337084 485832 337136
rect 426900 337016 426952 337068
rect 477592 337016 477644 337068
rect 475384 336948 475436 337000
rect 466552 336880 466604 336932
rect 470508 336880 470560 336932
rect 357348 336812 357400 336864
rect 362224 336812 362276 336864
rect 365168 336812 365220 336864
rect 381636 336812 381688 336864
rect 384764 336812 384816 336864
rect 396080 336812 396132 336864
rect 398104 336812 398156 336864
rect 420000 336812 420052 336864
rect 420736 336812 420788 336864
rect 424968 336812 425020 336864
rect 439504 336812 439556 336864
rect 451832 336812 451884 336864
rect 459192 336812 459244 336864
rect 460204 336812 460256 336864
rect 460388 336812 460440 336864
rect 460756 336812 460808 336864
rect 469220 336812 469272 336864
rect 351460 336744 351512 336796
rect 352564 336744 352616 336796
rect 357808 336744 357860 336796
rect 363604 336744 363656 336796
rect 364708 336744 364760 336796
rect 370504 336744 370556 336796
rect 372528 336744 372580 336796
rect 376024 336744 376076 336796
rect 376944 336744 376996 336796
rect 377680 336744 377732 336796
rect 378416 336744 378468 336796
rect 395068 336744 395120 336796
rect 395988 336744 396040 336796
rect 396540 336744 396592 336796
rect 398196 336744 398248 336796
rect 418528 336744 418580 336796
rect 419448 336744 419500 336796
rect 419540 336744 419592 336796
rect 420828 336744 420880 336796
rect 421472 336744 421524 336796
rect 422208 336744 422260 336796
rect 422484 336744 422536 336796
rect 424324 336744 424376 336796
rect 424416 336744 424468 336796
rect 457260 336744 457312 336796
rect 457996 336744 458048 336796
rect 458272 336744 458324 336796
rect 459468 336744 459520 336796
rect 459744 336744 459796 336796
rect 460848 336744 460900 336796
rect 461216 336744 461268 336796
rect 462136 336744 462188 336796
rect 462688 336744 462740 336796
rect 463516 336744 463568 336796
rect 464160 336744 464212 336796
rect 464988 336744 465040 336796
rect 465080 336744 465132 336796
rect 509884 336812 509936 336864
rect 424968 336676 425020 336728
rect 505744 336744 505796 336796
rect 247224 336404 247276 336456
rect 248144 336404 248196 336456
rect 251456 335792 251508 335844
rect 252468 335792 252520 335844
rect 236184 335656 236236 335708
rect 237012 335656 237064 335708
rect 302240 335656 302292 335708
rect 302700 335656 302752 335708
rect 332692 335656 332744 335708
rect 333428 335656 333480 335708
rect 334072 335656 334124 335708
rect 334900 335656 334952 335708
rect 390652 335656 390704 335708
rect 236092 335588 236144 335640
rect 236552 335588 236604 335640
rect 241612 335588 241664 335640
rect 242348 335588 242400 335640
rect 260932 335588 260984 335640
rect 261484 335588 261536 335640
rect 263692 335588 263744 335640
rect 264428 335588 264480 335640
rect 265072 335588 265124 335640
rect 265900 335588 265952 335640
rect 266452 335588 266504 335640
rect 267372 335588 267424 335640
rect 280252 335588 280304 335640
rect 280620 335588 280672 335640
rect 281540 335588 281592 335640
rect 282092 335588 282144 335640
rect 283012 335588 283064 335640
rect 283564 335588 283616 335640
rect 285680 335588 285732 335640
rect 285956 335588 286008 335640
rect 286048 335588 286100 335640
rect 286600 335588 286652 335640
rect 287060 335588 287112 335640
rect 287980 335588 288032 335640
rect 288440 335588 288492 335640
rect 289452 335588 289504 335640
rect 292764 335588 292816 335640
rect 293316 335588 293368 335640
rect 298284 335588 298336 335640
rect 298652 335588 298704 335640
rect 300860 335588 300912 335640
rect 301228 335588 301280 335640
rect 303620 335588 303672 335640
rect 304172 335588 304224 335640
rect 305000 335588 305052 335640
rect 305644 335588 305696 335640
rect 307760 335588 307812 335640
rect 308588 335588 308640 335640
rect 309140 335588 309192 335640
rect 310060 335588 310112 335640
rect 321652 335588 321704 335640
rect 322204 335588 322256 335640
rect 329840 335588 329892 335640
rect 330116 335588 330168 335640
rect 332600 335588 332652 335640
rect 333060 335588 333112 335640
rect 333980 335588 334032 335640
rect 334532 335588 334584 335640
rect 335360 335588 335412 335640
rect 336004 335588 336056 335640
rect 338120 335588 338172 335640
rect 338948 335588 339000 335640
rect 361672 335588 361724 335640
rect 362316 335588 362368 335640
rect 363052 335588 363104 335640
rect 363788 335588 363840 335640
rect 367284 335588 367336 335640
rect 367928 335588 367980 335640
rect 372620 335588 372672 335640
rect 373264 335588 373316 335640
rect 390652 335452 390704 335504
rect 265256 335291 265308 335300
rect 265256 335257 265265 335291
rect 265265 335257 265299 335291
rect 265299 335257 265308 335291
rect 265256 335248 265308 335257
rect 284484 335180 284536 335232
rect 248512 334908 248564 334960
rect 249524 334908 249576 334960
rect 278780 334772 278832 334824
rect 278964 334772 279016 334824
rect 302608 334704 302660 334756
rect 303068 334704 303120 334756
rect 258172 334568 258224 334620
rect 258540 334568 258592 334620
rect 234988 334500 235040 334552
rect 235632 334500 235684 334552
rect 336740 334500 336792 334552
rect 336924 334500 336976 334552
rect 250628 334432 250680 334484
rect 271236 334296 271288 334348
rect 272708 334296 272760 334348
rect 247868 333956 247920 334008
rect 248604 333956 248656 334008
rect 325976 333276 326028 333328
rect 326528 333276 326580 333328
rect 374092 333140 374144 333192
rect 374736 333140 374788 333192
rect 356152 332800 356204 332852
rect 356612 332800 356664 332852
rect 284668 332528 284720 332580
rect 285128 332528 285180 332580
rect 331220 332120 331272 332172
rect 331496 332120 331548 332172
rect 242992 332052 243044 332104
rect 243452 332052 243504 332104
rect 310520 332052 310572 332104
rect 311532 332052 311584 332104
rect 331312 331712 331364 331764
rect 331956 331712 332008 331764
rect 299572 331304 299624 331356
rect 328552 331304 328604 331356
rect 329012 331304 329064 331356
rect 259644 331168 259696 331220
rect 259828 331168 259880 331220
rect 336832 331236 336884 331288
rect 341156 331168 341208 331220
rect 341340 331168 341392 331220
rect 360292 331168 360344 331220
rect 360476 331168 360528 331220
rect 389272 331168 389324 331220
rect 389456 331168 389508 331220
rect 336832 331100 336884 331152
rect 299572 331032 299624 331084
rect 306472 331032 306524 331084
rect 306656 331032 306708 331084
rect 299480 330964 299532 331016
rect 299664 330964 299716 331016
rect 301136 330488 301188 330540
rect 301688 330488 301740 330540
rect 284300 329536 284352 329588
rect 284576 329536 284628 329588
rect 270776 328491 270828 328500
rect 270776 328457 270785 328491
rect 270785 328457 270819 328491
rect 270819 328457 270828 328491
rect 270776 328448 270828 328457
rect 272248 328491 272300 328500
rect 272248 328457 272257 328491
rect 272257 328457 272291 328491
rect 272291 328457 272300 328491
rect 272248 328448 272300 328457
rect 278872 328448 278924 328500
rect 279056 328448 279108 328500
rect 303896 328448 303948 328500
rect 304632 328448 304684 328500
rect 323308 328448 323360 328500
rect 323676 328448 323728 328500
rect 324688 328448 324740 328500
rect 325148 328448 325200 328500
rect 330208 328448 330260 328500
rect 330484 328448 330536 328500
rect 259828 328423 259880 328432
rect 259828 328389 259837 328423
rect 259837 328389 259871 328423
rect 259871 328389 259880 328423
rect 259828 328380 259880 328389
rect 295524 328380 295576 328432
rect 295708 328380 295760 328432
rect 296812 328380 296864 328432
rect 296996 328380 297048 328432
rect 302608 328423 302660 328432
rect 302608 328389 302617 328423
rect 302617 328389 302651 328423
rect 302651 328389 302660 328423
rect 302608 328380 302660 328389
rect 337384 328423 337436 328432
rect 337384 328389 337393 328423
rect 337393 328389 337427 328423
rect 337427 328389 337436 328423
rect 337384 328380 337436 328389
rect 341340 328423 341392 328432
rect 341340 328389 341349 328423
rect 341349 328389 341383 328423
rect 341383 328389 341392 328423
rect 341340 328380 341392 328389
rect 389456 328423 389508 328432
rect 389456 328389 389465 328423
rect 389465 328389 389499 328423
rect 389499 328389 389508 328423
rect 389456 328380 389508 328389
rect 470600 328423 470652 328432
rect 470600 328389 470609 328423
rect 470609 328389 470643 328423
rect 470643 328389 470652 328423
rect 470600 328380 470652 328389
rect 250168 327131 250220 327140
rect 250168 327097 250177 327131
rect 250177 327097 250211 327131
rect 250211 327097 250220 327131
rect 250168 327088 250220 327097
rect 327264 327131 327316 327140
rect 327264 327097 327273 327131
rect 327273 327097 327307 327131
rect 327307 327097 327316 327131
rect 327264 327088 327316 327097
rect 273628 327020 273680 327072
rect 284668 327020 284720 327072
rect 284760 327020 284812 327072
rect 286048 327020 286100 327072
rect 330116 327063 330168 327072
rect 330116 327029 330125 327063
rect 330125 327029 330159 327063
rect 330159 327029 330168 327063
rect 330116 327020 330168 327029
rect 357624 326476 357676 326528
rect 357900 326476 357952 326528
rect 358636 325728 358688 325780
rect 358728 325728 358780 325780
rect 262680 325660 262732 325712
rect 262864 325660 262916 325712
rect 265256 325703 265308 325712
rect 265256 325669 265265 325703
rect 265265 325669 265299 325703
rect 265299 325669 265308 325703
rect 265256 325660 265308 325669
rect 463700 325660 463752 325712
rect 463884 325660 463936 325712
rect 358544 325592 358596 325644
rect 358636 325592 358688 325644
rect 3332 324232 3384 324284
rect 14464 324232 14516 324284
rect 470048 322872 470100 322924
rect 579988 322872 580040 322924
rect 236460 321691 236512 321700
rect 236460 321657 236469 321691
rect 236469 321657 236503 321691
rect 236503 321657 236512 321691
rect 236460 321648 236512 321657
rect 244464 321580 244516 321632
rect 310796 321580 310848 321632
rect 337384 321623 337436 321632
rect 337384 321589 337393 321623
rect 337393 321589 337427 321623
rect 337427 321589 337436 321623
rect 337384 321580 337436 321589
rect 375840 321580 375892 321632
rect 377128 321580 377180 321632
rect 244372 321512 244424 321564
rect 273536 321555 273588 321564
rect 273536 321521 273545 321555
rect 273545 321521 273579 321555
rect 273579 321521 273588 321555
rect 273536 321512 273588 321521
rect 310888 321444 310940 321496
rect 375932 321376 375984 321428
rect 377220 321376 377272 321428
rect 359188 318860 359240 318912
rect 362316 318860 362368 318912
rect 236460 318835 236512 318844
rect 236460 318801 236469 318835
rect 236469 318801 236503 318835
rect 236503 318801 236512 318835
rect 236460 318792 236512 318801
rect 259920 318792 259972 318844
rect 299848 318792 299900 318844
rect 300216 318792 300268 318844
rect 302608 318835 302660 318844
rect 302608 318801 302617 318835
rect 302617 318801 302651 318835
rect 302651 318801 302660 318835
rect 302608 318792 302660 318801
rect 330208 318792 330260 318844
rect 337384 318835 337436 318844
rect 337384 318801 337393 318835
rect 337393 318801 337427 318835
rect 337427 318801 337436 318835
rect 337384 318792 337436 318801
rect 339776 318835 339828 318844
rect 339776 318801 339785 318835
rect 339785 318801 339819 318835
rect 339819 318801 339828 318835
rect 339776 318792 339828 318801
rect 341432 318792 341484 318844
rect 359096 318792 359148 318844
rect 362224 318792 362276 318844
rect 389548 318792 389600 318844
rect 424600 318792 424652 318844
rect 424692 318792 424744 318844
rect 470600 318835 470652 318844
rect 470600 318801 470609 318835
rect 470609 318801 470643 318835
rect 470643 318801 470652 318835
rect 470600 318792 470652 318801
rect 372712 318767 372764 318776
rect 372712 318733 372721 318767
rect 372721 318733 372755 318767
rect 372755 318733 372764 318767
rect 372712 318724 372764 318733
rect 288992 318588 289044 318640
rect 285956 317543 286008 317552
rect 285956 317509 285965 317543
rect 285965 317509 285999 317543
rect 285999 317509 286008 317543
rect 285956 317500 286008 317509
rect 306748 317475 306800 317484
rect 306748 317441 306757 317475
rect 306757 317441 306791 317475
rect 306791 317441 306800 317475
rect 306748 317432 306800 317441
rect 236276 317364 236328 317416
rect 236460 317364 236512 317416
rect 250168 317407 250220 317416
rect 250168 317373 250177 317407
rect 250177 317373 250211 317407
rect 250211 317373 250220 317407
rect 250168 317364 250220 317373
rect 251548 317407 251600 317416
rect 251548 317373 251557 317407
rect 251557 317373 251591 317407
rect 251591 317373 251600 317407
rect 251548 317364 251600 317373
rect 266636 317364 266688 317416
rect 266728 317364 266780 317416
rect 267740 317364 267792 317416
rect 267832 317364 267884 317416
rect 273260 317364 273312 317416
rect 273536 317364 273588 317416
rect 299848 317364 299900 317416
rect 325976 317364 326028 317416
rect 421196 317407 421248 317416
rect 421196 317373 421205 317407
rect 421205 317373 421239 317407
rect 421239 317373 421248 317407
rect 421196 317364 421248 317373
rect 245844 316004 245896 316056
rect 246120 316004 246172 316056
rect 265164 316004 265216 316056
rect 265348 316004 265400 316056
rect 301136 316004 301188 316056
rect 301320 316004 301372 316056
rect 306748 316047 306800 316056
rect 306748 316013 306757 316047
rect 306757 316013 306791 316047
rect 306791 316013 306800 316047
rect 306748 316004 306800 316013
rect 357440 316004 357492 316056
rect 357624 316004 357676 316056
rect 244372 315936 244424 315988
rect 244556 315800 244608 315852
rect 290096 313259 290148 313268
rect 290096 313225 290105 313259
rect 290105 313225 290139 313259
rect 290139 313225 290148 313259
rect 290096 313216 290148 313225
rect 239036 311856 239088 311908
rect 239220 311856 239272 311908
rect 284668 311856 284720 311908
rect 285956 311899 286008 311908
rect 285956 311865 285965 311899
rect 285965 311865 285999 311899
rect 285999 311865 286008 311899
rect 285956 311856 286008 311865
rect 302608 311924 302660 311976
rect 310888 311967 310940 311976
rect 310888 311933 310897 311967
rect 310897 311933 310931 311967
rect 310931 311933 310940 311967
rect 310888 311924 310940 311933
rect 323308 311924 323360 311976
rect 323216 311856 323268 311908
rect 337200 311856 337252 311908
rect 337384 311856 337436 311908
rect 341248 311856 341300 311908
rect 341432 311856 341484 311908
rect 360200 311856 360252 311908
rect 360568 311856 360620 311908
rect 424140 311856 424192 311908
rect 424600 311856 424652 311908
rect 302516 311788 302568 311840
rect 339684 311788 339736 311840
rect 339868 311788 339920 311840
rect 291476 309136 291528 309188
rect 291568 309136 291620 309188
rect 372712 309179 372764 309188
rect 372712 309145 372721 309179
rect 372721 309145 372755 309179
rect 372755 309145 372764 309179
rect 372712 309136 372764 309145
rect 389364 309136 389416 309188
rect 389548 309136 389600 309188
rect 239128 309111 239180 309120
rect 239128 309077 239137 309111
rect 239137 309077 239171 309111
rect 239171 309077 239180 309111
rect 239128 309068 239180 309077
rect 327172 309068 327224 309120
rect 327264 309068 327316 309120
rect 339868 309111 339920 309120
rect 339868 309077 339877 309111
rect 339877 309077 339911 309111
rect 339911 309077 339920 309111
rect 339868 309068 339920 309077
rect 341248 309068 341300 309120
rect 360200 309068 360252 309120
rect 360292 309068 360344 309120
rect 367008 309111 367060 309120
rect 367008 309077 367017 309111
rect 367017 309077 367051 309111
rect 367051 309077 367060 309111
rect 367008 309068 367060 309077
rect 470600 309111 470652 309120
rect 470600 309077 470609 309111
rect 470609 309077 470643 309111
rect 470643 309077 470652 309111
rect 470600 309068 470652 309077
rect 389364 309000 389416 309052
rect 2780 308796 2832 308848
rect 5356 308796 5408 308848
rect 288992 308388 289044 308440
rect 310704 307844 310756 307896
rect 250168 307819 250220 307828
rect 250168 307785 250177 307819
rect 250177 307785 250211 307819
rect 250211 307785 250220 307819
rect 250168 307776 250220 307785
rect 251548 307819 251600 307828
rect 251548 307785 251557 307819
rect 251557 307785 251591 307819
rect 251591 307785 251600 307819
rect 251548 307776 251600 307785
rect 259736 307776 259788 307828
rect 259920 307776 259972 307828
rect 301136 307776 301188 307828
rect 306748 307776 306800 307828
rect 325884 307819 325936 307828
rect 325884 307785 325893 307819
rect 325893 307785 325927 307819
rect 325927 307785 325936 307819
rect 325884 307776 325936 307785
rect 421196 307819 421248 307828
rect 421196 307785 421205 307819
rect 421205 307785 421239 307819
rect 421239 307785 421248 307819
rect 421196 307776 421248 307785
rect 232320 307751 232372 307760
rect 232320 307717 232329 307751
rect 232329 307717 232363 307751
rect 232363 307717 232372 307751
rect 232320 307708 232372 307717
rect 301228 307640 301280 307692
rect 310704 307751 310756 307760
rect 310704 307717 310713 307751
rect 310713 307717 310747 307751
rect 310747 307717 310756 307751
rect 310704 307708 310756 307717
rect 337200 307708 337252 307760
rect 306932 307640 306984 307692
rect 285772 306416 285824 306468
rect 267832 306348 267884 306400
rect 268016 306348 268068 306400
rect 273076 306348 273128 306400
rect 273260 306348 273312 306400
rect 284576 306391 284628 306400
rect 284576 306357 284585 306391
rect 284585 306357 284619 306391
rect 284619 306357 284628 306391
rect 284576 306348 284628 306357
rect 317512 306348 317564 306400
rect 317696 306348 317748 306400
rect 330208 306348 330260 306400
rect 330392 306348 330444 306400
rect 358544 306348 358596 306400
rect 358728 306348 358780 306400
rect 463700 306348 463752 306400
rect 463884 306348 463936 306400
rect 290188 306280 290240 306332
rect 294328 304920 294380 304972
rect 294236 304852 294288 304904
rect 245936 302447 245988 302456
rect 245936 302413 245945 302447
rect 245945 302413 245979 302447
rect 245979 302413 245988 302447
rect 245936 302404 245988 302413
rect 270684 302268 270736 302320
rect 272156 302268 272208 302320
rect 270776 302064 270828 302116
rect 330208 302268 330260 302320
rect 424140 302200 424192 302252
rect 424508 302200 424560 302252
rect 330116 302132 330168 302184
rect 272248 302064 272300 302116
rect 339868 299931 339920 299940
rect 339868 299897 339877 299931
rect 339877 299897 339911 299931
rect 339911 299897 339920 299931
rect 339868 299888 339920 299897
rect 239220 299480 239272 299532
rect 299848 299480 299900 299532
rect 302516 299480 302568 299532
rect 302608 299480 302660 299532
rect 306840 299523 306892 299532
rect 306840 299489 306849 299523
rect 306849 299489 306883 299523
rect 306883 299489 306892 299523
rect 306840 299480 306892 299489
rect 341156 299523 341208 299532
rect 341156 299489 341165 299523
rect 341165 299489 341199 299523
rect 341199 299489 341208 299523
rect 341156 299480 341208 299489
rect 367008 299523 367060 299532
rect 367008 299489 367017 299523
rect 367017 299489 367051 299523
rect 367051 299489 367060 299523
rect 367008 299480 367060 299489
rect 389272 299523 389324 299532
rect 389272 299489 389281 299523
rect 389281 299489 389315 299523
rect 389315 299489 389324 299523
rect 389272 299480 389324 299489
rect 470600 299523 470652 299532
rect 470600 299489 470609 299523
rect 470609 299489 470643 299523
rect 470643 299489 470652 299523
rect 470600 299480 470652 299489
rect 323308 299455 323360 299464
rect 323308 299421 323317 299455
rect 323317 299421 323351 299455
rect 323351 299421 323360 299455
rect 323308 299412 323360 299421
rect 324688 299455 324740 299464
rect 324688 299421 324697 299455
rect 324697 299421 324731 299455
rect 324731 299421 324740 299455
rect 324688 299412 324740 299421
rect 325884 299412 325936 299464
rect 372712 299455 372764 299464
rect 372712 299421 372721 299455
rect 372721 299421 372755 299455
rect 372755 299421 372764 299455
rect 372712 299412 372764 299421
rect 469956 299412 470008 299464
rect 579804 299412 579856 299464
rect 325976 299344 326028 299396
rect 232320 298163 232372 298172
rect 232320 298129 232329 298163
rect 232329 298129 232363 298163
rect 232363 298129 232372 298163
rect 232320 298120 232372 298129
rect 262496 298120 262548 298172
rect 262680 298120 262732 298172
rect 236276 298095 236328 298104
rect 236276 298061 236285 298095
rect 236285 298061 236319 298095
rect 236319 298061 236328 298095
rect 236276 298052 236328 298061
rect 250168 298095 250220 298104
rect 250168 298061 250177 298095
rect 250177 298061 250211 298095
rect 250211 298061 250220 298095
rect 250168 298052 250220 298061
rect 251548 298052 251600 298104
rect 295616 298188 295668 298240
rect 337016 298231 337068 298240
rect 337016 298197 337025 298231
rect 337025 298197 337059 298231
rect 337059 298197 337068 298231
rect 337016 298188 337068 298197
rect 358728 298188 358780 298240
rect 310888 298120 310940 298172
rect 358636 298120 358688 298172
rect 325976 298095 326028 298104
rect 325976 298061 325985 298095
rect 325985 298061 326019 298095
rect 326019 298061 326028 298095
rect 325976 298052 326028 298061
rect 327264 298052 327316 298104
rect 337016 298052 337068 298104
rect 359096 298052 359148 298104
rect 359188 298052 359240 298104
rect 421196 298095 421248 298104
rect 421196 298061 421205 298095
rect 421205 298061 421239 298095
rect 421239 298061 421248 298095
rect 421196 298052 421248 298061
rect 232320 297984 232372 298036
rect 246028 297984 246080 298036
rect 295524 297984 295576 298036
rect 273260 296692 273312 296744
rect 273536 296692 273588 296744
rect 285772 296692 285824 296744
rect 286048 296692 286100 296744
rect 296812 296692 296864 296744
rect 296904 296692 296956 296744
rect 301044 296692 301096 296744
rect 301412 296692 301464 296744
rect 306840 296735 306892 296744
rect 306840 296701 306849 296735
rect 306849 296701 306883 296735
rect 306883 296701 306892 296735
rect 306840 296692 306892 296701
rect 362224 296692 362276 296744
rect 362408 296692 362460 296744
rect 273628 296667 273680 296676
rect 273628 296633 273637 296667
rect 273637 296633 273671 296667
rect 273671 296633 273680 296667
rect 273628 296624 273680 296633
rect 299848 296624 299900 296676
rect 299940 296624 299992 296676
rect 302608 296624 302660 296676
rect 302700 296624 302752 296676
rect 310888 293063 310940 293072
rect 310888 293029 310897 293063
rect 310897 293029 310931 293063
rect 310931 293029 310940 293063
rect 310888 293020 310940 293029
rect 239036 292544 239088 292596
rect 239220 292544 239272 292596
rect 306840 292612 306892 292664
rect 306748 292476 306800 292528
rect 337200 292451 337252 292460
rect 337200 292417 337209 292451
rect 337209 292417 337243 292451
rect 337243 292417 337252 292451
rect 337200 292408 337252 292417
rect 285772 291864 285824 291916
rect 286048 291864 286100 291916
rect 288716 290003 288768 290012
rect 288716 289969 288725 290003
rect 288725 289969 288759 290003
rect 288759 289969 288768 290003
rect 288716 289960 288768 289969
rect 262496 289824 262548 289876
rect 262680 289824 262732 289876
rect 267832 289824 267884 289876
rect 267924 289824 267976 289876
rect 324688 289867 324740 289876
rect 324688 289833 324697 289867
rect 324697 289833 324731 289867
rect 324731 289833 324740 289867
rect 324688 289824 324740 289833
rect 372712 289867 372764 289876
rect 372712 289833 372721 289867
rect 372721 289833 372755 289867
rect 372755 289833 372764 289867
rect 372712 289824 372764 289833
rect 375840 289824 375892 289876
rect 375932 289824 375984 289876
rect 377128 289824 377180 289876
rect 377220 289824 377272 289876
rect 250168 289799 250220 289808
rect 250168 289765 250177 289799
rect 250177 289765 250211 289799
rect 250211 289765 250220 289799
rect 250168 289756 250220 289765
rect 270684 289756 270736 289808
rect 270776 289756 270828 289808
rect 272248 289756 272300 289808
rect 284576 289756 284628 289808
rect 288716 289756 288768 289808
rect 288808 289756 288860 289808
rect 341248 289756 341300 289808
rect 367008 289799 367060 289808
rect 367008 289765 367017 289799
rect 367017 289765 367051 289799
rect 367051 289765 367060 289799
rect 367008 289756 367060 289765
rect 389456 289756 389508 289808
rect 470600 289799 470652 289808
rect 470600 289765 470609 289799
rect 470609 289765 470643 289799
rect 470643 289765 470652 289799
rect 470600 289756 470652 289765
rect 284760 289688 284812 289740
rect 232228 288439 232280 288448
rect 232228 288405 232237 288439
rect 232237 288405 232271 288439
rect 232271 288405 232280 288439
rect 232228 288396 232280 288405
rect 236276 288439 236328 288448
rect 236276 288405 236285 288439
rect 236285 288405 236319 288439
rect 236319 288405 236328 288439
rect 236276 288396 236328 288405
rect 251364 288439 251416 288448
rect 251364 288405 251373 288439
rect 251373 288405 251407 288439
rect 251407 288405 251416 288439
rect 251364 288396 251416 288405
rect 323492 288396 323544 288448
rect 325976 288439 326028 288448
rect 325976 288405 325985 288439
rect 325985 288405 326019 288439
rect 326019 288405 326028 288439
rect 325976 288396 326028 288405
rect 327172 288439 327224 288448
rect 327172 288405 327181 288439
rect 327181 288405 327215 288439
rect 327215 288405 327224 288439
rect 327172 288396 327224 288405
rect 330300 288439 330352 288448
rect 330300 288405 330309 288439
rect 330309 288405 330343 288439
rect 330343 288405 330352 288439
rect 330300 288396 330352 288405
rect 357440 288396 357492 288448
rect 357624 288396 357676 288448
rect 358636 288396 358688 288448
rect 358728 288396 358780 288448
rect 421196 288439 421248 288448
rect 421196 288405 421205 288439
rect 421205 288405 421239 288439
rect 421239 288405 421248 288439
rect 421196 288396 421248 288405
rect 273628 287079 273680 287088
rect 273628 287045 273637 287079
rect 273637 287045 273671 287079
rect 273671 287045 273680 287079
rect 273628 287036 273680 287045
rect 330300 287079 330352 287088
rect 330300 287045 330309 287079
rect 330309 287045 330343 287079
rect 330343 287045 330352 287079
rect 330300 287036 330352 287045
rect 463700 287036 463752 287088
rect 463884 287036 463936 287088
rect 259552 285608 259604 285660
rect 259920 285608 259972 285660
rect 272340 283568 272392 283620
rect 236276 282888 236328 282940
rect 239128 282888 239180 282940
rect 337108 282931 337160 282940
rect 337108 282897 337117 282931
rect 337117 282897 337151 282931
rect 337151 282897 337160 282931
rect 337108 282888 337160 282897
rect 339684 282888 339736 282940
rect 339868 282888 339920 282940
rect 424508 282888 424560 282940
rect 424692 282888 424744 282940
rect 236460 282752 236512 282804
rect 239220 282752 239272 282804
rect 310888 282795 310940 282804
rect 310888 282761 310897 282795
rect 310897 282761 310931 282795
rect 310931 282761 310940 282795
rect 310888 282752 310940 282761
rect 232228 280168 232280 280220
rect 232320 280168 232372 280220
rect 341156 280211 341208 280220
rect 341156 280177 341165 280211
rect 341165 280177 341199 280211
rect 341199 280177 341208 280211
rect 341156 280168 341208 280177
rect 367008 280211 367060 280220
rect 367008 280177 367017 280211
rect 367017 280177 367051 280211
rect 367051 280177 367060 280211
rect 367008 280168 367060 280177
rect 389364 280211 389416 280220
rect 389364 280177 389373 280211
rect 389373 280177 389407 280211
rect 389407 280177 389416 280211
rect 389364 280168 389416 280177
rect 470600 280211 470652 280220
rect 470600 280177 470609 280211
rect 470609 280177 470643 280211
rect 470643 280177 470652 280211
rect 470600 280168 470652 280177
rect 250076 280100 250128 280152
rect 250168 280100 250220 280152
rect 270684 280143 270736 280152
rect 270684 280109 270693 280143
rect 270693 280109 270727 280143
rect 270727 280109 270736 280143
rect 270684 280100 270736 280109
rect 273536 280143 273588 280152
rect 273536 280109 273545 280143
rect 273545 280109 273579 280143
rect 273579 280109 273588 280143
rect 273536 280100 273588 280109
rect 284576 280100 284628 280152
rect 284760 280100 284812 280152
rect 288808 280100 288860 280152
rect 288900 280100 288952 280152
rect 323308 280100 323360 280152
rect 323400 280100 323452 280152
rect 372712 280143 372764 280152
rect 372712 280109 372721 280143
rect 372721 280109 372755 280143
rect 372755 280109 372764 280143
rect 372712 280100 372764 280109
rect 375840 280143 375892 280152
rect 375840 280109 375849 280143
rect 375849 280109 375883 280143
rect 375883 280109 375892 280143
rect 375840 280100 375892 280109
rect 377128 280143 377180 280152
rect 377128 280109 377137 280143
rect 377137 280109 377171 280143
rect 377171 280109 377180 280143
rect 377128 280100 377180 280109
rect 424600 280143 424652 280152
rect 424600 280109 424609 280143
rect 424609 280109 424643 280143
rect 424643 280109 424652 280143
rect 424600 280100 424652 280109
rect 265164 278740 265216 278792
rect 265256 278740 265308 278792
rect 267740 278740 267792 278792
rect 267832 278740 267884 278792
rect 285772 278740 285824 278792
rect 286048 278740 286100 278792
rect 295248 278740 295300 278792
rect 295524 278740 295576 278792
rect 301044 278740 301096 278792
rect 301228 278740 301280 278792
rect 327356 278740 327408 278792
rect 327540 278740 327592 278792
rect 337108 278783 337160 278792
rect 337108 278749 337117 278783
rect 337117 278749 337151 278783
rect 337151 278749 337160 278783
rect 337108 278740 337160 278749
rect 310888 278715 310940 278724
rect 310888 278681 310897 278715
rect 310897 278681 310931 278715
rect 310931 278681 310940 278715
rect 310888 278672 310940 278681
rect 324504 278715 324556 278724
rect 324504 278681 324513 278715
rect 324513 278681 324547 278715
rect 324547 278681 324556 278715
rect 324504 278672 324556 278681
rect 295524 277856 295576 277908
rect 295800 277856 295852 277908
rect 307024 277448 307076 277500
rect 290004 277380 290056 277432
rect 290096 277380 290148 277432
rect 296812 277380 296864 277432
rect 297088 277380 297140 277432
rect 306840 277380 306892 277432
rect 330116 277380 330168 277432
rect 330300 277380 330352 277432
rect 357716 277380 357768 277432
rect 357808 277380 357860 277432
rect 362224 277355 362276 277364
rect 362224 277321 362233 277355
rect 362233 277321 362267 277355
rect 362267 277321 362276 277355
rect 362224 277312 362276 277321
rect 330116 277287 330168 277296
rect 330116 277253 330125 277287
rect 330125 277253 330159 277287
rect 330159 277253 330168 277287
rect 330116 277244 330168 277253
rect 270684 275315 270736 275324
rect 270684 275281 270693 275315
rect 270693 275281 270727 275315
rect 270727 275281 270736 275315
rect 270684 275272 270736 275281
rect 236276 273232 236328 273284
rect 236460 273232 236512 273284
rect 239036 273232 239088 273284
rect 239220 273232 239272 273284
rect 301044 273232 301096 273284
rect 337108 273232 337160 273284
rect 301136 273164 301188 273216
rect 359004 273164 359056 273216
rect 359188 273164 359240 273216
rect 337200 273096 337252 273148
rect 357440 272552 357492 272604
rect 357900 272552 357952 272604
rect 294236 270580 294288 270632
rect 232228 270555 232280 270564
rect 232228 270521 232237 270555
rect 232237 270521 232271 270555
rect 232271 270521 232280 270555
rect 232228 270512 232280 270521
rect 251180 270512 251232 270564
rect 251456 270512 251508 270564
rect 273628 270512 273680 270564
rect 294144 270444 294196 270496
rect 372712 270555 372764 270564
rect 372712 270521 372721 270555
rect 372721 270521 372755 270555
rect 372755 270521 372764 270555
rect 372712 270512 372764 270521
rect 375840 270555 375892 270564
rect 375840 270521 375849 270555
rect 375849 270521 375883 270555
rect 375883 270521 375892 270555
rect 375840 270512 375892 270521
rect 377128 270555 377180 270564
rect 377128 270521 377137 270555
rect 377137 270521 377171 270555
rect 377171 270521 377180 270555
rect 377128 270512 377180 270521
rect 424784 270512 424836 270564
rect 301136 270444 301188 270496
rect 301228 270444 301280 270496
rect 327264 270444 327316 270496
rect 327356 270444 327408 270496
rect 341248 270444 341300 270496
rect 367008 270487 367060 270496
rect 367008 270453 367017 270487
rect 367017 270453 367051 270487
rect 367051 270453 367060 270487
rect 367008 270444 367060 270453
rect 389456 270444 389508 270496
rect 470600 270487 470652 270496
rect 470600 270453 470609 270487
rect 470609 270453 470643 270487
rect 470643 270453 470652 270487
rect 470600 270444 470652 270453
rect 232228 269127 232280 269136
rect 232228 269093 232237 269127
rect 232237 269093 232271 269127
rect 232271 269093 232280 269127
rect 232228 269084 232280 269093
rect 250076 269084 250128 269136
rect 250260 269084 250312 269136
rect 262588 269084 262640 269136
rect 262680 269084 262732 269136
rect 284576 269084 284628 269136
rect 284760 269084 284812 269136
rect 288808 269084 288860 269136
rect 288900 269084 288952 269136
rect 324596 269084 324648 269136
rect 421196 269084 421248 269136
rect 421380 269084 421432 269136
rect 267832 267724 267884 267776
rect 268016 267724 268068 267776
rect 299664 267724 299716 267776
rect 299848 267724 299900 267776
rect 463700 267724 463752 267776
rect 463884 267724 463936 267776
rect 236276 263576 236328 263628
rect 239128 263576 239180 263628
rect 270684 263576 270736 263628
rect 236460 263440 236512 263492
rect 325976 263644 326028 263696
rect 337108 263619 337160 263628
rect 337108 263585 337117 263619
rect 337117 263585 337151 263619
rect 337151 263585 337160 263619
rect 337108 263576 337160 263585
rect 339684 263576 339736 263628
rect 339868 263576 339920 263628
rect 360292 263576 360344 263628
rect 360476 263576 360528 263628
rect 325884 263508 325936 263560
rect 239220 263440 239272 263492
rect 270684 263440 270736 263492
rect 310888 263483 310940 263492
rect 310888 263449 310897 263483
rect 310897 263449 310931 263483
rect 310931 263449 310940 263483
rect 310888 263440 310940 263449
rect 362224 263483 362276 263492
rect 362224 263449 362233 263483
rect 362233 263449 362267 263483
rect 362267 263449 362276 263483
rect 362224 263440 362276 263449
rect 330116 263211 330168 263220
rect 330116 263177 330125 263211
rect 330125 263177 330159 263211
rect 330159 263177 330168 263211
rect 330116 263168 330168 263177
rect 264980 262896 265032 262948
rect 265164 262896 265216 262948
rect 306840 262939 306892 262948
rect 306840 262905 306849 262939
rect 306849 262905 306883 262939
rect 306883 262905 306892 262939
rect 306840 262896 306892 262905
rect 232228 260856 232280 260908
rect 232320 260856 232372 260908
rect 250076 260856 250128 260908
rect 250168 260856 250220 260908
rect 266728 260856 266780 260908
rect 270684 260831 270736 260840
rect 270684 260797 270693 260831
rect 270693 260797 270727 260831
rect 270727 260797 270736 260831
rect 270684 260788 270736 260797
rect 272340 260924 272392 260976
rect 284576 260856 284628 260908
rect 284760 260856 284812 260908
rect 341156 260899 341208 260908
rect 341156 260865 341165 260899
rect 341165 260865 341199 260899
rect 341199 260865 341208 260899
rect 341156 260856 341208 260865
rect 359096 260856 359148 260908
rect 359188 260856 359240 260908
rect 367008 260899 367060 260908
rect 367008 260865 367017 260899
rect 367017 260865 367051 260899
rect 367051 260865 367060 260899
rect 367008 260856 367060 260865
rect 389364 260899 389416 260908
rect 389364 260865 389373 260899
rect 389373 260865 389407 260899
rect 389407 260865 389416 260899
rect 389364 260856 389416 260865
rect 470600 260899 470652 260908
rect 470600 260865 470609 260899
rect 470609 260865 470643 260899
rect 470643 260865 470652 260899
rect 470600 260856 470652 260865
rect 273536 260831 273588 260840
rect 273536 260797 273545 260831
rect 273545 260797 273579 260831
rect 273579 260797 273588 260831
rect 273536 260788 273588 260797
rect 324596 260788 324648 260840
rect 372712 260831 372764 260840
rect 372712 260797 372721 260831
rect 372721 260797 372755 260831
rect 372755 260797 372764 260831
rect 372712 260788 372764 260797
rect 375840 260831 375892 260840
rect 375840 260797 375849 260831
rect 375849 260797 375883 260831
rect 375883 260797 375892 260831
rect 375840 260788 375892 260797
rect 377128 260831 377180 260840
rect 377128 260797 377137 260831
rect 377137 260797 377171 260831
rect 377171 260797 377180 260831
rect 377128 260788 377180 260797
rect 424600 260788 424652 260840
rect 463792 260788 463844 260840
rect 266728 260720 266780 260772
rect 272156 260720 272208 260772
rect 324688 260720 324740 260772
rect 267740 259428 267792 259480
rect 267832 259428 267884 259480
rect 296996 259428 297048 259480
rect 297088 259428 297140 259480
rect 337108 259471 337160 259480
rect 337108 259437 337117 259471
rect 337117 259437 337151 259471
rect 337151 259437 337160 259471
rect 337108 259428 337160 259437
rect 299848 259360 299900 259412
rect 300032 259360 300084 259412
rect 330116 259360 330168 259412
rect 330208 259360 330260 259412
rect 251180 259020 251232 259072
rect 251364 259020 251416 259072
rect 288808 258000 288860 258052
rect 288992 258000 289044 258052
rect 290096 258000 290148 258052
rect 294236 258043 294288 258052
rect 294236 258009 294245 258043
rect 294245 258009 294279 258043
rect 294279 258009 294288 258043
rect 294236 258000 294288 258009
rect 296996 258000 297048 258052
rect 297180 258000 297232 258052
rect 330208 258000 330260 258052
rect 330392 258000 330444 258052
rect 245844 257932 245896 257984
rect 245936 257932 245988 257984
rect 310888 256071 310940 256080
rect 310888 256037 310897 256071
rect 310897 256037 310931 256071
rect 310931 256037 310940 256071
rect 310888 256028 310940 256037
rect 270684 256003 270736 256012
rect 270684 255969 270693 256003
rect 270693 255969 270727 256003
rect 270727 255969 270736 256003
rect 270684 255960 270736 255969
rect 336740 254600 336792 254652
rect 337108 254600 337160 254652
rect 236276 253920 236328 253972
rect 236460 253920 236512 253972
rect 239036 253920 239088 253972
rect 239220 253920 239272 253972
rect 250076 253963 250128 253972
rect 250076 253929 250085 253963
rect 250085 253929 250119 253963
rect 250119 253929 250128 253963
rect 250076 253920 250128 253929
rect 362316 253920 362368 253972
rect 357532 253852 357584 253904
rect 357716 253852 357768 253904
rect 359004 253852 359056 253904
rect 359188 253852 359240 253904
rect 362224 253852 362276 253904
rect 323400 252739 323452 252748
rect 323400 252705 323409 252739
rect 323409 252705 323443 252739
rect 323443 252705 323452 252739
rect 323400 252696 323452 252705
rect 2780 252492 2832 252544
rect 5264 252492 5316 252544
rect 469864 252492 469916 252544
rect 580172 252492 580224 252544
rect 232320 251268 232372 251320
rect 310704 251268 310756 251320
rect 265164 251200 265216 251252
rect 265256 251200 265308 251252
rect 267740 251200 267792 251252
rect 267832 251200 267884 251252
rect 273628 251200 273680 251252
rect 291476 251200 291528 251252
rect 291568 251200 291620 251252
rect 372712 251243 372764 251252
rect 372712 251209 372721 251243
rect 372721 251209 372755 251243
rect 372755 251209 372764 251243
rect 372712 251200 372764 251209
rect 375840 251243 375892 251252
rect 375840 251209 375849 251243
rect 375849 251209 375883 251243
rect 375883 251209 375892 251243
rect 375840 251200 375892 251209
rect 377128 251243 377180 251252
rect 377128 251209 377137 251243
rect 377137 251209 377171 251243
rect 377171 251209 377180 251243
rect 377128 251200 377180 251209
rect 389180 251200 389232 251252
rect 389364 251200 389416 251252
rect 424508 251243 424560 251252
rect 424508 251209 424517 251243
rect 424517 251209 424551 251243
rect 424551 251209 424560 251243
rect 424508 251200 424560 251209
rect 463700 251243 463752 251252
rect 463700 251209 463709 251243
rect 463709 251209 463743 251243
rect 463743 251209 463752 251243
rect 463700 251200 463752 251209
rect 239128 251132 239180 251184
rect 239220 251132 239272 251184
rect 259736 251132 259788 251184
rect 262680 251132 262732 251184
rect 262772 251132 262824 251184
rect 266728 251132 266780 251184
rect 295524 251132 295576 251184
rect 295708 251132 295760 251184
rect 310704 251175 310756 251184
rect 310704 251141 310713 251175
rect 310713 251141 310747 251175
rect 310747 251141 310756 251175
rect 310704 251132 310756 251141
rect 325884 251175 325936 251184
rect 325884 251141 325893 251175
rect 325893 251141 325927 251175
rect 325927 251141 325936 251175
rect 325884 251132 325936 251141
rect 357624 251132 357676 251184
rect 357716 251132 357768 251184
rect 367008 251175 367060 251184
rect 367008 251141 367017 251175
rect 367017 251141 367051 251175
rect 367051 251141 367060 251175
rect 367008 251132 367060 251141
rect 470600 251175 470652 251184
rect 470600 251141 470609 251175
rect 470609 251141 470643 251175
rect 470643 251141 470652 251175
rect 470600 251132 470652 251141
rect 232228 251064 232280 251116
rect 266728 250996 266780 251048
rect 327356 249908 327408 249960
rect 284668 249840 284720 249892
rect 284760 249840 284812 249892
rect 324596 249840 324648 249892
rect 324688 249840 324740 249892
rect 327172 249840 327224 249892
rect 250076 249815 250128 249824
rect 250076 249781 250085 249815
rect 250085 249781 250119 249815
rect 250119 249781 250128 249815
rect 250076 249772 250128 249781
rect 285956 249772 286008 249824
rect 286048 249772 286100 249824
rect 306932 249772 306984 249824
rect 325884 249815 325936 249824
rect 325884 249781 325893 249815
rect 325893 249781 325927 249815
rect 325927 249781 325936 249815
rect 325884 249772 325936 249781
rect 358544 249772 358596 249824
rect 358728 249772 358780 249824
rect 421196 249772 421248 249824
rect 421380 249772 421432 249824
rect 284668 249747 284720 249756
rect 284668 249713 284677 249747
rect 284677 249713 284711 249747
rect 284711 249713 284720 249747
rect 284668 249704 284720 249713
rect 327172 249747 327224 249756
rect 327172 249713 327181 249747
rect 327181 249713 327215 249747
rect 327215 249713 327224 249747
rect 327172 249704 327224 249713
rect 290004 248455 290056 248464
rect 290004 248421 290013 248455
rect 290013 248421 290047 248455
rect 290047 248421 290056 248455
rect 290004 248412 290056 248421
rect 294236 248455 294288 248464
rect 294236 248421 294245 248455
rect 294245 248421 294279 248455
rect 294279 248421 294288 248455
rect 294236 248412 294288 248421
rect 291476 248387 291528 248396
rect 291476 248353 291485 248387
rect 291485 248353 291519 248387
rect 291519 248353 291528 248387
rect 291476 248344 291528 248353
rect 290004 245828 290056 245880
rect 290372 245828 290424 245880
rect 285956 244987 286008 244996
rect 285956 244953 285965 244987
rect 285965 244953 285999 244987
rect 285999 244953 286008 244987
rect 285956 244944 286008 244953
rect 272156 244332 272208 244384
rect 236276 244264 236328 244316
rect 270684 244307 270736 244316
rect 270684 244273 270693 244307
rect 270693 244273 270727 244307
rect 270727 244273 270736 244307
rect 270684 244264 270736 244273
rect 339684 244264 339736 244316
rect 339868 244264 339920 244316
rect 341248 244332 341300 244384
rect 360292 244264 360344 244316
rect 360476 244264 360528 244316
rect 272156 244196 272208 244248
rect 341156 244196 341208 244248
rect 236460 244128 236512 244180
rect 259644 242675 259696 242684
rect 259644 242641 259653 242675
rect 259653 242641 259687 242675
rect 259687 242641 259696 242675
rect 259644 242632 259696 242641
rect 358728 241612 358780 241664
rect 270684 241587 270736 241596
rect 270684 241553 270693 241587
rect 270693 241553 270727 241587
rect 270727 241553 270736 241587
rect 270684 241544 270736 241553
rect 388996 241544 389048 241596
rect 389272 241544 389324 241596
rect 250076 241476 250128 241528
rect 250168 241476 250220 241528
rect 251364 241519 251416 241528
rect 251364 241485 251373 241519
rect 251373 241485 251407 241519
rect 251407 241485 251416 241519
rect 251364 241476 251416 241485
rect 310888 241476 310940 241528
rect 323400 241519 323452 241528
rect 323400 241485 323409 241519
rect 323409 241485 323443 241519
rect 323443 241485 323452 241519
rect 323400 241476 323452 241485
rect 358728 241476 358780 241528
rect 359096 241476 359148 241528
rect 359188 241476 359240 241528
rect 367008 241519 367060 241528
rect 367008 241485 367017 241519
rect 367017 241485 367051 241519
rect 367051 241485 367060 241519
rect 367008 241476 367060 241485
rect 470600 241519 470652 241528
rect 470600 241485 470609 241519
rect 470609 241485 470643 241519
rect 470643 241485 470652 241519
rect 470600 241476 470652 241485
rect 270684 241451 270736 241460
rect 270684 241417 270693 241451
rect 270693 241417 270727 241451
rect 270727 241417 270736 241451
rect 270684 241408 270736 241417
rect 299480 241451 299532 241460
rect 299480 241417 299489 241451
rect 299489 241417 299523 241451
rect 299523 241417 299532 241451
rect 362224 241451 362276 241460
rect 299480 241408 299532 241417
rect 362224 241417 362233 241451
rect 362233 241417 362267 241451
rect 362267 241417 362276 241451
rect 362224 241408 362276 241417
rect 375840 241451 375892 241460
rect 375840 241417 375849 241451
rect 375849 241417 375883 241451
rect 375883 241417 375892 241451
rect 375840 241408 375892 241417
rect 389272 241451 389324 241460
rect 389272 241417 389281 241451
rect 389281 241417 389315 241451
rect 389315 241417 389324 241451
rect 389272 241408 389324 241417
rect 327172 240227 327224 240236
rect 327172 240193 327181 240227
rect 327181 240193 327215 240227
rect 327215 240193 327224 240227
rect 327172 240184 327224 240193
rect 232320 240116 232372 240168
rect 232504 240116 232556 240168
rect 244372 240116 244424 240168
rect 244464 240116 244516 240168
rect 245844 240116 245896 240168
rect 245936 240116 245988 240168
rect 251364 240159 251416 240168
rect 251364 240125 251373 240159
rect 251373 240125 251407 240159
rect 251407 240125 251416 240159
rect 251364 240116 251416 240125
rect 284852 240116 284904 240168
rect 299940 240116 299992 240168
rect 300032 240116 300084 240168
rect 302424 240116 302476 240168
rect 302700 240116 302752 240168
rect 306932 240116 306984 240168
rect 307116 240116 307168 240168
rect 324596 240116 324648 240168
rect 324688 240116 324740 240168
rect 325976 240116 326028 240168
rect 326160 240116 326212 240168
rect 337108 240116 337160 240168
rect 337292 240116 337344 240168
rect 291752 240048 291804 240100
rect 327172 240091 327224 240100
rect 327172 240057 327181 240091
rect 327181 240057 327215 240091
rect 327215 240057 327224 240091
rect 327172 240048 327224 240057
rect 330116 240048 330168 240100
rect 330208 240048 330260 240100
rect 330208 238688 330260 238740
rect 330392 238620 330444 238672
rect 3056 237328 3108 237380
rect 15844 237328 15896 237380
rect 244372 234855 244424 234864
rect 244372 234821 244381 234855
rect 244381 234821 244415 234855
rect 244415 234821 244424 234855
rect 244372 234812 244424 234821
rect 250076 234608 250128 234660
rect 310888 234676 310940 234728
rect 323400 234719 323452 234728
rect 323400 234685 323409 234719
rect 323409 234685 323443 234719
rect 323443 234685 323452 234719
rect 323400 234676 323452 234685
rect 389456 234608 389508 234660
rect 310796 234540 310848 234592
rect 285956 234515 286008 234524
rect 285956 234481 285965 234515
rect 285965 234481 285999 234515
rect 285999 234481 286008 234515
rect 285956 234472 286008 234481
rect 270684 232067 270736 232076
rect 270684 232033 270693 232067
rect 270693 232033 270727 232067
rect 270727 232033 270736 232067
rect 270684 232024 270736 232033
rect 302700 231956 302752 232008
rect 236276 231888 236328 231940
rect 236552 231888 236604 231940
rect 266728 231931 266780 231940
rect 266728 231897 266737 231931
rect 266737 231897 266771 231931
rect 266771 231897 266780 231931
rect 266728 231888 266780 231897
rect 262680 231820 262732 231872
rect 262772 231820 262824 231872
rect 265256 231820 265308 231872
rect 265348 231820 265400 231872
rect 299480 231863 299532 231872
rect 299480 231829 299489 231863
rect 299489 231829 299523 231863
rect 299523 231829 299532 231863
rect 299480 231820 299532 231829
rect 301136 231888 301188 231940
rect 366824 231888 366876 231940
rect 367008 231888 367060 231940
rect 306932 231820 306984 231872
rect 357624 231820 357676 231872
rect 357716 231820 357768 231872
rect 359096 231820 359148 231872
rect 359188 231820 359240 231872
rect 372528 231820 372580 231872
rect 372712 231820 372764 231872
rect 375840 231863 375892 231872
rect 375840 231829 375849 231863
rect 375849 231829 375883 231863
rect 375883 231829 375892 231863
rect 375840 231820 375892 231829
rect 376944 231820 376996 231872
rect 377128 231820 377180 231872
rect 301044 231752 301096 231804
rect 306748 231752 306800 231804
rect 310796 231795 310848 231804
rect 310796 231761 310805 231795
rect 310805 231761 310839 231795
rect 310839 231761 310848 231795
rect 310796 231752 310848 231761
rect 323400 231795 323452 231804
rect 323400 231761 323409 231795
rect 323409 231761 323443 231795
rect 323443 231761 323452 231795
rect 323400 231752 323452 231761
rect 324596 231752 324648 231804
rect 324780 231752 324832 231804
rect 367008 231795 367060 231804
rect 367008 231761 367017 231795
rect 367017 231761 367051 231795
rect 367051 231761 367060 231795
rect 367008 231752 367060 231761
rect 327172 230571 327224 230580
rect 327172 230537 327181 230571
rect 327181 230537 327215 230571
rect 327215 230537 327224 230571
rect 327172 230528 327224 230537
rect 337016 230528 337068 230580
rect 337200 230528 337252 230580
rect 244372 230503 244424 230512
rect 244372 230469 244381 230503
rect 244381 230469 244415 230503
rect 244415 230469 244424 230503
rect 244372 230460 244424 230469
rect 245936 230460 245988 230512
rect 246120 230460 246172 230512
rect 250168 230503 250220 230512
rect 250168 230469 250177 230503
rect 250177 230469 250211 230503
rect 250211 230469 250220 230503
rect 250168 230460 250220 230469
rect 251088 230460 251140 230512
rect 251364 230460 251416 230512
rect 259552 230460 259604 230512
rect 259828 230460 259880 230512
rect 266728 230503 266780 230512
rect 266728 230469 266737 230503
rect 266737 230469 266771 230503
rect 266771 230469 266780 230503
rect 266728 230460 266780 230469
rect 267924 230460 267976 230512
rect 268108 230460 268160 230512
rect 302608 230503 302660 230512
rect 302608 230469 302617 230503
rect 302617 230469 302651 230503
rect 302651 230469 302660 230503
rect 302608 230460 302660 230469
rect 341248 230460 341300 230512
rect 341432 230460 341484 230512
rect 358544 230460 358596 230512
rect 358728 230460 358780 230512
rect 362408 230460 362460 230512
rect 421196 230460 421248 230512
rect 421380 230460 421432 230512
rect 244280 229032 244332 229084
rect 244372 229032 244424 229084
rect 284852 225020 284904 225072
rect 236276 224952 236328 225004
rect 270684 224995 270736 225004
rect 270684 224961 270693 224995
rect 270693 224961 270727 224995
rect 270727 224961 270736 224995
rect 270684 224952 270736 224961
rect 339684 224952 339736 225004
rect 339868 224952 339920 225004
rect 341248 225020 341300 225072
rect 360292 224952 360344 225004
rect 360476 224952 360528 225004
rect 284852 224884 284904 224936
rect 341156 224884 341208 224936
rect 236460 224816 236512 224868
rect 329932 224204 329984 224256
rect 330208 224204 330260 224256
rect 358728 222300 358780 222352
rect 265256 222232 265308 222284
rect 270684 222275 270736 222284
rect 270684 222241 270693 222275
rect 270693 222241 270727 222275
rect 270727 222241 270736 222275
rect 270684 222232 270736 222241
rect 245844 222164 245896 222216
rect 246028 222164 246080 222216
rect 265164 222164 265216 222216
rect 295524 222164 295576 222216
rect 295616 222164 295668 222216
rect 296812 222164 296864 222216
rect 296904 222164 296956 222216
rect 306748 222164 306800 222216
rect 306932 222164 306984 222216
rect 310888 222164 310940 222216
rect 358728 222164 358780 222216
rect 362224 222164 362276 222216
rect 362408 222164 362460 222216
rect 367008 222207 367060 222216
rect 367008 222173 367017 222207
rect 367017 222173 367051 222207
rect 367051 222173 367060 222207
rect 367008 222164 367060 222173
rect 389272 222164 389324 222216
rect 389548 222164 389600 222216
rect 463792 222164 463844 222216
rect 464068 222164 464120 222216
rect 470416 222164 470468 222216
rect 470600 222164 470652 222216
rect 270684 222139 270736 222148
rect 270684 222105 270693 222139
rect 270693 222105 270727 222139
rect 270727 222105 270736 222139
rect 270684 222096 270736 222105
rect 299480 222139 299532 222148
rect 299480 222105 299489 222139
rect 299489 222105 299523 222139
rect 299523 222105 299532 222139
rect 375840 222139 375892 222148
rect 299480 222096 299532 222105
rect 375840 222105 375849 222139
rect 375849 222105 375883 222139
rect 375883 222105 375892 222139
rect 375840 222096 375892 222105
rect 337108 220872 337160 220924
rect 337384 220872 337436 220924
rect 232320 220804 232372 220856
rect 232504 220804 232556 220856
rect 251548 220804 251600 220856
rect 251640 220804 251692 220856
rect 267740 220804 267792 220856
rect 267924 220804 267976 220856
rect 290188 220804 290240 220856
rect 290372 220804 290424 220856
rect 291660 220804 291712 220856
rect 291844 220804 291896 220856
rect 294328 220804 294380 220856
rect 294420 220804 294472 220856
rect 325884 220804 325936 220856
rect 326068 220804 326120 220856
rect 327356 220804 327408 220856
rect 327540 220804 327592 220856
rect 337108 220736 337160 220788
rect 337292 220736 337344 220788
rect 341156 220779 341208 220788
rect 341156 220745 341165 220779
rect 341165 220745 341199 220779
rect 341199 220745 341208 220779
rect 341156 220736 341208 220745
rect 244464 219376 244516 219428
rect 244556 219376 244608 219428
rect 317512 219376 317564 219428
rect 317696 219376 317748 219428
rect 330116 219419 330168 219428
rect 330116 219385 330125 219419
rect 330125 219385 330159 219419
rect 330159 219385 330168 219419
rect 330116 219376 330168 219385
rect 244464 217991 244516 218000
rect 244464 217957 244473 217991
rect 244473 217957 244507 217991
rect 244507 217957 244516 217991
rect 244464 217948 244516 217957
rect 310888 215364 310940 215416
rect 362316 215296 362368 215348
rect 389548 215364 389600 215416
rect 464068 215364 464120 215416
rect 310796 215228 310848 215280
rect 341156 215271 341208 215280
rect 341156 215237 341165 215271
rect 341165 215237 341199 215271
rect 341199 215237 341208 215271
rect 341156 215228 341208 215237
rect 357532 215228 357584 215280
rect 357716 215228 357768 215280
rect 359004 215228 359056 215280
rect 359188 215228 359240 215280
rect 389456 215228 389508 215280
rect 463976 215228 464028 215280
rect 270684 212755 270736 212764
rect 270684 212721 270693 212755
rect 270693 212721 270727 212755
rect 270727 212721 270736 212755
rect 270684 212712 270736 212721
rect 236276 212576 236328 212628
rect 236460 212576 236512 212628
rect 239128 212576 239180 212628
rect 239404 212576 239456 212628
rect 290188 212576 290240 212628
rect 291660 212576 291712 212628
rect 245844 212508 245896 212560
rect 245936 212508 245988 212560
rect 250076 212508 250128 212560
rect 250260 212508 250312 212560
rect 265164 212508 265216 212560
rect 265256 212508 265308 212560
rect 266636 212508 266688 212560
rect 266820 212508 266872 212560
rect 267740 212508 267792 212560
rect 267832 212508 267884 212560
rect 272156 212551 272208 212560
rect 272156 212517 272165 212551
rect 272165 212517 272199 212551
rect 272199 212517 272208 212551
rect 272156 212508 272208 212517
rect 299480 212551 299532 212560
rect 299480 212517 299489 212551
rect 299489 212517 299523 212551
rect 299523 212517 299532 212551
rect 299480 212508 299532 212517
rect 301136 212576 301188 212628
rect 306932 212576 306984 212628
rect 324688 212508 324740 212560
rect 324780 212508 324832 212560
rect 325884 212508 325936 212560
rect 325976 212508 326028 212560
rect 372528 212508 372580 212560
rect 372712 212508 372764 212560
rect 375840 212551 375892 212560
rect 375840 212517 375849 212551
rect 375849 212517 375883 212551
rect 375883 212517 375892 212551
rect 375840 212508 375892 212517
rect 376944 212508 376996 212560
rect 377128 212508 377180 212560
rect 284668 212440 284720 212492
rect 284852 212440 284904 212492
rect 290188 212440 290240 212492
rect 291660 212440 291712 212492
rect 301044 212440 301096 212492
rect 306748 212440 306800 212492
rect 310796 212483 310848 212492
rect 310796 212449 310805 212483
rect 310805 212449 310839 212483
rect 310839 212449 310848 212483
rect 310796 212440 310848 212449
rect 232320 211216 232372 211268
rect 272156 211191 272208 211200
rect 272156 211157 272165 211191
rect 272165 211157 272199 211191
rect 272199 211157 272208 211191
rect 272156 211148 272208 211157
rect 358544 211148 358596 211200
rect 358636 211148 358688 211200
rect 362132 211191 362184 211200
rect 362132 211157 362141 211191
rect 362141 211157 362175 211191
rect 362175 211157 362184 211191
rect 362132 211148 362184 211157
rect 239036 211080 239088 211132
rect 239312 211080 239364 211132
rect 265256 211123 265308 211132
rect 265256 211089 265265 211123
rect 265265 211089 265299 211123
rect 265299 211089 265308 211123
rect 265256 211080 265308 211089
rect 284668 211080 284720 211132
rect 284944 211080 284996 211132
rect 294236 211080 294288 211132
rect 294328 211080 294380 211132
rect 288808 210944 288860 210996
rect 289176 210944 289228 210996
rect 232228 209831 232280 209840
rect 232228 209797 232237 209831
rect 232237 209797 232271 209831
rect 232271 209797 232280 209831
rect 232228 209788 232280 209797
rect 317512 209788 317564 209840
rect 317696 209788 317748 209840
rect 330116 209831 330168 209840
rect 330116 209797 330125 209831
rect 330125 209797 330159 209831
rect 330159 209797 330168 209831
rect 330116 209788 330168 209797
rect 284668 209720 284720 209772
rect 284760 209720 284812 209772
rect 330208 209763 330260 209772
rect 330208 209729 330217 209763
rect 330217 209729 330251 209763
rect 330251 209729 330260 209763
rect 330208 209720 330260 209729
rect 250076 205640 250128 205692
rect 323308 205640 323360 205692
rect 339684 205640 339736 205692
rect 339868 205640 339920 205692
rect 360292 205640 360344 205692
rect 360476 205640 360528 205692
rect 250168 205572 250220 205624
rect 323400 205504 323452 205556
rect 245844 202852 245896 202904
rect 245936 202852 245988 202904
rect 267740 202852 267792 202904
rect 267832 202852 267884 202904
rect 285956 202852 286008 202904
rect 286140 202852 286192 202904
rect 295524 202852 295576 202904
rect 295616 202852 295668 202904
rect 296812 202852 296864 202904
rect 296904 202852 296956 202904
rect 306748 202852 306800 202904
rect 306932 202852 306984 202904
rect 310888 202852 310940 202904
rect 324596 202852 324648 202904
rect 324688 202852 324740 202904
rect 325884 202852 325936 202904
rect 325976 202852 326028 202904
rect 341156 202852 341208 202904
rect 341248 202852 341300 202904
rect 358636 202852 358688 202904
rect 358728 202852 358780 202904
rect 359096 202852 359148 202904
rect 359188 202852 359240 202904
rect 362132 202852 362184 202904
rect 362224 202852 362276 202904
rect 389272 202852 389324 202904
rect 389548 202852 389600 202904
rect 421196 202852 421248 202904
rect 421380 202852 421432 202904
rect 424600 202852 424652 202904
rect 424876 202852 424928 202904
rect 463792 202852 463844 202904
rect 464068 202852 464120 202904
rect 470416 202852 470468 202904
rect 470600 202852 470652 202904
rect 299480 202827 299532 202836
rect 299480 202793 299489 202827
rect 299489 202793 299523 202827
rect 299523 202793 299532 202827
rect 299480 202784 299532 202793
rect 330116 202784 330168 202836
rect 336924 202827 336976 202836
rect 336924 202793 336933 202827
rect 336933 202793 336967 202827
rect 336967 202793 336976 202827
rect 336924 202784 336976 202793
rect 375840 202827 375892 202836
rect 375840 202793 375849 202827
rect 375849 202793 375883 202827
rect 375883 202793 375892 202827
rect 375840 202784 375892 202793
rect 265256 202759 265308 202768
rect 265256 202725 265265 202759
rect 265265 202725 265299 202759
rect 265299 202725 265308 202759
rect 265256 202716 265308 202725
rect 264980 201424 265032 201476
rect 265256 201424 265308 201476
rect 266636 201424 266688 201476
rect 266820 201424 266872 201476
rect 358728 201424 358780 201476
rect 421104 201424 421156 201476
rect 421196 201424 421248 201476
rect 244464 200175 244516 200184
rect 244464 200141 244473 200175
rect 244473 200141 244507 200175
rect 244507 200141 244516 200175
rect 244464 200132 244516 200141
rect 284668 200064 284720 200116
rect 284852 200064 284904 200116
rect 291660 200064 291712 200116
rect 317512 200064 317564 200116
rect 317696 200064 317748 200116
rect 284668 198679 284720 198688
rect 284668 198645 284677 198679
rect 284677 198645 284711 198679
rect 284711 198645 284720 198679
rect 284668 198636 284720 198645
rect 285772 198024 285824 198076
rect 285956 198024 286008 198076
rect 294236 198024 294288 198076
rect 294420 198024 294472 198076
rect 362224 198067 362276 198076
rect 362224 198033 362233 198067
rect 362233 198033 362267 198067
rect 362267 198033 362276 198067
rect 362224 198024 362276 198033
rect 290004 196596 290056 196648
rect 290188 196596 290240 196648
rect 262588 195984 262640 196036
rect 310888 196052 310940 196104
rect 389548 196052 389600 196104
rect 424692 195984 424744 196036
rect 424876 195984 424928 196036
rect 464068 196052 464120 196104
rect 262680 195916 262732 195968
rect 310796 195916 310848 195968
rect 389456 195916 389508 195968
rect 463976 195916 464028 195968
rect 236276 193332 236328 193384
rect 245844 193332 245896 193384
rect 236276 193196 236328 193248
rect 239128 193196 239180 193248
rect 239220 193196 239272 193248
rect 250076 193196 250128 193248
rect 250260 193196 250312 193248
rect 259736 193196 259788 193248
rect 259920 193196 259972 193248
rect 299480 193239 299532 193248
rect 299480 193205 299489 193239
rect 299489 193205 299523 193239
rect 299523 193205 299532 193239
rect 299480 193196 299532 193205
rect 302700 193264 302752 193316
rect 366824 193264 366876 193316
rect 367008 193264 367060 193316
rect 323308 193196 323360 193248
rect 323492 193196 323544 193248
rect 324596 193196 324648 193248
rect 324688 193196 324740 193248
rect 336924 193239 336976 193248
rect 336924 193205 336933 193239
rect 336933 193205 336967 193239
rect 336967 193205 336976 193239
rect 336924 193196 336976 193205
rect 337200 193196 337252 193248
rect 337384 193196 337436 193248
rect 341248 193196 341300 193248
rect 341432 193196 341484 193248
rect 357624 193196 357676 193248
rect 357716 193196 357768 193248
rect 359096 193196 359148 193248
rect 359188 193196 359240 193248
rect 362316 193196 362368 193248
rect 372528 193196 372580 193248
rect 372712 193196 372764 193248
rect 375840 193239 375892 193248
rect 375840 193205 375849 193239
rect 375849 193205 375883 193239
rect 375883 193205 375892 193239
rect 375840 193196 375892 193205
rect 376944 193196 376996 193248
rect 377128 193196 377180 193248
rect 245844 193128 245896 193180
rect 302516 193128 302568 193180
rect 367008 193171 367060 193180
rect 367008 193137 367017 193171
rect 367017 193137 367051 193171
rect 367051 193137 367060 193171
rect 367008 193128 367060 193137
rect 358636 191879 358688 191888
rect 358636 191845 358645 191879
rect 358645 191845 358679 191879
rect 358679 191845 358688 191879
rect 358636 191836 358688 191845
rect 239128 191768 239180 191820
rect 239404 191768 239456 191820
rect 251548 191768 251600 191820
rect 251640 191768 251692 191820
rect 324688 191768 324740 191820
rect 324872 191768 324924 191820
rect 288808 190476 288860 190528
rect 288900 190476 288952 190528
rect 291476 190519 291528 190528
rect 291476 190485 291485 190519
rect 291485 190485 291519 190519
rect 291519 190485 291528 190519
rect 291476 190476 291528 190485
rect 317512 190476 317564 190528
rect 317696 190476 317748 190528
rect 288808 190340 288860 190392
rect 288992 190340 289044 190392
rect 264980 189932 265032 189984
rect 265164 189932 265216 189984
rect 299848 188479 299900 188488
rect 299848 188445 299857 188479
rect 299857 188445 299891 188479
rect 299891 188445 299900 188479
rect 299848 188436 299900 188445
rect 306840 188479 306892 188488
rect 306840 188445 306849 188479
rect 306849 188445 306883 188479
rect 306883 188445 306892 188479
rect 306840 188436 306892 188445
rect 244464 186940 244516 186992
rect 267740 186371 267792 186380
rect 267740 186337 267749 186371
rect 267749 186337 267783 186371
rect 267783 186337 267792 186371
rect 267740 186328 267792 186337
rect 270684 186371 270736 186380
rect 270684 186337 270693 186371
rect 270693 186337 270727 186371
rect 270727 186337 270736 186371
rect 270684 186328 270736 186337
rect 295616 186396 295668 186448
rect 296904 186396 296956 186448
rect 325976 186396 326028 186448
rect 330116 186328 330168 186380
rect 295524 186260 295576 186312
rect 296812 186260 296864 186312
rect 325884 186260 325936 186312
rect 330116 186192 330168 186244
rect 285956 183676 286008 183728
rect 302516 183608 302568 183660
rect 267740 183583 267792 183592
rect 267740 183549 267749 183583
rect 267749 183549 267783 183583
rect 267783 183549 267792 183583
rect 267740 183540 267792 183549
rect 270684 183583 270736 183592
rect 270684 183549 270693 183583
rect 270693 183549 270727 183583
rect 270727 183549 270736 183583
rect 270684 183540 270736 183549
rect 272156 183540 272208 183592
rect 285956 183540 286008 183592
rect 294236 183540 294288 183592
rect 294420 183540 294472 183592
rect 299848 183583 299900 183592
rect 299848 183549 299857 183583
rect 299857 183549 299891 183583
rect 299891 183549 299900 183583
rect 299848 183540 299900 183549
rect 301044 183540 301096 183592
rect 301228 183540 301280 183592
rect 302608 183540 302660 183592
rect 306840 183583 306892 183592
rect 306840 183549 306849 183583
rect 306849 183549 306883 183583
rect 306883 183549 306892 183583
rect 306840 183540 306892 183549
rect 310888 183540 310940 183592
rect 311072 183540 311124 183592
rect 358636 183540 358688 183592
rect 358728 183540 358780 183592
rect 367008 183583 367060 183592
rect 367008 183549 367017 183583
rect 367017 183549 367051 183583
rect 367051 183549 367060 183583
rect 367008 183540 367060 183549
rect 389272 183540 389324 183592
rect 389548 183540 389600 183592
rect 424048 183540 424100 183592
rect 424692 183540 424744 183592
rect 463792 183540 463844 183592
rect 464068 183540 464120 183592
rect 470416 183540 470468 183592
rect 470600 183540 470652 183592
rect 272248 183472 272300 183524
rect 284668 183515 284720 183524
rect 284668 183481 284677 183515
rect 284677 183481 284711 183515
rect 284711 183481 284720 183515
rect 284668 183472 284720 183481
rect 337108 183515 337160 183524
rect 337108 183481 337117 183515
rect 337117 183481 337151 183515
rect 337151 183481 337160 183515
rect 337108 183472 337160 183481
rect 375840 183515 375892 183524
rect 375840 183481 375849 183515
rect 375849 183481 375883 183515
rect 375883 183481 375892 183515
rect 375840 183472 375892 183481
rect 424048 183447 424100 183456
rect 424048 183413 424057 183447
rect 424057 183413 424091 183447
rect 424091 183413 424100 183447
rect 424048 183404 424100 183413
rect 339684 182996 339736 183048
rect 339868 182996 339920 183048
rect 362224 182180 362276 182232
rect 362316 182180 362368 182232
rect 251456 182112 251508 182164
rect 251732 182112 251784 182164
rect 299848 182112 299900 182164
rect 299940 182112 299992 182164
rect 327356 182112 327408 182164
rect 327540 182112 327592 182164
rect 329932 182112 329984 182164
rect 330116 182112 330168 182164
rect 339500 182112 339552 182164
rect 339684 182112 339736 182164
rect 341156 182112 341208 182164
rect 341432 182112 341484 182164
rect 358544 182112 358596 182164
rect 358728 182112 358780 182164
rect 421196 182112 421248 182164
rect 421380 182112 421432 182164
rect 244372 180863 244424 180872
rect 244372 180829 244381 180863
rect 244381 180829 244415 180863
rect 244415 180829 244424 180863
rect 244372 180820 244424 180829
rect 251180 180752 251232 180804
rect 251456 180752 251508 180804
rect 265164 180752 265216 180804
rect 265256 180752 265308 180804
rect 284668 180795 284720 180804
rect 284668 180761 284677 180795
rect 284677 180761 284711 180795
rect 284711 180761 284720 180795
rect 284668 180752 284720 180761
rect 285956 180795 286008 180804
rect 285956 180761 285965 180795
rect 285965 180761 285999 180795
rect 285999 180761 286008 180795
rect 285956 180752 286008 180761
rect 288716 180795 288768 180804
rect 288716 180761 288725 180795
rect 288725 180761 288759 180795
rect 288759 180761 288768 180795
rect 288716 180752 288768 180761
rect 317512 180752 317564 180804
rect 317696 180752 317748 180804
rect 265256 179324 265308 179376
rect 359004 179367 359056 179376
rect 359004 179333 359013 179367
rect 359013 179333 359047 179367
rect 359047 179333 359056 179367
rect 359004 179324 359056 179333
rect 294236 178712 294288 178764
rect 294420 178712 294472 178764
rect 295524 178712 295576 178764
rect 295708 178712 295760 178764
rect 337200 178712 337252 178764
rect 289084 177828 289136 177880
rect 232228 176672 232280 176724
rect 301044 176672 301096 176724
rect 232320 176604 232372 176656
rect 302608 176740 302660 176792
rect 306840 176740 306892 176792
rect 310888 176740 310940 176792
rect 389548 176740 389600 176792
rect 463884 176672 463936 176724
rect 464068 176672 464120 176724
rect 302516 176604 302568 176656
rect 306748 176604 306800 176656
rect 310796 176604 310848 176656
rect 389456 176604 389508 176656
rect 301136 176536 301188 176588
rect 424232 176536 424284 176588
rect 285956 175967 286008 175976
rect 285956 175933 285965 175967
rect 285965 175933 285999 175967
rect 285999 175933 286008 175967
rect 285956 175924 286008 175933
rect 236276 173952 236328 174004
rect 266728 174020 266780 174072
rect 270500 173952 270552 174004
rect 270684 173952 270736 174004
rect 372620 173952 372672 174004
rect 372804 173952 372856 174004
rect 244372 173884 244424 173936
rect 244464 173884 244516 173936
rect 245844 173884 245896 173936
rect 245936 173884 245988 173936
rect 250076 173884 250128 173936
rect 250260 173884 250312 173936
rect 259644 173927 259696 173936
rect 259644 173893 259653 173927
rect 259653 173893 259687 173927
rect 259687 173893 259696 173927
rect 259644 173884 259696 173893
rect 262588 173884 262640 173936
rect 262680 173884 262732 173936
rect 266636 173884 266688 173936
rect 267832 173884 267884 173936
rect 267924 173884 267976 173936
rect 323308 173884 323360 173936
rect 323492 173884 323544 173936
rect 325884 173884 325936 173936
rect 325976 173884 326028 173936
rect 336740 173884 336792 173936
rect 336924 173884 336976 173936
rect 375840 173927 375892 173936
rect 375840 173893 375849 173927
rect 375849 173893 375883 173927
rect 375883 173893 375892 173927
rect 375840 173884 375892 173893
rect 376944 173884 376996 173936
rect 377128 173884 377180 173936
rect 236276 173816 236328 173868
rect 239128 172592 239180 172644
rect 239404 172592 239456 172644
rect 259644 172567 259696 172576
rect 259644 172533 259653 172567
rect 259653 172533 259687 172567
rect 259687 172533 259696 172567
rect 259644 172524 259696 172533
rect 296904 172456 296956 172508
rect 296996 172456 297048 172508
rect 324688 172456 324740 172508
rect 360292 171071 360344 171080
rect 360292 171037 360301 171071
rect 360301 171037 360335 171071
rect 360335 171037 360344 171071
rect 360292 171028 360344 171037
rect 362316 171028 362368 171080
rect 359096 169736 359148 169788
rect 289084 169711 289136 169720
rect 289084 169677 289093 169711
rect 289093 169677 289127 169711
rect 289127 169677 289136 169711
rect 289084 169668 289136 169677
rect 302516 169532 302568 169584
rect 302792 169532 302844 169584
rect 306748 169532 306800 169584
rect 307024 169532 307076 169584
rect 270500 169056 270552 169108
rect 270684 169056 270736 169108
rect 272156 167016 272208 167068
rect 310796 167016 310848 167068
rect 272248 166948 272300 167000
rect 424232 166948 424284 167000
rect 310888 166880 310940 166932
rect 424416 166880 424468 166932
rect 2780 165452 2832 165504
rect 5172 165452 5224 165504
rect 330116 164296 330168 164348
rect 330208 164296 330260 164348
rect 239128 164228 239180 164280
rect 244372 164160 244424 164212
rect 244556 164160 244608 164212
rect 372804 164203 372856 164212
rect 372804 164169 372813 164203
rect 372813 164169 372847 164203
rect 372847 164169 372856 164203
rect 372804 164160 372856 164169
rect 375840 164203 375892 164212
rect 375840 164169 375849 164203
rect 375849 164169 375883 164203
rect 375883 164169 375892 164203
rect 375840 164160 375892 164169
rect 376944 164160 376996 164212
rect 377128 164160 377180 164212
rect 424416 164160 424468 164212
rect 424508 164160 424560 164212
rect 463792 164160 463844 164212
rect 464068 164160 464120 164212
rect 239312 164092 239364 164144
rect 284668 162911 284720 162920
rect 284668 162877 284677 162911
rect 284677 162877 284711 162911
rect 284711 162877 284720 162911
rect 284668 162868 284720 162877
rect 294328 162868 294380 162920
rect 294420 162868 294472 162920
rect 324596 162911 324648 162920
rect 324596 162877 324605 162911
rect 324605 162877 324639 162911
rect 324639 162877 324648 162911
rect 324596 162868 324648 162877
rect 236276 162800 236328 162852
rect 236460 162800 236512 162852
rect 245844 162843 245896 162852
rect 245844 162809 245853 162843
rect 245853 162809 245887 162843
rect 245887 162809 245896 162843
rect 245844 162800 245896 162809
rect 250076 162800 250128 162852
rect 272064 162843 272116 162852
rect 272064 162809 272073 162843
rect 272073 162809 272107 162843
rect 272107 162809 272116 162843
rect 272064 162800 272116 162809
rect 302608 162800 302660 162852
rect 306748 162800 306800 162852
rect 306840 162800 306892 162852
rect 327172 162800 327224 162852
rect 327448 162800 327500 162852
rect 358636 162800 358688 162852
rect 358728 162800 358780 162852
rect 359004 162800 359056 162852
rect 359096 162800 359148 162852
rect 421196 162843 421248 162852
rect 421196 162809 421205 162843
rect 421205 162809 421239 162843
rect 421239 162809 421248 162843
rect 421196 162800 421248 162809
rect 239036 162732 239088 162784
rect 239312 162732 239364 162784
rect 250352 162732 250404 162784
rect 259552 161440 259604 161492
rect 259644 161440 259696 161492
rect 265164 161483 265216 161492
rect 265164 161449 265173 161483
rect 265173 161449 265207 161483
rect 265207 161449 265216 161483
rect 265164 161440 265216 161449
rect 360476 161440 360528 161492
rect 362224 161483 362276 161492
rect 362224 161449 362233 161483
rect 362233 161449 362267 161483
rect 362267 161449 362276 161483
rect 362224 161440 362276 161449
rect 250352 161415 250404 161424
rect 250352 161381 250361 161415
rect 250361 161381 250395 161415
rect 250395 161381 250404 161415
rect 250352 161372 250404 161381
rect 359096 161415 359148 161424
rect 359096 161381 359105 161415
rect 359105 161381 359139 161415
rect 359139 161381 359148 161415
rect 359096 161372 359148 161381
rect 289084 160123 289136 160132
rect 289084 160089 289093 160123
rect 289093 160089 289127 160123
rect 289127 160089 289136 160123
rect 289084 160080 289136 160089
rect 299756 159332 299808 159384
rect 299940 159332 299992 159384
rect 341064 159332 341116 159384
rect 341248 159332 341300 159384
rect 417884 157564 417936 157616
rect 418252 157564 418304 157616
rect 298008 157496 298060 157548
rect 306288 157496 306340 157548
rect 437204 157496 437256 157548
rect 437480 157496 437532 157548
rect 456524 157496 456576 157548
rect 456892 157496 456944 157548
rect 273536 157428 273588 157480
rect 307576 157428 307628 157480
rect 315948 157428 316000 157480
rect 267740 157360 267792 157412
rect 295524 157360 295576 157412
rect 295708 157360 295760 157412
rect 296812 157360 296864 157412
rect 296996 157360 297048 157412
rect 337108 157360 337160 157412
rect 273536 157292 273588 157344
rect 267740 157224 267792 157276
rect 325976 157224 326028 157276
rect 372804 157335 372856 157344
rect 372804 157301 372813 157335
rect 372813 157301 372847 157335
rect 372847 157301 372856 157335
rect 372804 157292 372856 157301
rect 337200 157224 337252 157276
rect 270684 157156 270736 157208
rect 270776 157088 270828 157140
rect 325976 157088 326028 157140
rect 375840 154615 375892 154624
rect 375840 154581 375849 154615
rect 375849 154581 375883 154615
rect 375883 154581 375892 154615
rect 375840 154572 375892 154581
rect 232320 154547 232372 154556
rect 232320 154513 232329 154547
rect 232329 154513 232363 154547
rect 232363 154513 232372 154547
rect 232320 154504 232372 154513
rect 272248 154504 272300 154556
rect 341064 154504 341116 154556
rect 341248 154504 341300 154556
rect 389456 154504 389508 154556
rect 389640 154504 389692 154556
rect 470416 154504 470468 154556
rect 470600 154504 470652 154556
rect 245936 154436 245988 154488
rect 301044 154436 301096 154488
rect 301228 154436 301280 154488
rect 302516 153255 302568 153264
rect 302516 153221 302525 153255
rect 302525 153221 302559 153255
rect 302559 153221 302568 153255
rect 302516 153212 302568 153221
rect 421196 153255 421248 153264
rect 421196 153221 421205 153255
rect 421205 153221 421239 153255
rect 421239 153221 421248 153255
rect 421196 153212 421248 153221
rect 245936 153187 245988 153196
rect 245936 153153 245945 153187
rect 245945 153153 245979 153187
rect 245979 153153 245988 153187
rect 245936 153144 245988 153153
rect 265164 153144 265216 153196
rect 265348 153144 265400 153196
rect 266636 153187 266688 153196
rect 266636 153153 266645 153187
rect 266645 153153 266679 153187
rect 266679 153153 266688 153187
rect 266636 153144 266688 153153
rect 285956 153144 286008 153196
rect 286048 153144 286100 153196
rect 310796 153187 310848 153196
rect 310796 153153 310805 153187
rect 310805 153153 310839 153187
rect 310839 153153 310848 153187
rect 310796 153144 310848 153153
rect 337200 153144 337252 153196
rect 302516 153076 302568 153128
rect 302792 153076 302844 153128
rect 250352 151827 250404 151836
rect 250352 151793 250361 151827
rect 250361 151793 250395 151827
rect 250395 151793 250404 151827
rect 250352 151784 250404 151793
rect 359188 151784 359240 151836
rect 3332 151716 3384 151768
rect 17224 151716 17276 151768
rect 288992 150356 289044 150408
rect 284668 147704 284720 147756
rect 284668 147568 284720 147620
rect 310796 147611 310848 147620
rect 310796 147577 310805 147611
rect 310805 147577 310839 147611
rect 310839 147577 310848 147611
rect 310796 147568 310848 147577
rect 232320 144959 232372 144968
rect 232320 144925 232329 144959
rect 232329 144925 232363 144959
rect 232363 144925 232372 144959
rect 232320 144916 232372 144925
rect 250352 144916 250404 144968
rect 250168 144848 250220 144900
rect 262588 144848 262640 144900
rect 262772 144848 262824 144900
rect 266636 144891 266688 144900
rect 266636 144857 266645 144891
rect 266645 144857 266679 144891
rect 266679 144857 266688 144891
rect 266636 144848 266688 144857
rect 267740 144848 267792 144900
rect 267924 144848 267976 144900
rect 270684 144848 270736 144900
rect 270960 144848 271012 144900
rect 272156 144848 272208 144900
rect 272432 144848 272484 144900
rect 273536 144891 273588 144900
rect 273536 144857 273545 144891
rect 273545 144857 273579 144891
rect 273579 144857 273588 144891
rect 273536 144848 273588 144857
rect 323308 144848 323360 144900
rect 323400 144848 323452 144900
rect 324596 144848 324648 144900
rect 324780 144848 324832 144900
rect 325884 144848 325936 144900
rect 326068 144848 326120 144900
rect 327172 144848 327224 144900
rect 327264 144848 327316 144900
rect 359188 144848 359240 144900
rect 359280 144848 359332 144900
rect 362132 144848 362184 144900
rect 362316 144848 362368 144900
rect 367008 144891 367060 144900
rect 367008 144857 367017 144891
rect 367017 144857 367051 144891
rect 367051 144857 367060 144891
rect 367008 144848 367060 144857
rect 375840 144891 375892 144900
rect 375840 144857 375849 144891
rect 375849 144857 375883 144891
rect 375883 144857 375892 144891
rect 375840 144848 375892 144857
rect 376944 144848 376996 144900
rect 377128 144848 377180 144900
rect 329932 144304 329984 144356
rect 330392 144304 330444 144356
rect 245936 143599 245988 143608
rect 245936 143565 245945 143599
rect 245945 143565 245979 143599
rect 245979 143565 245988 143599
rect 245936 143556 245988 143565
rect 337108 143599 337160 143608
rect 337108 143565 337117 143599
rect 337117 143565 337151 143599
rect 337151 143565 337160 143599
rect 337108 143556 337160 143565
rect 232320 143531 232372 143540
rect 232320 143497 232329 143531
rect 232329 143497 232363 143531
rect 232363 143497 232372 143531
rect 232320 143488 232372 143497
rect 244464 143531 244516 143540
rect 244464 143497 244473 143531
rect 244473 143497 244507 143531
rect 244507 143497 244516 143531
rect 244464 143488 244516 143497
rect 250168 143488 250220 143540
rect 250260 143488 250312 143540
rect 270960 143531 271012 143540
rect 270960 143497 270969 143531
rect 270969 143497 271003 143531
rect 271003 143497 271012 143531
rect 270960 143488 271012 143497
rect 272340 143488 272392 143540
rect 272432 143488 272484 143540
rect 302424 143488 302476 143540
rect 302608 143488 302660 143540
rect 323308 143488 323360 143540
rect 323492 143488 323544 143540
rect 327264 143531 327316 143540
rect 327264 143497 327273 143531
rect 327273 143497 327307 143531
rect 327307 143497 327316 143531
rect 327264 143488 327316 143497
rect 358728 143531 358780 143540
rect 358728 143497 358737 143531
rect 358737 143497 358771 143531
rect 358771 143497 358780 143531
rect 358728 143488 358780 143497
rect 362316 143488 362368 143540
rect 362500 143488 362552 143540
rect 421196 143531 421248 143540
rect 421196 143497 421205 143531
rect 421205 143497 421239 143531
rect 421239 143497 421248 143531
rect 421196 143488 421248 143497
rect 424140 142808 424192 142860
rect 424600 142808 424652 142860
rect 317512 142128 317564 142180
rect 317696 142128 317748 142180
rect 250260 142060 250312 142112
rect 259644 142103 259696 142112
rect 259644 142069 259653 142103
rect 259653 142069 259687 142103
rect 259687 142069 259696 142103
rect 259644 142060 259696 142069
rect 286140 142060 286192 142112
rect 296996 142060 297048 142112
rect 288808 140811 288860 140820
rect 288808 140777 288817 140811
rect 288817 140777 288851 140811
rect 288851 140777 288860 140811
rect 288808 140768 288860 140777
rect 295708 140743 295760 140752
rect 295708 140709 295717 140743
rect 295717 140709 295751 140743
rect 295751 140709 295760 140743
rect 295708 140700 295760 140709
rect 291568 139340 291620 139392
rect 291752 139340 291804 139392
rect 310888 138660 310940 138712
rect 372804 138116 372856 138168
rect 251456 138023 251508 138032
rect 251456 137989 251465 138023
rect 251465 137989 251499 138023
rect 251499 137989 251508 138023
rect 251456 137980 251508 137989
rect 301044 137980 301096 138032
rect 337108 137980 337160 138032
rect 389364 137980 389416 138032
rect 244464 137955 244516 137964
rect 244464 137921 244473 137955
rect 244473 137921 244507 137955
rect 244507 137921 244516 137955
rect 244464 137912 244516 137921
rect 273536 137955 273588 137964
rect 273536 137921 273545 137955
rect 273545 137921 273579 137955
rect 273579 137921 273588 137955
rect 273536 137912 273588 137921
rect 291752 137912 291804 137964
rect 301136 137912 301188 137964
rect 317512 137912 317564 137964
rect 317788 137912 317840 137964
rect 329932 137912 329984 137964
rect 330208 137912 330260 137964
rect 337200 137912 337252 137964
rect 389456 137912 389508 137964
rect 2780 136484 2832 136536
rect 5080 136484 5132 136536
rect 367008 135303 367060 135312
rect 367008 135269 367017 135303
rect 367017 135269 367051 135303
rect 367051 135269 367060 135303
rect 367008 135260 367060 135269
rect 372712 135303 372764 135312
rect 372712 135269 372721 135303
rect 372721 135269 372755 135303
rect 372755 135269 372764 135303
rect 372712 135260 372764 135269
rect 375840 135303 375892 135312
rect 375840 135269 375849 135303
rect 375849 135269 375883 135303
rect 375883 135269 375892 135303
rect 375840 135260 375892 135269
rect 239128 135192 239180 135244
rect 239312 135192 239364 135244
rect 267740 135192 267792 135244
rect 267832 135192 267884 135244
rect 324596 135192 324648 135244
rect 324688 135192 324740 135244
rect 327264 135235 327316 135244
rect 327264 135201 327273 135235
rect 327273 135201 327307 135235
rect 327307 135201 327316 135235
rect 327264 135192 327316 135201
rect 340880 135192 340932 135244
rect 341248 135192 341300 135244
rect 357440 135235 357492 135244
rect 357440 135201 357449 135235
rect 357449 135201 357483 135235
rect 357483 135201 357492 135235
rect 357440 135192 357492 135201
rect 470416 135192 470468 135244
rect 470600 135192 470652 135244
rect 270960 135099 271012 135108
rect 270960 135065 270969 135099
rect 270969 135065 271003 135099
rect 271003 135065 271012 135099
rect 270960 135056 271012 135065
rect 251456 133943 251508 133952
rect 251456 133909 251465 133943
rect 251465 133909 251499 133943
rect 251499 133909 251508 133943
rect 251456 133900 251508 133909
rect 358728 133943 358780 133952
rect 358728 133909 358737 133943
rect 358737 133909 358771 133943
rect 358771 133909 358780 133943
rect 421196 133943 421248 133952
rect 358728 133900 358780 133909
rect 421196 133909 421205 133943
rect 421205 133909 421239 133943
rect 421239 133909 421248 133943
rect 421196 133900 421248 133909
rect 337200 133875 337252 133884
rect 337200 133841 337209 133875
rect 337209 133841 337243 133875
rect 337243 133841 337252 133875
rect 337200 133832 337252 133841
rect 389456 133875 389508 133884
rect 389456 133841 389465 133875
rect 389465 133841 389499 133875
rect 389499 133841 389508 133875
rect 389456 133832 389508 133841
rect 249984 132515 250036 132524
rect 249984 132481 249993 132515
rect 249993 132481 250027 132515
rect 250027 132481 250036 132515
rect 249984 132472 250036 132481
rect 259736 132472 259788 132524
rect 286048 132515 286100 132524
rect 286048 132481 286057 132515
rect 286057 132481 286091 132515
rect 286091 132481 286100 132515
rect 286048 132472 286100 132481
rect 296904 132515 296956 132524
rect 296904 132481 296913 132515
rect 296913 132481 296947 132515
rect 296947 132481 296956 132515
rect 296904 132472 296956 132481
rect 299756 132472 299808 132524
rect 299848 132472 299900 132524
rect 302424 132472 302476 132524
rect 302608 132472 302660 132524
rect 284668 132447 284720 132456
rect 284668 132413 284677 132447
rect 284677 132413 284711 132447
rect 284711 132413 284720 132447
rect 284668 132404 284720 132413
rect 306748 132447 306800 132456
rect 306748 132413 306757 132447
rect 306757 132413 306791 132447
rect 306791 132413 306800 132447
rect 306748 132404 306800 132413
rect 288808 131180 288860 131232
rect 288716 131112 288768 131164
rect 295616 131112 295668 131164
rect 463884 130364 463936 130416
rect 464068 130364 464120 130416
rect 306840 129888 306892 129940
rect 325976 128392 326028 128444
rect 339684 128324 339736 128376
rect 339868 128324 339920 128376
rect 360292 128324 360344 128376
rect 360476 128324 360528 128376
rect 424140 128324 424192 128376
rect 424508 128324 424560 128376
rect 310796 128299 310848 128308
rect 310796 128265 310805 128299
rect 310805 128265 310839 128299
rect 310839 128265 310848 128299
rect 310796 128256 310848 128265
rect 325884 128256 325936 128308
rect 357532 128188 357584 128240
rect 232320 125715 232372 125724
rect 232320 125681 232329 125715
rect 232329 125681 232363 125715
rect 232363 125681 232372 125715
rect 232320 125672 232372 125681
rect 265164 125536 265216 125588
rect 265348 125536 265400 125588
rect 267740 125536 267792 125588
rect 267924 125536 267976 125588
rect 270684 125536 270736 125588
rect 270960 125536 271012 125588
rect 272156 125536 272208 125588
rect 272432 125536 272484 125588
rect 273536 125579 273588 125588
rect 273536 125545 273545 125579
rect 273545 125545 273579 125579
rect 273579 125545 273588 125579
rect 273536 125536 273588 125545
rect 323216 125536 323268 125588
rect 323400 125536 323452 125588
rect 324596 125536 324648 125588
rect 324780 125536 324832 125588
rect 325884 125536 325936 125588
rect 326068 125536 326120 125588
rect 327172 125536 327224 125588
rect 341064 125536 341116 125588
rect 357532 125536 357584 125588
rect 367008 125579 367060 125588
rect 367008 125545 367017 125579
rect 367017 125545 367051 125579
rect 367051 125545 367060 125579
rect 367008 125536 367060 125545
rect 310888 125468 310940 125520
rect 327264 125468 327316 125520
rect 357624 125468 357676 125520
rect 337292 124176 337344 124228
rect 232320 124151 232372 124160
rect 232320 124117 232329 124151
rect 232329 124117 232363 124151
rect 232363 124117 232372 124151
rect 232320 124108 232372 124117
rect 249984 124151 250036 124160
rect 249984 124117 249993 124151
rect 249993 124117 250027 124151
rect 250027 124117 250036 124151
rect 249984 124108 250036 124117
rect 272432 124108 272484 124160
rect 358728 124151 358780 124160
rect 358728 124117 358737 124151
rect 358737 124117 358771 124151
rect 358771 124117 358780 124151
rect 358728 124108 358780 124117
rect 421196 124151 421248 124160
rect 421196 124117 421205 124151
rect 421205 124117 421239 124151
rect 421239 124117 421248 124151
rect 421196 124108 421248 124117
rect 284852 122816 284904 122868
rect 290004 122816 290056 122868
rect 296904 122816 296956 122868
rect 297088 122816 297140 122868
rect 389180 122816 389232 122868
rect 290096 122680 290148 122732
rect 2780 122272 2832 122324
rect 4988 122272 5040 122324
rect 306840 121388 306892 121440
rect 330208 121388 330260 121440
rect 330576 121388 330628 121440
rect 324780 120572 324832 120624
rect 291568 120139 291620 120148
rect 291568 120105 291577 120139
rect 291577 120105 291611 120139
rect 291611 120105 291620 120139
rect 291568 120096 291620 120105
rect 330576 120071 330628 120080
rect 330576 120037 330585 120071
rect 330585 120037 330619 120071
rect 330619 120037 330628 120071
rect 330576 120028 330628 120037
rect 251456 118736 251508 118788
rect 299848 118736 299900 118788
rect 339868 118736 339920 118788
rect 337108 118668 337160 118720
rect 337292 118668 337344 118720
rect 377128 118668 377180 118720
rect 463884 118668 463936 118720
rect 251456 118600 251508 118652
rect 299848 118600 299900 118652
rect 341156 118643 341208 118652
rect 341156 118609 341165 118643
rect 341165 118609 341199 118643
rect 341199 118609 341208 118643
rect 341156 118600 341208 118609
rect 463976 118600 464028 118652
rect 377128 118532 377180 118584
rect 326068 118396 326120 118448
rect 326068 118260 326120 118312
rect 273536 115991 273588 116000
rect 273536 115957 273545 115991
rect 273545 115957 273579 115991
rect 273579 115957 273588 115991
rect 273536 115948 273588 115957
rect 339776 115991 339828 116000
rect 339776 115957 339785 115991
rect 339785 115957 339819 115991
rect 339819 115957 339828 115991
rect 339776 115948 339828 115957
rect 367008 115991 367060 116000
rect 367008 115957 367017 115991
rect 367017 115957 367051 115991
rect 367051 115957 367060 115991
rect 367008 115948 367060 115957
rect 270684 115880 270736 115932
rect 270960 115880 271012 115932
rect 341248 115880 341300 115932
rect 341432 115880 341484 115932
rect 377128 115880 377180 115932
rect 424600 115880 424652 115932
rect 424692 115880 424744 115932
rect 366824 115812 366876 115864
rect 367008 115812 367060 115864
rect 291568 115200 291620 115252
rect 310888 114588 310940 114640
rect 232320 114563 232372 114572
rect 232320 114529 232329 114563
rect 232329 114529 232363 114563
rect 232363 114529 232372 114563
rect 232320 114520 232372 114529
rect 250260 114520 250312 114572
rect 272156 114563 272208 114572
rect 272156 114529 272165 114563
rect 272165 114529 272199 114563
rect 272199 114529 272208 114563
rect 272156 114520 272208 114529
rect 358728 114563 358780 114572
rect 358728 114529 358737 114563
rect 358737 114529 358771 114563
rect 358771 114529 358780 114563
rect 358728 114520 358780 114529
rect 421196 114563 421248 114572
rect 421196 114529 421205 114563
rect 421205 114529 421239 114563
rect 421239 114529 421248 114563
rect 421196 114520 421248 114529
rect 267832 114495 267884 114504
rect 267832 114461 267841 114495
rect 267841 114461 267875 114495
rect 267875 114461 267884 114495
rect 267832 114452 267884 114461
rect 285956 114452 286008 114504
rect 286232 114452 286284 114504
rect 310796 114495 310848 114504
rect 310796 114461 310805 114495
rect 310805 114461 310839 114495
rect 310839 114461 310848 114495
rect 310796 114452 310848 114461
rect 424600 114452 424652 114504
rect 301044 113228 301096 113280
rect 259644 113160 259696 113212
rect 259736 113160 259788 113212
rect 296996 113160 297048 113212
rect 297088 113160 297140 113212
rect 301136 113160 301188 113212
rect 324596 113203 324648 113212
rect 324596 113169 324605 113203
rect 324605 113169 324639 113203
rect 324639 113169 324648 113203
rect 324596 113160 324648 113169
rect 299848 113092 299900 113144
rect 299940 113092 299992 113144
rect 306840 111843 306892 111852
rect 306840 111809 306849 111843
rect 306849 111809 306883 111843
rect 306883 111809 306892 111843
rect 306840 111800 306892 111809
rect 330576 111775 330628 111784
rect 330576 111741 330585 111775
rect 330585 111741 330619 111775
rect 330619 111741 330628 111775
rect 330576 111732 330628 111741
rect 368204 110644 368256 110696
rect 376668 110644 376720 110696
rect 456524 110644 456576 110696
rect 458824 110644 458876 110696
rect 414020 110576 414072 110628
rect 423496 110576 423548 110628
rect 437204 110576 437256 110628
rect 437480 110576 437532 110628
rect 347780 110508 347832 110560
rect 357348 110508 357400 110560
rect 324596 109692 324648 109744
rect 324596 109556 324648 109608
rect 266636 109012 266688 109064
rect 362224 109080 362276 109132
rect 463792 109012 463844 109064
rect 463976 109012 464028 109064
rect 266728 108944 266780 108996
rect 278780 108944 278832 108996
rect 279056 108944 279108 108996
rect 362132 108944 362184 108996
rect 330576 106700 330628 106752
rect 284852 106292 284904 106344
rect 358728 106335 358780 106344
rect 358728 106301 358737 106335
rect 358737 106301 358771 106335
rect 358771 106301 358780 106335
rect 358728 106292 358780 106301
rect 377036 106335 377088 106344
rect 377036 106301 377045 106335
rect 377045 106301 377079 106335
rect 377079 106301 377088 106335
rect 377036 106292 377088 106301
rect 236460 106224 236512 106276
rect 236644 106224 236696 106276
rect 239128 106224 239180 106276
rect 239312 106224 239364 106276
rect 259552 106224 259604 106276
rect 259828 106224 259880 106276
rect 270684 106224 270736 106276
rect 270960 106224 271012 106276
rect 272156 106224 272208 106276
rect 272432 106224 272484 106276
rect 273536 106267 273588 106276
rect 273536 106233 273545 106267
rect 273545 106233 273579 106267
rect 273579 106233 273588 106267
rect 273536 106224 273588 106233
rect 284760 106224 284812 106276
rect 375840 106267 375892 106276
rect 375840 106233 375849 106267
rect 375849 106233 375883 106267
rect 375883 106233 375892 106267
rect 375840 106224 375892 106233
rect 377128 106267 377180 106276
rect 377128 106233 377137 106267
rect 377137 106233 377171 106267
rect 377171 106233 377180 106267
rect 377128 106224 377180 106233
rect 358728 104975 358780 104984
rect 358728 104941 358737 104975
rect 358737 104941 358771 104975
rect 358771 104941 358780 104975
rect 358728 104932 358780 104941
rect 265256 104864 265308 104916
rect 265348 104864 265400 104916
rect 288808 104864 288860 104916
rect 288992 104864 289044 104916
rect 310888 104864 310940 104916
rect 424508 104907 424560 104916
rect 424508 104873 424517 104907
rect 424517 104873 424551 104907
rect 424551 104873 424560 104907
rect 424508 104864 424560 104873
rect 232320 104839 232372 104848
rect 232320 104805 232329 104839
rect 232329 104805 232363 104839
rect 232363 104805 232372 104839
rect 232320 104796 232372 104805
rect 295524 104796 295576 104848
rect 295616 104796 295668 104848
rect 302608 104839 302660 104848
rect 302608 104805 302617 104839
rect 302617 104805 302651 104839
rect 302651 104805 302660 104839
rect 302608 104796 302660 104805
rect 323400 104839 323452 104848
rect 323400 104805 323409 104839
rect 323409 104805 323443 104839
rect 323443 104805 323452 104839
rect 323400 104796 323452 104805
rect 324596 104839 324648 104848
rect 324596 104805 324605 104839
rect 324605 104805 324639 104839
rect 324639 104805 324648 104839
rect 324596 104796 324648 104805
rect 337292 104796 337344 104848
rect 339500 104796 339552 104848
rect 339776 104796 339828 104848
rect 358728 104796 358780 104848
rect 421196 104839 421248 104848
rect 421196 104805 421205 104839
rect 421205 104805 421239 104839
rect 421239 104805 421248 104839
rect 421196 104796 421248 104805
rect 291476 103547 291528 103556
rect 291476 103513 291485 103547
rect 291485 103513 291519 103547
rect 291519 103513 291528 103547
rect 291476 103504 291528 103513
rect 272432 103479 272484 103488
rect 272432 103445 272441 103479
rect 272441 103445 272475 103479
rect 272475 103445 272484 103479
rect 327172 103479 327224 103488
rect 272432 103436 272484 103445
rect 327172 103445 327181 103479
rect 327181 103445 327215 103479
rect 327215 103445 327224 103479
rect 327172 103436 327224 103445
rect 339500 103436 339552 103488
rect 330208 102187 330260 102196
rect 330208 102153 330217 102187
rect 330217 102153 330251 102187
rect 330251 102153 330260 102187
rect 330208 102144 330260 102153
rect 288808 102076 288860 102128
rect 294236 100036 294288 100088
rect 294420 100036 294472 100088
rect 244464 99424 244516 99476
rect 245936 99424 245988 99476
rect 310888 99424 310940 99476
rect 251456 99399 251508 99408
rect 251456 99365 251465 99399
rect 251465 99365 251499 99399
rect 251499 99365 251508 99399
rect 251456 99356 251508 99365
rect 278872 99356 278924 99408
rect 279056 99356 279108 99408
rect 424508 99356 424560 99408
rect 244464 99288 244516 99340
rect 245936 99288 245988 99340
rect 273536 99331 273588 99340
rect 273536 99297 273545 99331
rect 273545 99297 273579 99331
rect 273579 99297 273588 99331
rect 273536 99288 273588 99297
rect 310888 99288 310940 99340
rect 377128 99331 377180 99340
rect 377128 99297 377137 99331
rect 377137 99297 377171 99331
rect 377171 99297 377180 99331
rect 377128 99288 377180 99297
rect 424692 99288 424744 99340
rect 389456 99152 389508 99204
rect 327172 98719 327224 98728
rect 327172 98685 327181 98719
rect 327181 98685 327215 98719
rect 327215 98685 327224 98719
rect 327172 98676 327224 98685
rect 270500 98064 270552 98116
rect 270960 98064 271012 98116
rect 375840 97835 375892 97844
rect 375840 97801 375849 97835
rect 375849 97801 375883 97835
rect 375883 97801 375892 97835
rect 375840 97792 375892 97801
rect 330208 97248 330260 97300
rect 250076 96636 250128 96688
rect 250260 96636 250312 96688
rect 251456 96679 251508 96688
rect 251456 96645 251465 96679
rect 251465 96645 251499 96679
rect 251499 96645 251508 96679
rect 251456 96636 251508 96645
rect 367008 96611 367060 96620
rect 367008 96577 367017 96611
rect 367017 96577 367051 96611
rect 367051 96577 367060 96611
rect 367008 96568 367060 96577
rect 372620 96568 372672 96620
rect 372712 96568 372764 96620
rect 232320 95251 232372 95260
rect 232320 95217 232329 95251
rect 232329 95217 232363 95251
rect 232363 95217 232372 95251
rect 232320 95208 232372 95217
rect 285956 95208 286008 95260
rect 286048 95208 286100 95260
rect 302608 95251 302660 95260
rect 302608 95217 302617 95251
rect 302617 95217 302651 95251
rect 302651 95217 302660 95251
rect 302608 95208 302660 95217
rect 323400 95251 323452 95260
rect 323400 95217 323409 95251
rect 323409 95217 323443 95251
rect 323443 95217 323452 95251
rect 323400 95208 323452 95217
rect 324596 95251 324648 95260
rect 324596 95217 324605 95251
rect 324605 95217 324639 95251
rect 324639 95217 324648 95251
rect 324596 95208 324648 95217
rect 325884 95208 325936 95260
rect 325976 95208 326028 95260
rect 337200 95251 337252 95260
rect 337200 95217 337209 95251
rect 337209 95217 337243 95251
rect 337243 95217 337252 95251
rect 337200 95208 337252 95217
rect 339500 95208 339552 95260
rect 358636 95251 358688 95260
rect 358636 95217 358645 95251
rect 358645 95217 358679 95251
rect 358679 95217 358688 95251
rect 358636 95208 358688 95217
rect 266636 95183 266688 95192
rect 266636 95149 266645 95183
rect 266645 95149 266679 95183
rect 266679 95149 266688 95183
rect 266636 95140 266688 95149
rect 284760 95183 284812 95192
rect 284760 95149 284769 95183
rect 284769 95149 284803 95183
rect 284803 95149 284812 95183
rect 284760 95140 284812 95149
rect 310796 95183 310848 95192
rect 310796 95149 310805 95183
rect 310805 95149 310839 95183
rect 310839 95149 310848 95183
rect 310796 95140 310848 95149
rect 362316 95183 362368 95192
rect 362316 95149 362325 95183
rect 362325 95149 362359 95183
rect 362359 95149 362368 95183
rect 362316 95140 362368 95149
rect 267740 93848 267792 93900
rect 272340 93848 272392 93900
rect 284760 93891 284812 93900
rect 284760 93857 284769 93891
rect 284769 93857 284803 93891
rect 284803 93857 284812 93891
rect 284760 93848 284812 93857
rect 463700 93848 463752 93900
rect 463884 93848 463936 93900
rect 291476 93780 291528 93832
rect 306840 92556 306892 92608
rect 288716 92531 288768 92540
rect 288716 92497 288725 92531
rect 288725 92497 288759 92531
rect 288759 92497 288768 92531
rect 288716 92488 288768 92497
rect 306748 92488 306800 92540
rect 317788 89700 317840 89752
rect 424508 89700 424560 89752
rect 424692 89700 424744 89752
rect 317880 89564 317932 89616
rect 291384 88995 291436 89004
rect 291384 88961 291393 88995
rect 291393 88961 291427 88995
rect 291427 88961 291436 88995
rect 291384 88952 291436 88961
rect 389364 87907 389416 87916
rect 389364 87873 389373 87907
rect 389373 87873 389407 87907
rect 389407 87873 389416 87907
rect 389364 87864 389416 87873
rect 395896 87184 395948 87236
rect 395988 87184 396040 87236
rect 251180 87048 251232 87100
rect 260656 87048 260708 87100
rect 297548 87048 297600 87100
rect 306288 87048 306340 87100
rect 376760 87048 376812 87100
rect 386236 87048 386288 87100
rect 386420 87048 386472 87100
rect 395804 87048 395856 87100
rect 437204 87116 437256 87168
rect 437480 87116 437532 87168
rect 456524 87116 456576 87168
rect 456984 87116 457036 87168
rect 494612 87116 494664 87168
rect 502248 87116 502300 87168
rect 262588 86980 262640 87032
rect 262680 86980 262732 87032
rect 294420 86980 294472 87032
rect 347780 86980 347832 87032
rect 357348 86980 357400 87032
rect 367008 87023 367060 87032
rect 367008 86989 367017 87023
rect 367017 86989 367051 87023
rect 367051 86989 367060 87023
rect 367008 86980 367060 86989
rect 395896 86980 395948 87032
rect 395988 86980 396040 87032
rect 421196 87023 421248 87032
rect 421196 86989 421205 87023
rect 421205 86989 421239 87023
rect 421239 86989 421248 87023
rect 421196 86980 421248 86989
rect 251456 86955 251508 86964
rect 251456 86921 251465 86955
rect 251465 86921 251499 86955
rect 251499 86921 251508 86955
rect 251456 86912 251508 86921
rect 324596 86912 324648 86964
rect 327172 86912 327224 86964
rect 327264 86912 327316 86964
rect 336924 86912 336976 86964
rect 341156 86912 341208 86964
rect 294420 86844 294472 86896
rect 324688 86844 324740 86896
rect 336924 86776 336976 86828
rect 265256 85552 265308 85604
rect 265348 85552 265400 85604
rect 266728 85552 266780 85604
rect 267740 85552 267792 85604
rect 267832 85552 267884 85604
rect 272156 85552 272208 85604
rect 272340 85552 272392 85604
rect 299848 85552 299900 85604
rect 299940 85552 299992 85604
rect 301136 85552 301188 85604
rect 301228 85552 301280 85604
rect 306748 85552 306800 85604
rect 306840 85552 306892 85604
rect 310796 85595 310848 85604
rect 310796 85561 310805 85595
rect 310805 85561 310839 85595
rect 310839 85561 310848 85595
rect 310796 85552 310848 85561
rect 323032 85552 323084 85604
rect 323400 85552 323452 85604
rect 325884 85552 325936 85604
rect 325976 85552 326028 85604
rect 339500 85552 339552 85604
rect 339868 85552 339920 85604
rect 362408 85552 362460 85604
rect 232320 85484 232372 85536
rect 317880 85484 317932 85536
rect 360384 85484 360436 85536
rect 421196 85484 421248 85536
rect 266728 84167 266780 84176
rect 266728 84133 266737 84167
rect 266737 84133 266771 84167
rect 266771 84133 266780 84167
rect 266728 84124 266780 84133
rect 267832 84124 267884 84176
rect 284760 84124 284812 84176
rect 286048 84124 286100 84176
rect 288716 84167 288768 84176
rect 288716 84133 288725 84167
rect 288725 84133 288759 84167
rect 288759 84133 288768 84167
rect 288716 84124 288768 84133
rect 289912 84167 289964 84176
rect 289912 84133 289921 84167
rect 289921 84133 289955 84167
rect 289955 84133 289964 84167
rect 289912 84124 289964 84133
rect 296996 84167 297048 84176
rect 296996 84133 297005 84167
rect 297005 84133 297039 84167
rect 297039 84133 297048 84167
rect 296996 84124 297048 84133
rect 306840 84124 306892 84176
rect 330300 82900 330352 82952
rect 357716 80112 357768 80164
rect 303896 80044 303948 80096
rect 357624 80044 357676 80096
rect 372896 80112 372948 80164
rect 389364 80044 389416 80096
rect 463792 80044 463844 80096
rect 372712 79976 372764 80028
rect 375840 79976 375892 80028
rect 377128 79976 377180 80028
rect 303896 79908 303948 79960
rect 375932 79908 375984 79960
rect 377220 79908 377272 79960
rect 389456 79908 389508 79960
rect 463792 79908 463844 79960
rect 2780 79772 2832 79824
rect 4896 79772 4948 79824
rect 250076 77392 250128 77444
rect 236276 77256 236328 77308
rect 236460 77256 236512 77308
rect 249984 77256 250036 77308
rect 301228 77367 301280 77376
rect 301228 77333 301237 77367
rect 301237 77333 301271 77367
rect 301271 77333 301280 77367
rect 301228 77324 301280 77333
rect 251456 77299 251508 77308
rect 251456 77265 251465 77299
rect 251465 77265 251499 77299
rect 251499 77265 251508 77299
rect 251456 77256 251508 77265
rect 262588 77256 262640 77308
rect 262680 77256 262732 77308
rect 299756 77256 299808 77308
rect 299848 77256 299900 77308
rect 302516 77256 302568 77308
rect 302608 77256 302660 77308
rect 341064 77299 341116 77308
rect 341064 77265 341073 77299
rect 341073 77265 341107 77299
rect 341107 77265 341116 77299
rect 341064 77256 341116 77265
rect 303896 77188 303948 77240
rect 303988 77188 304040 77240
rect 389456 77188 389508 77240
rect 341064 77163 341116 77172
rect 341064 77129 341073 77163
rect 341073 77129 341107 77163
rect 341107 77129 341116 77163
rect 341064 77120 341116 77129
rect 294236 76440 294288 76492
rect 294420 76440 294472 76492
rect 367100 76168 367152 76220
rect 376668 76168 376720 76220
rect 396080 76032 396132 76084
rect 399392 76032 399444 76084
rect 437204 76032 437256 76084
rect 437480 76032 437532 76084
rect 456524 76032 456576 76084
rect 456800 76032 456852 76084
rect 232228 75939 232280 75948
rect 232228 75905 232237 75939
rect 232237 75905 232271 75939
rect 232271 75905 232280 75939
rect 232228 75896 232280 75905
rect 270500 75896 270552 75948
rect 270684 75896 270736 75948
rect 306380 75896 306432 75948
rect 311256 75896 311308 75948
rect 317696 75939 317748 75948
rect 317696 75905 317705 75939
rect 317705 75905 317739 75939
rect 317739 75905 317748 75939
rect 317696 75896 317748 75905
rect 323032 75896 323084 75948
rect 323308 75896 323360 75948
rect 358728 75896 358780 75948
rect 359004 75896 359056 75948
rect 360200 75939 360252 75948
rect 360200 75905 360209 75939
rect 360209 75905 360243 75939
rect 360243 75905 360252 75939
rect 360200 75896 360252 75905
rect 362224 75896 362276 75948
rect 362408 75896 362460 75948
rect 421012 75939 421064 75948
rect 421012 75905 421021 75939
rect 421021 75905 421055 75939
rect 421055 75905 421064 75939
rect 421012 75896 421064 75905
rect 301228 75871 301280 75880
rect 301228 75837 301237 75871
rect 301237 75837 301271 75871
rect 301271 75837 301280 75871
rect 301228 75828 301280 75837
rect 310796 75871 310848 75880
rect 310796 75837 310805 75871
rect 310805 75837 310839 75871
rect 310839 75837 310848 75871
rect 310796 75828 310848 75837
rect 330208 75871 330260 75880
rect 330208 75837 330217 75871
rect 330217 75837 330251 75871
rect 330251 75837 330260 75871
rect 330208 75828 330260 75837
rect 288900 75760 288952 75812
rect 306748 75803 306800 75812
rect 306748 75769 306757 75803
rect 306757 75769 306791 75803
rect 306791 75769 306800 75803
rect 306748 75760 306800 75769
rect 266820 74536 266872 74588
rect 267740 74579 267792 74588
rect 267740 74545 267749 74579
rect 267749 74545 267783 74579
rect 267783 74545 267792 74579
rect 267740 74536 267792 74545
rect 290004 74536 290056 74588
rect 296904 74536 296956 74588
rect 359096 74536 359148 74588
rect 359188 74536 359240 74588
rect 362224 74468 362276 74520
rect 362408 74468 362460 74520
rect 296904 74400 296956 74452
rect 272248 72428 272300 72480
rect 357624 70499 357676 70508
rect 357624 70465 357633 70499
rect 357633 70465 357667 70499
rect 357667 70465 357676 70499
rect 357624 70456 357676 70465
rect 341156 70252 341208 70304
rect 330208 69955 330260 69964
rect 330208 69921 330217 69955
rect 330217 69921 330251 69955
rect 330251 69921 330260 69955
rect 330208 69912 330260 69921
rect 302516 67668 302568 67720
rect 272156 67643 272208 67652
rect 272156 67609 272165 67643
rect 272165 67609 272199 67643
rect 272199 67609 272208 67643
rect 272156 67600 272208 67609
rect 302424 67600 302476 67652
rect 325884 67600 325936 67652
rect 325976 67600 326028 67652
rect 389364 67643 389416 67652
rect 389364 67609 389373 67643
rect 389373 67609 389407 67643
rect 389407 67609 389416 67643
rect 389364 67600 389416 67609
rect 236276 67575 236328 67584
rect 236276 67541 236285 67575
rect 236285 67541 236319 67575
rect 236319 67541 236328 67575
rect 236276 67532 236328 67541
rect 273628 67575 273680 67584
rect 273628 67541 273637 67575
rect 273637 67541 273671 67575
rect 273671 67541 273680 67575
rect 273628 67532 273680 67541
rect 270684 66308 270736 66360
rect 310796 66351 310848 66360
rect 310796 66317 310805 66351
rect 310805 66317 310839 66351
rect 310839 66317 310848 66351
rect 310796 66308 310848 66317
rect 266636 66240 266688 66292
rect 266820 66240 266872 66292
rect 270776 66240 270828 66292
rect 284668 66283 284720 66292
rect 284668 66249 284677 66283
rect 284677 66249 284711 66283
rect 284711 66249 284720 66283
rect 284668 66240 284720 66249
rect 285956 66283 286008 66292
rect 285956 66249 285965 66283
rect 285965 66249 285999 66283
rect 285999 66249 286008 66283
rect 285956 66240 286008 66249
rect 301044 66240 301096 66292
rect 301228 66240 301280 66292
rect 306656 66240 306708 66292
rect 306748 66240 306800 66292
rect 357624 66283 357676 66292
rect 357624 66249 357633 66283
rect 357633 66249 357667 66283
rect 357667 66249 357676 66283
rect 357624 66240 357676 66249
rect 232320 66172 232372 66224
rect 250076 66215 250128 66224
rect 250076 66181 250085 66215
rect 250085 66181 250119 66215
rect 250119 66181 250128 66215
rect 250076 66172 250128 66181
rect 265164 66172 265216 66224
rect 310796 66215 310848 66224
rect 310796 66181 310805 66215
rect 310805 66181 310839 66215
rect 310839 66181 310848 66215
rect 310796 66172 310848 66181
rect 325884 66172 325936 66224
rect 327172 66215 327224 66224
rect 327172 66181 327181 66215
rect 327181 66181 327215 66215
rect 327215 66181 327224 66215
rect 327172 66172 327224 66181
rect 336924 66215 336976 66224
rect 336924 66181 336933 66215
rect 336933 66181 336967 66215
rect 336967 66181 336976 66215
rect 336924 66172 336976 66181
rect 421196 66172 421248 66224
rect 296812 64923 296864 64932
rect 296812 64889 296821 64923
rect 296821 64889 296855 64923
rect 296855 64889 296864 64923
rect 296812 64880 296864 64889
rect 3332 64812 3384 64864
rect 24124 64812 24176 64864
rect 267740 64855 267792 64864
rect 267740 64821 267749 64855
rect 267749 64821 267783 64855
rect 267783 64821 267792 64855
rect 294236 64855 294288 64864
rect 267740 64812 267792 64821
rect 294236 64821 294245 64855
rect 294245 64821 294279 64855
rect 294279 64821 294288 64855
rect 294236 64812 294288 64821
rect 324872 64812 324924 64864
rect 324964 64812 325016 64864
rect 359096 64855 359148 64864
rect 359096 64821 359105 64855
rect 359105 64821 359139 64855
rect 359139 64821 359148 64855
rect 359096 64812 359148 64821
rect 362500 64812 362552 64864
rect 414020 63724 414072 63776
rect 418896 63724 418948 63776
rect 437204 63656 437256 63708
rect 437480 63656 437532 63708
rect 456524 63656 456576 63708
rect 456892 63656 456944 63708
rect 266636 61455 266688 61464
rect 266636 61421 266645 61455
rect 266645 61421 266679 61455
rect 266679 61421 266688 61455
rect 266636 61412 266688 61421
rect 323308 61455 323360 61464
rect 323308 61421 323317 61455
rect 323317 61421 323351 61455
rect 323351 61421 323360 61455
rect 323308 61412 323360 61421
rect 250076 60707 250128 60716
rect 250076 60673 250085 60707
rect 250085 60673 250119 60707
rect 250119 60673 250128 60707
rect 250076 60664 250128 60673
rect 259644 60664 259696 60716
rect 259828 60664 259880 60716
rect 262588 60664 262640 60716
rect 262772 60664 262824 60716
rect 339684 60664 339736 60716
rect 339868 60664 339920 60716
rect 341156 60664 341208 60716
rect 341340 60664 341392 60716
rect 360292 60664 360344 60716
rect 360476 60664 360528 60716
rect 306656 59984 306708 60036
rect 311072 59984 311124 60036
rect 272156 58012 272208 58064
rect 236276 57987 236328 57996
rect 236276 57953 236285 57987
rect 236285 57953 236319 57987
rect 236319 57953 236328 57987
rect 236276 57944 236328 57953
rect 273628 57987 273680 57996
rect 273628 57953 273637 57987
rect 273637 57953 273671 57987
rect 273671 57953 273680 57987
rect 273628 57944 273680 57953
rect 299756 57944 299808 57996
rect 299848 57944 299900 57996
rect 302424 57944 302476 57996
rect 302516 57944 302568 57996
rect 303896 57944 303948 57996
rect 303988 57944 304040 57996
rect 245568 57876 245620 57928
rect 245936 57876 245988 57928
rect 272156 57876 272208 57928
rect 290004 57876 290056 57928
rect 290096 57876 290148 57928
rect 291476 57876 291528 57928
rect 291568 57876 291620 57928
rect 301044 57919 301096 57928
rect 301044 57885 301053 57919
rect 301053 57885 301087 57919
rect 301087 57885 301096 57919
rect 301044 57876 301096 57885
rect 339868 57876 339920 57928
rect 367008 57919 367060 57928
rect 367008 57885 367017 57919
rect 367017 57885 367051 57919
rect 367051 57885 367060 57919
rect 367008 57876 367060 57885
rect 389180 57919 389232 57928
rect 389180 57885 389189 57919
rect 389189 57885 389223 57919
rect 389223 57885 389232 57919
rect 389180 57876 389232 57885
rect 470600 57919 470652 57928
rect 470600 57885 470609 57919
rect 470609 57885 470643 57919
rect 470643 57885 470652 57919
rect 470600 57876 470652 57885
rect 284668 57035 284720 57044
rect 284668 57001 284677 57035
rect 284677 57001 284711 57035
rect 284711 57001 284720 57035
rect 284668 56992 284720 57001
rect 421104 56695 421156 56704
rect 421104 56661 421113 56695
rect 421113 56661 421147 56695
rect 421147 56661 421156 56695
rect 421104 56652 421156 56661
rect 327264 56584 327316 56636
rect 336924 56627 336976 56636
rect 336924 56593 336933 56627
rect 336933 56593 336967 56627
rect 336967 56593 336976 56627
rect 336924 56584 336976 56593
rect 286048 56559 286100 56568
rect 286048 56525 286057 56559
rect 286057 56525 286091 56559
rect 286091 56525 286100 56559
rect 337292 56559 337344 56568
rect 286048 56516 286100 56525
rect 337292 56525 337301 56559
rect 337301 56525 337335 56559
rect 337335 56525 337344 56559
rect 337292 56516 337344 56525
rect 359096 56559 359148 56568
rect 359096 56525 359105 56559
rect 359105 56525 359139 56559
rect 359139 56525 359148 56559
rect 359096 56516 359148 56525
rect 421104 56516 421156 56568
rect 268108 55224 268160 55276
rect 294236 55267 294288 55276
rect 294236 55233 294245 55267
rect 294245 55233 294279 55267
rect 294279 55233 294288 55267
rect 294236 55224 294288 55233
rect 317512 55224 317564 55276
rect 317696 55224 317748 55276
rect 362224 55267 362276 55276
rect 362224 55233 362233 55267
rect 362233 55233 362267 55267
rect 362267 55233 362276 55267
rect 362224 55224 362276 55233
rect 424508 53839 424560 53848
rect 424508 53805 424517 53839
rect 424517 53805 424551 53839
rect 424551 53805 424560 53839
rect 424508 53796 424560 53805
rect 262588 52232 262640 52284
rect 262772 52232 262824 52284
rect 307024 51960 307076 52012
rect 301044 51799 301096 51808
rect 301044 51765 301053 51799
rect 301053 51765 301087 51799
rect 301087 51765 301096 51799
rect 301044 51756 301096 51765
rect 244464 51076 244516 51128
rect 244372 51008 244424 51060
rect 250076 50983 250128 50992
rect 250076 50949 250085 50983
rect 250085 50949 250119 50983
rect 250119 50949 250128 50983
rect 250076 50940 250128 50949
rect 2780 50464 2832 50516
rect 4804 50464 4856 50516
rect 232228 48331 232280 48340
rect 232228 48297 232237 48331
rect 232237 48297 232271 48331
rect 232271 48297 232280 48331
rect 232228 48288 232280 48297
rect 250076 48331 250128 48340
rect 250076 48297 250085 48331
rect 250085 48297 250119 48331
rect 250119 48297 250128 48331
rect 250076 48288 250128 48297
rect 266636 48331 266688 48340
rect 266636 48297 266645 48331
rect 266645 48297 266679 48331
rect 266679 48297 266688 48331
rect 266636 48288 266688 48297
rect 284760 48288 284812 48340
rect 323308 48331 323360 48340
rect 323308 48297 323317 48331
rect 323317 48297 323351 48331
rect 323351 48297 323360 48331
rect 323308 48288 323360 48297
rect 339776 48331 339828 48340
rect 339776 48297 339785 48331
rect 339785 48297 339819 48331
rect 339819 48297 339828 48331
rect 339776 48288 339828 48297
rect 358636 48288 358688 48340
rect 358728 48288 358780 48340
rect 367008 48331 367060 48340
rect 367008 48297 367017 48331
rect 367017 48297 367051 48331
rect 367051 48297 367060 48331
rect 367008 48288 367060 48297
rect 389272 48288 389324 48340
rect 424692 48288 424744 48340
rect 470600 48331 470652 48340
rect 470600 48297 470609 48331
rect 470609 48297 470643 48331
rect 470643 48297 470652 48331
rect 470600 48288 470652 48297
rect 236276 48263 236328 48272
rect 236276 48229 236285 48263
rect 236285 48229 236319 48263
rect 236319 48229 236328 48263
rect 236276 48220 236328 48229
rect 273536 48263 273588 48272
rect 273536 48229 273545 48263
rect 273545 48229 273579 48263
rect 273579 48229 273588 48263
rect 273536 48220 273588 48229
rect 326068 48152 326120 48204
rect 265256 46971 265308 46980
rect 265256 46937 265265 46971
rect 265265 46937 265299 46971
rect 265299 46937 265308 46971
rect 265256 46928 265308 46937
rect 285956 46928 286008 46980
rect 337108 46928 337160 46980
rect 421012 46971 421064 46980
rect 421012 46937 421021 46971
rect 421021 46937 421055 46971
rect 421055 46937 421064 46971
rect 421012 46928 421064 46937
rect 234988 46903 235040 46912
rect 234988 46869 234997 46903
rect 234997 46869 235031 46903
rect 235031 46869 235040 46903
rect 234988 46860 235040 46869
rect 259644 46860 259696 46912
rect 259736 46860 259788 46912
rect 301044 46860 301096 46912
rect 301320 46860 301372 46912
rect 302516 46860 302568 46912
rect 302608 46860 302660 46912
rect 327264 46903 327316 46912
rect 327264 46869 327273 46903
rect 327273 46869 327307 46903
rect 327307 46869 327316 46903
rect 327264 46860 327316 46869
rect 330116 46903 330168 46912
rect 330116 46869 330125 46903
rect 330125 46869 330159 46903
rect 330159 46869 330168 46903
rect 330116 46860 330168 46869
rect 336924 46903 336976 46912
rect 336924 46869 336933 46903
rect 336933 46869 336967 46903
rect 336967 46869 336976 46903
rect 336924 46860 336976 46869
rect 341432 46860 341484 46912
rect 358728 46860 358780 46912
rect 359096 46903 359148 46912
rect 359096 46869 359105 46903
rect 359105 46869 359139 46903
rect 359139 46869 359148 46903
rect 359096 46860 359148 46869
rect 268108 45908 268160 45960
rect 310888 45636 310940 45688
rect 311072 45636 311124 45688
rect 267832 45611 267884 45620
rect 267832 45577 267841 45611
rect 267841 45577 267875 45611
rect 267875 45577 267884 45611
rect 267832 45568 267884 45577
rect 265256 45543 265308 45552
rect 265256 45509 265265 45543
rect 265265 45509 265299 45543
rect 265299 45509 265308 45543
rect 265256 45500 265308 45509
rect 290096 45500 290148 45552
rect 291568 45500 291620 45552
rect 296812 45543 296864 45552
rect 296812 45509 296821 45543
rect 296821 45509 296855 45543
rect 296855 45509 296864 45543
rect 296812 45500 296864 45509
rect 301320 45543 301372 45552
rect 301320 45509 301329 45543
rect 301329 45509 301363 45543
rect 301363 45509 301372 45543
rect 301320 45500 301372 45509
rect 307024 45543 307076 45552
rect 307024 45509 307033 45543
rect 307033 45509 307067 45543
rect 307067 45509 307076 45543
rect 307024 45500 307076 45509
rect 310888 45500 310940 45552
rect 311072 45500 311124 45552
rect 317512 45500 317564 45552
rect 317696 45500 317748 45552
rect 288808 45432 288860 45484
rect 289084 45432 289136 45484
rect 290188 45432 290240 45484
rect 291660 45432 291712 45484
rect 299756 42032 299808 42084
rect 300124 42032 300176 42084
rect 421012 42032 421064 42084
rect 251456 41420 251508 41472
rect 284760 41420 284812 41472
rect 362224 41463 362276 41472
rect 362224 41429 362233 41463
rect 362233 41429 362267 41463
rect 362267 41429 362276 41463
rect 362224 41420 362276 41429
rect 251364 41352 251416 41404
rect 284668 41352 284720 41404
rect 360292 41352 360344 41404
rect 360476 41352 360528 41404
rect 388996 41352 389048 41404
rect 389364 41352 389416 41404
rect 239128 41327 239180 41336
rect 239128 41293 239137 41327
rect 239137 41293 239171 41327
rect 239171 41293 239180 41327
rect 239128 41284 239180 41293
rect 377128 41327 377180 41336
rect 377128 41293 377137 41327
rect 377137 41293 377171 41327
rect 377171 41293 377180 41327
rect 377128 41284 377180 41293
rect 396080 40196 396132 40248
rect 399024 40196 399076 40248
rect 437204 40196 437256 40248
rect 437480 40196 437532 40248
rect 303804 40171 303856 40180
rect 303804 40137 303813 40171
rect 303813 40137 303847 40171
rect 303847 40137 303856 40171
rect 303804 40128 303856 40137
rect 306380 40128 306432 40180
rect 315948 40128 316000 40180
rect 417884 40128 417936 40180
rect 418252 40128 418304 40180
rect 456524 40128 456576 40180
rect 456892 40128 456944 40180
rect 232320 38700 232372 38752
rect 232412 38700 232464 38752
rect 244372 38700 244424 38752
rect 377036 38700 377088 38752
rect 244464 38632 244516 38684
rect 245568 38632 245620 38684
rect 245936 38632 245988 38684
rect 270684 38632 270736 38684
rect 270776 38632 270828 38684
rect 272156 38632 272208 38684
rect 272248 38632 272300 38684
rect 273536 38675 273588 38684
rect 273536 38641 273545 38675
rect 273545 38641 273579 38675
rect 273579 38641 273588 38675
rect 273536 38632 273588 38641
rect 323308 38632 323360 38684
rect 296812 38607 296864 38616
rect 296812 38573 296821 38607
rect 296821 38573 296855 38607
rect 296855 38573 296864 38607
rect 296812 38564 296864 38573
rect 362224 38607 362276 38616
rect 362224 38573 362233 38607
rect 362233 38573 362267 38607
rect 362267 38573 362276 38607
rect 362224 38564 362276 38573
rect 367008 38607 367060 38616
rect 367008 38573 367017 38607
rect 367017 38573 367051 38607
rect 367051 38573 367060 38607
rect 367008 38564 367060 38573
rect 424508 38607 424560 38616
rect 424508 38573 424517 38607
rect 424517 38573 424551 38607
rect 424551 38573 424560 38607
rect 424508 38564 424560 38573
rect 323400 38496 323452 38548
rect 235080 37272 235132 37324
rect 236276 37315 236328 37324
rect 236276 37281 236285 37315
rect 236285 37281 236319 37315
rect 236319 37281 236328 37315
rect 236276 37272 236328 37281
rect 239128 37315 239180 37324
rect 239128 37281 239137 37315
rect 239137 37281 239171 37315
rect 239171 37281 239180 37315
rect 239128 37272 239180 37281
rect 325976 37272 326028 37324
rect 326068 37272 326120 37324
rect 327264 37315 327316 37324
rect 327264 37281 327273 37315
rect 327273 37281 327307 37315
rect 327307 37281 327316 37315
rect 327264 37272 327316 37281
rect 330116 37315 330168 37324
rect 330116 37281 330125 37315
rect 330125 37281 330159 37315
rect 330159 37281 330168 37315
rect 330116 37272 330168 37281
rect 336924 37315 336976 37324
rect 336924 37281 336933 37315
rect 336933 37281 336967 37315
rect 336967 37281 336976 37315
rect 336924 37272 336976 37281
rect 341248 37315 341300 37324
rect 341248 37281 341257 37315
rect 341257 37281 341291 37315
rect 341291 37281 341300 37315
rect 341248 37272 341300 37281
rect 357532 37272 357584 37324
rect 357716 37272 357768 37324
rect 358636 37315 358688 37324
rect 358636 37281 358645 37315
rect 358645 37281 358679 37315
rect 358679 37281 358688 37315
rect 358636 37272 358688 37281
rect 359188 37272 359240 37324
rect 244464 37204 244516 37256
rect 245936 37204 245988 37256
rect 267832 37204 267884 37256
rect 268016 37204 268068 37256
rect 337200 37204 337252 37256
rect 265256 35955 265308 35964
rect 265256 35921 265265 35955
rect 265265 35921 265299 35955
rect 265299 35921 265308 35955
rect 265256 35912 265308 35921
rect 294144 35912 294196 35964
rect 294236 35912 294288 35964
rect 301320 35955 301372 35964
rect 301320 35921 301329 35955
rect 301329 35921 301363 35955
rect 301363 35921 301372 35955
rect 301320 35912 301372 35921
rect 307024 35955 307076 35964
rect 307024 35921 307033 35955
rect 307033 35921 307067 35955
rect 307067 35921 307076 35955
rect 307024 35912 307076 35921
rect 3148 35844 3200 35896
rect 6184 35844 6236 35896
rect 336740 33804 336792 33856
rect 336924 33804 336976 33856
rect 303896 32376 303948 32428
rect 377128 31968 377180 32020
rect 377312 31968 377364 32020
rect 265256 31764 265308 31816
rect 317512 31764 317564 31816
rect 317696 31764 317748 31816
rect 327264 31764 327316 31816
rect 265256 31628 265308 31680
rect 389364 31696 389416 31748
rect 389548 31696 389600 31748
rect 266636 31560 266688 31612
rect 266820 31560 266872 31612
rect 327264 31560 327316 31612
rect 289084 29792 289136 29844
rect 267740 29180 267792 29232
rect 277308 29180 277360 29232
rect 456524 29180 456576 29232
rect 456984 29180 457036 29232
rect 238760 29112 238812 29164
rect 256608 29112 256660 29164
rect 437204 29112 437256 29164
rect 437480 29112 437532 29164
rect 286048 29044 286100 29096
rect 347780 29044 347832 29096
rect 357348 29044 357400 29096
rect 359188 29044 359240 29096
rect 367008 29087 367060 29096
rect 367008 29053 367017 29087
rect 367017 29053 367051 29087
rect 367051 29053 367060 29087
rect 367008 29044 367060 29053
rect 492772 29044 492824 29096
rect 502248 29044 502300 29096
rect 232228 28976 232280 29028
rect 232412 28976 232464 29028
rect 284668 28976 284720 29028
rect 284760 28976 284812 29028
rect 285956 28976 286008 29028
rect 325976 28976 326028 29028
rect 326068 28976 326120 29028
rect 358636 28976 358688 29028
rect 358728 28976 358780 29028
rect 424600 28976 424652 29028
rect 295524 28908 295576 28960
rect 295616 28908 295668 28960
rect 323308 28908 323360 28960
rect 323400 28908 323452 28960
rect 324596 28908 324648 28960
rect 324688 28908 324740 28960
rect 359188 28908 359240 28960
rect 367008 28951 367060 28960
rect 367008 28917 367017 28951
rect 367017 28917 367051 28951
rect 367051 28917 367060 28951
rect 367008 28908 367060 28917
rect 389548 28908 389600 28960
rect 306380 28772 306432 28824
rect 315948 28772 316000 28824
rect 244372 28067 244424 28076
rect 244372 28033 244381 28067
rect 244381 28033 244415 28067
rect 244415 28033 244424 28067
rect 244372 28024 244424 28033
rect 245844 27659 245896 27668
rect 245844 27625 245853 27659
rect 245853 27625 245887 27659
rect 245887 27625 245896 27659
rect 245844 27616 245896 27625
rect 268016 27684 268068 27736
rect 341248 27684 341300 27736
rect 337108 27659 337160 27668
rect 337108 27625 337117 27659
rect 337117 27625 337151 27659
rect 337151 27625 337160 27659
rect 337108 27616 337160 27625
rect 341156 27616 341208 27668
rect 421012 27616 421064 27668
rect 236276 27591 236328 27600
rect 236276 27557 236285 27591
rect 236285 27557 236319 27591
rect 236319 27557 236328 27591
rect 236276 27548 236328 27557
rect 265256 27591 265308 27600
rect 265256 27557 265265 27591
rect 265265 27557 265299 27591
rect 265299 27557 265308 27591
rect 265256 27548 265308 27557
rect 267924 27548 267976 27600
rect 284760 27548 284812 27600
rect 285956 27591 286008 27600
rect 285956 27557 285965 27591
rect 285965 27557 285999 27591
rect 285999 27557 286008 27591
rect 285956 27548 286008 27557
rect 299756 27548 299808 27600
rect 299940 27548 299992 27600
rect 301136 27548 301188 27600
rect 301228 27548 301280 27600
rect 306932 27548 306984 27600
rect 358728 27548 358780 27600
rect 306840 27480 306892 27532
rect 244372 26188 244424 26240
rect 245844 26231 245896 26240
rect 245844 26197 245853 26231
rect 245853 26197 245887 26231
rect 245887 26197 245896 26231
rect 245844 26188 245896 26197
rect 249984 26188 250036 26240
rect 250168 26188 250220 26240
rect 267924 26188 267976 26240
rect 299756 26231 299808 26240
rect 299756 26197 299765 26231
rect 299765 26197 299799 26231
rect 299799 26197 299808 26231
rect 299756 26188 299808 26197
rect 341156 26188 341208 26240
rect 421012 22720 421064 22772
rect 270500 22108 270552 22160
rect 270776 22108 270828 22160
rect 377036 22108 377088 22160
rect 424600 22108 424652 22160
rect 424508 22040 424560 22092
rect 377128 21972 377180 22024
rect 232412 19320 232464 19372
rect 302516 19320 302568 19372
rect 302608 19320 302660 19372
rect 336740 19320 336792 19372
rect 336924 19320 336976 19372
rect 367008 19363 367060 19372
rect 367008 19329 367017 19363
rect 367017 19329 367051 19363
rect 367051 19329 367060 19363
rect 367008 19320 367060 19329
rect 389456 19363 389508 19372
rect 389456 19329 389465 19363
rect 389465 19329 389499 19363
rect 389499 19329 389508 19363
rect 389456 19320 389508 19329
rect 265256 19295 265308 19304
rect 265256 19261 265265 19295
rect 265265 19261 265299 19295
rect 265299 19261 265308 19295
rect 265256 19252 265308 19261
rect 288808 19295 288860 19304
rect 288808 19261 288817 19295
rect 288817 19261 288851 19295
rect 288851 19261 288860 19295
rect 288808 19252 288860 19261
rect 325976 19252 326028 19304
rect 327264 19252 327316 19304
rect 366916 19295 366968 19304
rect 366916 19261 366925 19295
rect 366925 19261 366959 19295
rect 366959 19261 366968 19295
rect 366916 19252 366968 19261
rect 232504 19184 232556 19236
rect 325976 19116 326028 19168
rect 327264 19116 327316 19168
rect 362316 18028 362368 18080
rect 236276 18003 236328 18012
rect 236276 17969 236285 18003
rect 236285 17969 236319 18003
rect 236319 17969 236328 18003
rect 236276 17960 236328 17969
rect 270592 17960 270644 18012
rect 271972 17960 272024 18012
rect 284576 18003 284628 18012
rect 284576 17969 284585 18003
rect 284585 17969 284619 18003
rect 284619 17969 284628 18003
rect 284576 17960 284628 17969
rect 285956 18003 286008 18012
rect 285956 17969 285965 18003
rect 285965 17969 285999 18003
rect 285999 17969 286008 18003
rect 285956 17960 286008 17969
rect 294144 17960 294196 18012
rect 294236 17960 294288 18012
rect 265256 17892 265308 17944
rect 265440 17892 265492 17944
rect 273444 17935 273496 17944
rect 273444 17901 273453 17935
rect 273453 17901 273487 17935
rect 273487 17901 273496 17935
rect 273444 17892 273496 17901
rect 377128 17892 377180 17944
rect 270592 17824 270644 17876
rect 271972 17824 272024 17876
rect 271880 17756 271932 17808
rect 272340 17756 272392 17808
rect 395988 17144 396040 17196
rect 306380 17008 306432 17060
rect 315948 17008 316000 17060
rect 395988 16940 396040 16992
rect 347780 16872 347832 16924
rect 352656 16872 352708 16924
rect 385132 16804 385184 16856
rect 395896 16804 395948 16856
rect 417884 16804 417936 16856
rect 418252 16804 418304 16856
rect 456524 16804 456576 16856
rect 458824 16804 458876 16856
rect 289268 16736 289320 16788
rect 289912 16736 289964 16788
rect 437204 16736 437256 16788
rect 437480 16736 437532 16788
rect 310980 16668 311032 16720
rect 244188 16643 244240 16652
rect 244188 16609 244197 16643
rect 244197 16609 244231 16643
rect 244231 16609 244240 16643
rect 244188 16600 244240 16609
rect 246028 16600 246080 16652
rect 299756 16643 299808 16652
rect 299756 16609 299765 16643
rect 299765 16609 299799 16643
rect 299799 16609 299808 16643
rect 299756 16600 299808 16609
rect 310796 16600 310848 16652
rect 298100 16532 298152 16584
rect 298468 16532 298520 16584
rect 110328 15104 110380 15156
rect 274732 15104 274784 15156
rect 107476 15036 107528 15088
rect 273352 15036 273404 15088
rect 103428 14968 103480 15020
rect 271972 14968 272024 15020
rect 99288 14900 99340 14952
rect 270592 14900 270644 14952
rect 96528 14832 96580 14884
rect 269212 14832 269264 14884
rect 92388 14764 92440 14816
rect 266452 14764 266504 14816
rect 89628 14696 89680 14748
rect 265072 14696 265124 14748
rect 85488 14628 85540 14680
rect 263692 14628 263744 14680
rect 82728 14560 82780 14612
rect 262588 14560 262640 14612
rect 78588 14492 78640 14544
rect 260932 14492 260984 14544
rect 74448 14424 74500 14476
rect 259644 14424 259696 14476
rect 114468 14356 114520 14408
rect 276112 14356 276164 14408
rect 366824 14356 366876 14408
rect 367008 14356 367060 14408
rect 117228 14288 117280 14340
rect 277676 14288 277728 14340
rect 121368 14220 121420 14272
rect 278780 14220 278832 14272
rect 125416 14152 125468 14204
rect 280252 14152 280304 14204
rect 232136 14084 232188 14136
rect 232504 14084 232556 14136
rect 183468 13744 183520 13796
rect 303896 13744 303948 13796
rect 186228 13676 186280 13728
rect 306564 13676 306616 13728
rect 179328 13608 179380 13660
rect 302516 13608 302568 13660
rect 176568 13540 176620 13592
rect 301136 13540 301188 13592
rect 172428 13472 172480 13524
rect 299756 13472 299808 13524
rect 168288 13404 168340 13456
rect 298284 13404 298336 13456
rect 165528 13336 165580 13388
rect 296904 13336 296956 13388
rect 160008 13268 160060 13320
rect 294236 13268 294288 13320
rect 155868 13200 155920 13252
rect 292764 13200 292816 13252
rect 71688 13132 71740 13184
rect 258172 13132 258224 13184
rect 31668 13064 31720 13116
rect 241612 13064 241664 13116
rect 245844 13064 245896 13116
rect 246028 13064 246080 13116
rect 190368 12996 190420 13048
rect 307944 12996 307996 13048
rect 206928 12928 206980 12980
rect 314844 12928 314896 12980
rect 211068 12860 211120 12912
rect 316224 12860 316276 12912
rect 213828 12792 213880 12844
rect 317604 12792 317656 12844
rect 217968 12724 218020 12776
rect 318984 12724 319036 12776
rect 220728 12656 220780 12708
rect 320272 12656 320324 12708
rect 224868 12588 224920 12640
rect 321744 12588 321796 12640
rect 229008 12520 229060 12572
rect 323124 12520 323176 12572
rect 295616 12495 295668 12504
rect 295616 12461 295625 12495
rect 295625 12461 295659 12495
rect 295659 12461 295668 12495
rect 295616 12452 295668 12461
rect 173808 12384 173860 12436
rect 300952 12384 301004 12436
rect 392124 12384 392176 12436
rect 393044 12384 393096 12436
rect 426440 12384 426492 12436
rect 427544 12384 427596 12436
rect 169668 12316 169720 12368
rect 299572 12316 299624 12368
rect 166908 12248 166960 12300
rect 298192 12248 298244 12300
rect 162768 12180 162820 12232
rect 151728 12112 151780 12164
rect 291568 12112 291620 12164
rect 148968 12044 149020 12096
rect 290280 12044 290332 12096
rect 144828 11976 144880 12028
rect 288808 11976 288860 12028
rect 142068 11908 142120 11960
rect 287336 11908 287388 11960
rect 128268 11840 128320 11892
rect 281540 11840 281592 11892
rect 126888 11772 126940 11824
rect 281632 11772 281684 11824
rect 23388 11704 23440 11756
rect 238944 11704 238996 11756
rect 176476 11636 176528 11688
rect 302332 11636 302384 11688
rect 180708 11568 180760 11620
rect 303712 11568 303764 11620
rect 184848 11500 184900 11552
rect 305092 11500 305144 11552
rect 187608 11432 187660 11484
rect 306472 11432 306524 11484
rect 191748 11364 191800 11416
rect 308036 11364 308088 11416
rect 194508 11296 194560 11348
rect 309416 11296 309468 11348
rect 198648 11228 198700 11280
rect 307576 11228 307628 11280
rect 337108 11203 337160 11212
rect 337108 11169 337117 11203
rect 337117 11169 337151 11203
rect 337151 11169 337160 11203
rect 337108 11160 337160 11169
rect 113088 10956 113140 11008
rect 276020 10956 276072 11008
rect 108948 10888 109000 10940
rect 106188 10820 106240 10872
rect 271880 10820 271932 10872
rect 102048 10752 102100 10804
rect 270500 10752 270552 10804
rect 99196 10684 99248 10736
rect 269304 10684 269356 10736
rect 95148 10616 95200 10668
rect 91008 10548 91060 10600
rect 266728 10548 266780 10600
rect 64788 10480 64840 10532
rect 255596 10480 255648 10532
rect 60648 10412 60700 10464
rect 254032 10412 254084 10464
rect 56508 10344 56560 10396
rect 252652 10344 252704 10396
rect 53748 10276 53800 10328
rect 251272 10276 251324 10328
rect 117136 10208 117188 10260
rect 277584 10208 277636 10260
rect 119988 10140 120040 10192
rect 278964 10140 279016 10192
rect 124128 10072 124180 10124
rect 280344 10072 280396 10124
rect 366916 10115 366968 10124
rect 366916 10081 366925 10115
rect 366925 10081 366959 10115
rect 366959 10081 366968 10115
rect 366916 10072 366968 10081
rect 143448 10004 143500 10056
rect 288532 10004 288584 10056
rect 147588 9936 147640 9988
rect 289820 9936 289872 9988
rect 151636 9868 151688 9920
rect 291292 9868 291344 9920
rect 154488 9800 154540 9852
rect 292856 9800 292908 9852
rect 158628 9732 158680 9784
rect 294052 9732 294104 9784
rect 161388 9664 161440 9716
rect 295432 9664 295484 9716
rect 306656 9664 306708 9716
rect 306932 9664 306984 9716
rect 341248 9707 341300 9716
rect 341248 9673 341257 9707
rect 341257 9673 341291 9707
rect 341291 9673 341300 9707
rect 341248 9664 341300 9673
rect 358544 9707 358596 9716
rect 358544 9673 358553 9707
rect 358553 9673 358587 9707
rect 358587 9673 358596 9707
rect 358544 9664 358596 9673
rect 421472 9664 421524 9716
rect 203892 9596 203944 9648
rect 313372 9596 313424 9648
rect 330208 9639 330260 9648
rect 330208 9605 330217 9639
rect 330217 9605 330251 9639
rect 330251 9605 330260 9639
rect 330208 9596 330260 9605
rect 336924 9639 336976 9648
rect 336924 9605 336933 9639
rect 336933 9605 336967 9639
rect 336967 9605 336976 9639
rect 336924 9596 336976 9605
rect 389548 9596 389600 9648
rect 200396 9528 200448 9580
rect 311992 9528 312044 9580
rect 196808 9460 196860 9512
rect 310612 9460 310664 9512
rect 193220 9392 193272 9444
rect 309232 9392 309284 9444
rect 139676 9324 139728 9376
rect 287152 9324 287204 9376
rect 136088 9256 136140 9308
rect 285864 9256 285916 9308
rect 49332 9188 49384 9240
rect 249892 9188 249944 9240
rect 253848 9188 253900 9240
rect 334164 9188 334216 9240
rect 44548 9120 44600 9172
rect 247224 9120 247276 9172
rect 250352 9120 250404 9172
rect 332784 9120 332836 9172
rect 27896 9052 27948 9104
rect 233884 9052 233936 9104
rect 243176 9052 243228 9104
rect 330024 9052 330076 9104
rect 18328 8984 18380 9036
rect 236184 8984 236236 9036
rect 239588 8984 239640 9036
rect 328644 8984 328696 9036
rect 13636 8916 13688 8968
rect 234804 8916 234856 8968
rect 236000 8916 236052 8968
rect 325976 8916 326028 8968
rect 207480 8848 207532 8900
rect 314936 8848 314988 8900
rect 210976 8780 211028 8832
rect 316132 8780 316184 8832
rect 214656 8712 214708 8764
rect 317512 8712 317564 8764
rect 218152 8644 218204 8696
rect 318892 8644 318944 8696
rect 221740 8576 221792 8628
rect 320180 8576 320232 8628
rect 225328 8508 225380 8560
rect 321652 8508 321704 8560
rect 228916 8440 228968 8492
rect 323308 8440 323360 8492
rect 232504 8372 232556 8424
rect 324596 8372 324648 8424
rect 234896 8304 234948 8356
rect 235080 8304 235132 8356
rect 246764 8304 246816 8356
rect 331404 8304 331456 8356
rect 362224 8347 362276 8356
rect 362224 8313 362233 8347
rect 362233 8313 362267 8347
rect 362267 8313 362276 8347
rect 362224 8304 362276 8313
rect 376760 8347 376812 8356
rect 376760 8313 376769 8347
rect 376769 8313 376803 8347
rect 376803 8313 376812 8347
rect 376760 8304 376812 8313
rect 468760 8304 468812 8356
rect 469036 8304 469088 8356
rect 87328 8236 87380 8288
rect 265164 8236 265216 8288
rect 270500 8236 270552 8288
rect 340972 8236 341024 8288
rect 445484 8236 445536 8288
rect 523868 8236 523920 8288
rect 83832 8168 83884 8220
rect 263876 8168 263928 8220
rect 267004 8168 267056 8220
rect 339592 8168 339644 8220
rect 446956 8168 447008 8220
rect 527456 8168 527508 8220
rect 80244 8100 80296 8152
rect 262404 8100 262456 8152
rect 263416 8100 263468 8152
rect 338304 8100 338356 8152
rect 448244 8100 448296 8152
rect 531044 8100 531096 8152
rect 40960 8032 41012 8084
rect 245936 8032 245988 8084
rect 259828 8032 259880 8084
rect 451004 8032 451056 8084
rect 534540 8032 534592 8084
rect 37372 7964 37424 8016
rect 244188 7964 244240 8016
rect 256240 7964 256292 8016
rect 334072 7964 334124 8016
rect 452476 7964 452528 8016
rect 538128 7964 538180 8016
rect 33876 7896 33928 7948
rect 242992 7896 243044 7948
rect 252652 7896 252704 7948
rect 332692 7896 332744 7948
rect 453764 7896 453816 7948
rect 541716 7896 541768 7948
rect 30288 7828 30340 7880
rect 241796 7828 241848 7880
rect 249156 7828 249208 7880
rect 331312 7828 331364 7880
rect 455236 7828 455288 7880
rect 545304 7828 545356 7880
rect 26700 7760 26752 7812
rect 240416 7760 240468 7812
rect 245568 7760 245620 7812
rect 456616 7760 456668 7812
rect 548892 7760 548944 7812
rect 21916 7692 21968 7744
rect 238852 7692 238904 7744
rect 241980 7692 242032 7744
rect 328552 7692 328604 7744
rect 457996 7692 458048 7744
rect 552388 7692 552440 7744
rect 8852 7624 8904 7676
rect 4068 7556 4120 7608
rect 230664 7624 230716 7676
rect 234804 7624 234856 7676
rect 325792 7624 325844 7676
rect 459376 7624 459428 7676
rect 555976 7624 556028 7676
rect 227720 7556 227772 7608
rect 229008 7556 229060 7608
rect 231308 7556 231360 7608
rect 324412 7556 324464 7608
rect 460756 7556 460808 7608
rect 559564 7556 559616 7608
rect 134892 7488 134944 7540
rect 284576 7488 284628 7540
rect 444196 7488 444248 7540
rect 520280 7488 520332 7540
rect 138480 7420 138532 7472
rect 285956 7420 286008 7472
rect 442816 7420 442868 7472
rect 516784 7420 516836 7472
rect 141976 7352 142028 7404
rect 287060 7352 287112 7404
rect 441436 7352 441488 7404
rect 513196 7352 513248 7404
rect 145656 7284 145708 7336
rect 288440 7284 288492 7336
rect 440056 7284 440108 7336
rect 509608 7284 509660 7336
rect 149244 7216 149296 7268
rect 291200 7216 291252 7268
rect 152740 7148 152792 7200
rect 292580 7148 292632 7200
rect 156328 7080 156380 7132
rect 293960 7080 294012 7132
rect 159916 7012 159968 7064
rect 295340 7012 295392 7064
rect 233424 6944 233476 6996
rect 238392 6944 238444 6996
rect 327264 6944 327316 6996
rect 516692 6876 516744 6928
rect 516876 6876 516928 6928
rect 170588 6808 170640 6860
rect 299480 6808 299532 6860
rect 433248 6808 433300 6860
rect 491760 6808 491812 6860
rect 167092 6740 167144 6792
rect 298376 6740 298428 6792
rect 431776 6740 431828 6792
rect 490564 6740 490616 6792
rect 163504 6672 163556 6724
rect 296720 6672 296772 6724
rect 297364 6672 297416 6724
rect 336832 6672 336884 6724
rect 434628 6672 434680 6724
rect 495348 6672 495400 6724
rect 131396 6604 131448 6656
rect 283012 6604 283064 6656
rect 298100 6604 298152 6656
rect 338396 6604 338448 6656
rect 433156 6604 433208 6656
rect 494152 6604 494204 6656
rect 76656 6536 76708 6588
rect 261024 6536 261076 6588
rect 295892 6536 295944 6588
rect 335452 6536 335504 6588
rect 435916 6536 435968 6588
rect 497740 6536 497792 6588
rect 73068 6468 73120 6520
rect 259460 6468 259512 6520
rect 289820 6468 289872 6520
rect 339684 6468 339736 6520
rect 436008 6468 436060 6520
rect 498936 6468 498988 6520
rect 69480 6400 69532 6452
rect 258264 6400 258316 6452
rect 288440 6400 288492 6452
rect 341248 6400 341300 6452
rect 437296 6400 437348 6452
rect 501236 6400 501288 6452
rect 65984 6332 66036 6384
rect 256792 6332 256844 6384
rect 288532 6332 288584 6384
rect 343640 6332 343692 6384
rect 437388 6332 437440 6384
rect 502432 6332 502484 6384
rect 62396 6264 62448 6316
rect 255504 6264 255556 6316
rect 294328 6264 294380 6316
rect 350632 6264 350684 6316
rect 438768 6264 438820 6316
rect 504824 6264 504876 6316
rect 58808 6196 58860 6248
rect 253940 6196 253992 6248
rect 280068 6196 280120 6248
rect 345204 6196 345256 6248
rect 438676 6196 438728 6248
rect 506020 6196 506072 6248
rect 55220 6128 55272 6180
rect 251364 6128 251416 6180
rect 274088 6128 274140 6180
rect 342352 6128 342404 6180
rect 440148 6128 440200 6180
rect 508412 6128 508464 6180
rect 174176 6060 174228 6112
rect 300860 6060 300912 6112
rect 430396 6060 430448 6112
rect 486976 6060 487028 6112
rect 177764 5992 177816 6044
rect 302240 5992 302292 6044
rect 431868 5992 431920 6044
rect 488172 5992 488224 6044
rect 181352 5924 181404 5976
rect 303620 5924 303672 5976
rect 429108 5924 429160 5976
rect 483480 5924 483532 5976
rect 184848 5856 184900 5908
rect 305000 5856 305052 5908
rect 430488 5856 430540 5908
rect 484584 5856 484636 5908
rect 188436 5788 188488 5840
rect 306656 5788 306708 5840
rect 427728 5788 427780 5840
rect 479892 5788 479944 5840
rect 192024 5720 192076 5772
rect 307760 5720 307812 5772
rect 426348 5720 426400 5772
rect 476304 5720 476356 5772
rect 195612 5652 195664 5704
rect 309140 5652 309192 5704
rect 199200 5584 199252 5636
rect 310520 5584 310572 5636
rect 470600 5584 470652 5636
rect 202696 5516 202748 5568
rect 313280 5516 313332 5568
rect 468944 5516 468996 5568
rect 137284 5448 137336 5500
rect 285680 5448 285732 5500
rect 297824 5448 297876 5500
rect 352104 5448 352156 5500
rect 452568 5448 452620 5500
rect 540520 5448 540572 5500
rect 133788 5380 133840 5432
rect 284300 5380 284352 5432
rect 290740 5380 290792 5432
rect 349344 5380 349396 5432
rect 408408 5380 408460 5432
rect 433524 5380 433576 5432
rect 453856 5380 453908 5432
rect 544108 5380 544160 5432
rect 130200 5312 130252 5364
rect 283196 5312 283248 5364
rect 287152 5312 287204 5364
rect 347964 5312 348016 5364
rect 412364 5312 412416 5364
rect 440608 5312 440660 5364
rect 455328 5312 455380 5364
rect 547696 5312 547748 5364
rect 67180 5244 67232 5296
rect 256976 5244 257028 5296
rect 283656 5244 283708 5296
rect 346584 5244 346636 5296
rect 413836 5244 413888 5296
rect 444196 5244 444248 5296
rect 459468 5244 459520 5296
rect 48136 5176 48188 5228
rect 248512 5176 248564 5228
rect 251456 5176 251508 5228
rect 332600 5176 332652 5228
rect 415308 5176 415360 5228
rect 447784 5176 447836 5228
rect 460848 5176 460900 5228
rect 551192 5244 551244 5296
rect 17224 5108 17276 5160
rect 236092 5108 236144 5160
rect 247960 5108 248012 5160
rect 331220 5108 331272 5160
rect 416504 5108 416556 5160
rect 451280 5108 451332 5160
rect 12440 5040 12492 5092
rect 234712 5040 234764 5092
rect 244372 5040 244424 5092
rect 321652 5040 321704 5092
rect 327080 5040 327132 5092
rect 329840 5040 329892 5092
rect 337108 5040 337160 5092
rect 368572 5040 368624 5092
rect 381544 5040 381596 5092
rect 417976 5040 418028 5092
rect 454868 5040 454920 5092
rect 458088 5040 458140 5092
rect 7656 4972 7708 5024
rect 232136 4972 232188 5024
rect 240784 4972 240836 5024
rect 328736 4972 328788 5024
rect 333612 4972 333664 5024
rect 367192 4972 367244 5024
rect 419448 4972 419500 5024
rect 458456 4972 458508 5024
rect 2872 4904 2924 4956
rect 572 4836 624 4888
rect 229100 4904 229152 4956
rect 237196 4904 237248 4956
rect 321652 4904 321704 4956
rect 327080 4904 327132 4956
rect 361672 4904 361724 4956
rect 380164 4904 380216 4956
rect 420736 4904 420788 4956
rect 462044 4972 462096 5024
rect 463516 5108 463568 5160
rect 554780 5176 554832 5228
rect 464988 5040 465040 5092
rect 558368 5108 558420 5160
rect 465632 4972 465684 5024
rect 561956 5040 562008 5092
rect 466184 4904 466236 4956
rect 565544 4972 565596 5024
rect 230112 4836 230164 4888
rect 324320 4836 324372 4888
rect 326344 4836 326396 4888
rect 360292 4836 360344 4888
rect 422208 4836 422260 4888
rect 1676 4768 1728 4820
rect 230756 4768 230808 4820
rect 233700 4768 233752 4820
rect 325700 4768 325752 4820
rect 328460 4768 328512 4820
rect 363052 4768 363104 4820
rect 423588 4768 423640 4820
rect 469128 4836 469180 4888
rect 569040 4904 569092 4956
rect 572628 4836 572680 4888
rect 462136 4768 462188 4820
rect 579804 4768 579856 4820
rect 212264 4700 212316 4752
rect 316040 4700 316092 4752
rect 318708 4700 318760 4752
rect 215852 4632 215904 4684
rect 317420 4632 317472 4684
rect 323308 4700 323360 4752
rect 359188 4700 359240 4752
rect 451096 4700 451148 4752
rect 536932 4700 536984 4752
rect 333980 4632 334032 4684
rect 449808 4632 449860 4684
rect 533436 4632 533488 4684
rect 219348 4564 219400 4616
rect 318800 4564 318852 4616
rect 222936 4496 222988 4548
rect 321376 4564 321428 4616
rect 322756 4564 322808 4616
rect 448336 4564 448388 4616
rect 529848 4564 529900 4616
rect 320364 4496 320416 4548
rect 335360 4496 335412 4548
rect 447048 4496 447100 4548
rect 526260 4496 526312 4548
rect 226524 4428 226576 4480
rect 322940 4428 322992 4480
rect 325148 4428 325200 4480
rect 338120 4428 338172 4480
rect 445576 4428 445628 4480
rect 522672 4428 522724 4480
rect 201500 4360 201552 4412
rect 271144 4360 271196 4412
rect 301412 4360 301464 4412
rect 353484 4360 353536 4412
rect 444288 4360 444340 4412
rect 519084 4360 519136 4412
rect 205088 4292 205140 4344
rect 272524 4292 272576 4344
rect 305000 4292 305052 4344
rect 354956 4292 355008 4344
rect 442908 4292 442960 4344
rect 515588 4292 515640 4344
rect 230572 4224 230624 4276
rect 308588 4224 308640 4276
rect 356152 4224 356204 4276
rect 441528 4224 441580 4276
rect 512000 4224 512052 4276
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 140872 4156 140924 4208
rect 142068 4156 142120 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 160008 4156 160060 4208
rect 175372 4156 175424 4208
rect 176568 4156 176620 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 34980 4088 35032 4140
rect 50344 4088 50396 4140
rect 57612 4088 57664 4140
rect 250444 4088 250496 4140
rect 268108 4088 268160 4140
rect 269028 4088 269080 4140
rect 284760 4088 284812 4140
rect 285588 4088 285640 4140
rect 312176 4156 312228 4208
rect 357716 4156 357768 4208
rect 424968 4156 425020 4208
rect 472716 4156 472768 4208
rect 20720 4020 20772 4072
rect 28264 4020 28316 4072
rect 50528 4020 50580 4072
rect 249064 4020 249116 4072
rect 295892 4088 295944 4140
rect 296720 4088 296772 4140
rect 297916 4088 297968 4140
rect 300308 4088 300360 4140
rect 332416 4088 332468 4140
rect 333244 4088 333296 4140
rect 334716 4088 334768 4140
rect 335268 4088 335320 4140
rect 338764 4088 338816 4140
rect 339500 4088 339552 4140
rect 340788 4088 340840 4140
rect 345664 4088 345716 4140
rect 347872 4088 347924 4140
rect 349068 4088 349120 4140
rect 351184 4088 351236 4140
rect 351368 4088 351420 4140
rect 351828 4088 351880 4140
rect 354956 4088 355008 4140
rect 355968 4088 356020 4140
rect 358084 4088 358136 4140
rect 362132 4088 362184 4140
rect 362868 4088 362920 4140
rect 363328 4088 363380 4140
rect 364248 4088 364300 4140
rect 365720 4088 365772 4140
rect 366916 4088 366968 4140
rect 369216 4088 369268 4140
rect 369768 4088 369820 4140
rect 370412 4088 370464 4140
rect 371148 4088 371200 4140
rect 377588 4088 377640 4140
rect 378048 4088 378100 4140
rect 378784 4088 378836 4140
rect 385316 4088 385368 4140
rect 390560 4088 390612 4140
rect 391848 4088 391900 4140
rect 393136 4088 393188 4140
rect 395436 4088 395488 4140
rect 398104 4088 398156 4140
rect 403716 4088 403768 4140
rect 438216 4088 438268 4140
rect 442264 4088 442316 4140
rect 445668 4088 445720 4140
rect 521476 4088 521528 4140
rect 529204 4088 529256 4140
rect 575020 4088 575072 4140
rect 298100 4020 298152 4072
rect 302608 4020 302660 4072
rect 309784 4020 309836 4072
rect 313372 4020 313424 4072
rect 46940 3952 46992 4004
rect 248696 3952 248748 4004
rect 257436 3952 257488 4004
rect 297364 3952 297416 4004
rect 314568 3952 314620 4004
rect 374000 4020 374052 4072
rect 376760 4020 376812 4072
rect 383568 4020 383620 4072
rect 384304 4020 384356 4072
rect 393228 4020 393280 4072
rect 396632 4020 396684 4072
rect 411168 4020 411220 4072
rect 439412 4020 439464 4072
rect 439596 4020 439648 4072
rect 448428 4020 448480 4072
rect 528652 4020 528704 4072
rect 530584 4020 530636 4072
rect 582196 4020 582248 4072
rect 358820 3952 358872 4004
rect 359740 3952 359792 4004
rect 402888 3952 402940 4004
rect 419172 3952 419224 4004
rect 420276 3952 420328 4004
rect 423956 3952 424008 4004
rect 424600 3952 424652 4004
rect 425152 3952 425204 4004
rect 450176 3952 450228 4004
rect 451188 3952 451240 4004
rect 535736 3952 535788 4004
rect 45744 3884 45796 3936
rect 247684 3884 247736 3936
rect 282460 3884 282512 3936
rect 39764 3816 39816 3868
rect 245752 3816 245804 3868
rect 264612 3816 264664 3868
rect 19524 3748 19576 3800
rect 32404 3748 32456 3800
rect 38568 3748 38620 3800
rect 245660 3748 245712 3800
rect 278872 3748 278924 3800
rect 289544 3816 289596 3868
rect 365812 3884 365864 3936
rect 371608 3884 371660 3936
rect 412456 3884 412508 3936
rect 441620 3884 441672 3936
rect 453672 3884 453724 3936
rect 453948 3884 454000 3936
rect 542912 3884 542964 3936
rect 285956 3748 286008 3800
rect 335820 3748 335872 3800
rect 342904 3816 342956 3868
rect 343088 3816 343140 3868
rect 369124 3816 369176 3868
rect 372804 3816 372856 3868
rect 373908 3816 373960 3868
rect 413928 3816 413980 3868
rect 445392 3816 445444 3868
rect 550088 3816 550140 3868
rect 341524 3748 341576 3800
rect 341892 3748 341944 3800
rect 370136 3748 370188 3800
rect 374000 3748 374052 3800
rect 375288 3748 375340 3800
rect 399484 3748 399536 3800
rect 408500 3748 408552 3800
rect 411076 3748 411128 3800
rect 32680 3680 32732 3732
rect 243084 3680 243136 3732
rect 326436 3680 326488 3732
rect 328460 3680 328512 3732
rect 331220 3680 331272 3732
rect 338304 3680 338356 3732
rect 368664 3680 368716 3732
rect 375196 3680 375248 3732
rect 383844 3680 383896 3732
rect 400128 3680 400180 3732
rect 412088 3680 412140 3732
rect 412548 3680 412600 3732
rect 443000 3748 443052 3800
rect 24308 3612 24360 3664
rect 239036 3612 239088 3664
rect 262220 3612 262272 3664
rect 11244 3544 11296 3596
rect 19984 3544 20036 3596
rect 25504 3544 25556 3596
rect 240324 3544 240376 3596
rect 265808 3544 265860 3596
rect 325148 3612 325200 3664
rect 325240 3612 325292 3664
rect 322848 3544 322900 3596
rect 327080 3544 327132 3596
rect 358912 3612 358964 3664
rect 360936 3612 360988 3664
rect 377404 3612 377456 3664
rect 400036 3612 400088 3664
rect 413192 3612 413244 3664
rect 416688 3612 416740 3664
rect 421564 3612 421616 3664
rect 427084 3612 427136 3664
rect 431132 3612 431184 3664
rect 442356 3612 442408 3664
rect 443644 3612 443696 3664
rect 446588 3612 446640 3664
rect 452476 3748 452528 3800
rect 456708 3748 456760 3800
rect 460112 3748 460164 3800
rect 460296 3748 460348 3800
rect 463240 3748 463292 3800
rect 449164 3612 449216 3664
rect 16028 3476 16080 3528
rect 236276 3476 236328 3528
rect 258632 3476 258684 3528
rect 320364 3476 320416 3528
rect 320456 3476 320508 3528
rect 321192 3476 321244 3528
rect 321652 3476 321704 3528
rect 361856 3544 361908 3596
rect 402244 3544 402296 3596
rect 415676 3544 415728 3596
rect 418068 3544 418120 3596
rect 457260 3544 457312 3596
rect 460204 3680 460256 3732
rect 557172 3748 557224 3800
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 14832 3408 14884 3460
rect 234988 3408 235040 3460
rect 255044 3408 255096 3460
rect 318708 3408 318760 3460
rect 322756 3408 322808 3460
rect 324044 3408 324096 3460
rect 363144 3476 363196 3528
rect 363604 3408 363656 3460
rect 368020 3408 368072 3460
rect 379980 3476 380032 3528
rect 380808 3476 380860 3528
rect 381176 3476 381228 3528
rect 382188 3476 382240 3528
rect 388260 3476 388312 3528
rect 389088 3476 389140 3528
rect 395988 3476 396040 3528
rect 401324 3476 401376 3528
rect 402796 3476 402848 3528
rect 413284 3476 413336 3528
rect 414480 3476 414532 3528
rect 420828 3476 420880 3528
rect 460848 3476 460900 3528
rect 462228 3544 462280 3596
rect 564348 3680 564400 3732
rect 463608 3612 463660 3664
rect 566740 3612 566792 3664
rect 463516 3544 463568 3596
rect 466368 3544 466420 3596
rect 571432 3544 571484 3596
rect 466276 3476 466328 3528
rect 573824 3476 573876 3528
rect 379704 3408 379756 3460
rect 382372 3408 382424 3460
rect 386604 3408 386656 3460
rect 395896 3408 395948 3460
rect 402520 3408 402572 3460
rect 403624 3408 403676 3460
rect 407304 3408 407356 3460
rect 29092 3340 29144 3392
rect 35164 3340 35216 3392
rect 36176 3340 36228 3392
rect 39304 3340 39356 3392
rect 10048 3272 10100 3324
rect 13084 3272 13136 3324
rect 42156 3272 42208 3324
rect 57244 3272 57296 3324
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 61384 3272 61436 3324
rect 52828 3204 52880 3256
rect 53748 3204 53800 3256
rect 54024 3204 54076 3256
rect 43352 3136 43404 3188
rect 64788 3204 64840 3256
rect 251824 3340 251876 3392
rect 289820 3340 289872 3392
rect 299112 3340 299164 3392
rect 302884 3340 302936 3392
rect 310980 3340 311032 3392
rect 341524 3340 341576 3392
rect 71872 3272 71924 3324
rect 253204 3272 253256 3324
rect 61200 3136 61252 3188
rect 66904 3068 66956 3120
rect 68284 3136 68336 3188
rect 71044 3068 71096 3120
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 75460 3136 75512 3188
rect 79324 3136 79376 3188
rect 82636 3136 82688 3188
rect 84844 3204 84896 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 88524 3204 88576 3256
rect 89628 3204 89680 3256
rect 254584 3204 254636 3256
rect 269304 3204 269356 3256
rect 89720 3068 89772 3120
rect 255964 3136 256016 3188
rect 272892 3136 272944 3188
rect 288440 3272 288492 3324
rect 303804 3272 303856 3324
rect 344284 3272 344336 3324
rect 353760 3340 353812 3392
rect 375656 3340 375708 3392
rect 404268 3340 404320 3392
rect 422760 3408 422812 3460
rect 424324 3408 424376 3460
rect 467932 3408 467984 3460
rect 469036 3408 469088 3460
rect 578608 3408 578660 3460
rect 409788 3340 409840 3392
rect 433984 3340 434036 3392
rect 435824 3340 435876 3392
rect 438124 3340 438176 3392
rect 348424 3272 348476 3324
rect 349068 3272 349120 3324
rect 365536 3272 365588 3324
rect 394516 3272 394568 3324
rect 399024 3272 399076 3324
rect 405004 3272 405056 3324
rect 416872 3272 416924 3324
rect 420184 3272 420236 3324
rect 446588 3272 446640 3324
rect 503628 3272 503680 3324
rect 514024 3340 514076 3392
rect 517888 3340 517940 3392
rect 514392 3272 514444 3324
rect 516876 3272 516928 3324
rect 525064 3340 525116 3392
rect 527824 3340 527876 3392
rect 567844 3340 567896 3392
rect 276480 3204 276532 3256
rect 288532 3204 288584 3256
rect 291936 3204 291988 3256
rect 316684 3204 316736 3256
rect 318064 3204 318116 3256
rect 345756 3204 345808 3256
rect 350264 3204 350316 3256
rect 355324 3204 355376 3256
rect 357348 3204 357400 3256
rect 376024 3204 376076 3256
rect 394608 3204 394660 3256
rect 400220 3204 400272 3256
rect 409144 3204 409196 3256
rect 432328 3204 432380 3256
rect 437020 3204 437072 3256
rect 446220 3204 446272 3256
rect 496544 3204 496596 3256
rect 512644 3204 512696 3256
rect 577412 3272 577464 3324
rect 570236 3204 570288 3256
rect 277676 3136 277728 3188
rect 290464 3136 290516 3188
rect 309784 3136 309836 3188
rect 336004 3136 336056 3188
rect 340696 3136 340748 3188
rect 346676 3136 346728 3188
rect 370504 3136 370556 3188
rect 407028 3136 407080 3188
rect 429936 3136 429988 3188
rect 431224 3136 431276 3188
rect 94504 3068 94556 3120
rect 95148 3068 95200 3120
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 98092 3068 98144 3120
rect 99196 3068 99248 3120
rect 101588 3068 101640 3120
rect 102048 3068 102100 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 105176 3068 105228 3120
rect 106188 3068 106240 3120
rect 106372 3068 106424 3120
rect 107476 3068 107528 3120
rect 77944 3000 77996 3052
rect 93308 3000 93360 3052
rect 102600 3000 102652 3052
rect 79048 2932 79100 2984
rect 86132 2932 86184 2984
rect 96896 2932 96948 2984
rect 257344 3068 257396 3120
rect 295524 3068 295576 3120
rect 319444 3068 319496 3120
rect 327724 3068 327776 3120
rect 328828 3068 328880 3120
rect 359464 3068 359516 3120
rect 372988 3068 373040 3120
rect 405648 3068 405700 3120
rect 426348 3068 426400 3120
rect 428464 3068 428516 3120
rect 475108 3068 475160 3120
rect 475384 3068 475436 3120
rect 477500 3068 477552 3120
rect 505744 3136 505796 3188
rect 563152 3136 563204 3188
rect 482284 3068 482336 3120
rect 524972 3068 525024 3120
rect 560760 3068 560812 3120
rect 103980 2864 104032 2916
rect 258724 3000 258776 3052
rect 293132 3000 293184 3052
rect 312544 3000 312596 3052
rect 315764 3000 315816 3052
rect 323308 3000 323360 3052
rect 327632 3000 327684 3052
rect 336188 3000 336240 3052
rect 112352 2932 112404 2984
rect 113088 2932 113140 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 115940 2932 115992 2984
rect 116952 2932 117004 2984
rect 119436 2932 119488 2984
rect 119988 2932 120040 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 111156 2864 111208 2916
rect 258816 2932 258868 2984
rect 316960 2932 317012 2984
rect 336004 2932 336056 2984
rect 352472 2932 352524 2984
rect 352564 2932 352616 2984
rect 364524 3000 364576 3052
rect 365536 3000 365588 3052
rect 376392 3000 376444 3052
rect 381636 3000 381688 3052
rect 406384 3000 406436 3052
rect 410892 3000 410944 3052
rect 420368 3000 420420 3052
rect 431316 3000 431368 3052
rect 459652 3000 459704 3052
rect 489368 3000 489420 3052
rect 509884 3000 509936 3052
rect 523684 3000 523736 3052
rect 553584 3000 553636 3052
rect 95884 2796 95936 2848
rect 114744 2796 114796 2848
rect 260104 2864 260156 2916
rect 275284 2864 275336 2916
rect 275928 2864 275980 2916
rect 319260 2864 319312 2916
rect 326344 2864 326396 2916
rect 335912 2864 335964 2916
rect 336188 2864 336240 2916
rect 340972 2864 341024 2916
rect 344284 2864 344336 2916
rect 121828 2796 121880 2848
rect 261484 2796 261536 2848
rect 330024 2796 330076 2848
rect 344376 2796 344428 2848
rect 356704 2864 356756 2916
rect 374092 2932 374144 2984
rect 398196 2932 398248 2984
rect 404912 2932 404964 2984
rect 417424 2932 417476 2984
rect 428740 2932 428792 2984
rect 429844 2932 429896 2984
rect 448980 2932 449032 2984
rect 367284 2864 367336 2916
rect 385868 2864 385920 2916
rect 387064 2864 387116 2916
rect 416596 2864 416648 2916
rect 356152 2796 356204 2848
rect 356796 2796 356848 2848
rect 357072 2796 357124 2848
rect 375840 2796 375892 2848
rect 388444 2796 388496 2848
rect 439504 2796 439556 2848
rect 481088 2932 481140 2984
rect 521016 2932 521068 2984
rect 546500 2932 546552 2984
rect 473912 2864 473964 2916
rect 520924 2864 520976 2916
rect 539324 2864 539376 2916
rect 466828 2796 466880 2848
rect 518164 2796 518216 2848
rect 532240 2796 532292 2848
rect 362224 2728 362276 2780
rect 387064 2728 387116 2780
rect 261024 1096 261076 1148
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 164700 552 164752 604
rect 165528 552 165580 604
rect 165896 552 165948 604
rect 166908 552 166960 604
rect 169392 552 169444 604
rect 169668 552 169720 604
rect 182548 552 182600 604
rect 183468 552 183520 604
rect 183744 552 183796 604
rect 184756 552 184808 604
rect 187240 552 187292 604
rect 187608 552 187660 604
rect 189632 552 189684 604
rect 190368 552 190420 604
rect 281264 552 281316 604
rect 281448 552 281500 604
rect 389456 595 389508 604
rect 389456 561 389465 595
rect 389465 561 389499 595
rect 389499 561 389508 595
rect 389456 552 389508 561
rect 393596 552 393648 604
rect 394240 552 394292 604
rect 397460 552 397512 604
rect 397828 552 397880 604
rect 405924 552 405976 604
rect 406108 552 406160 604
rect 463700 552 463752 604
rect 464436 552 464488 604
rect 469220 552 469272 604
rect 470324 552 470376 604
rect 471520 595 471572 604
rect 471520 561 471529 595
rect 471529 561 471563 595
rect 471563 561 471572 595
rect 471520 552 471572 561
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700670 137876 703520
rect 154132 700738 154160 703520
rect 170324 700942 170352 703520
rect 202800 701010 202828 703520
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 170312 700936 170364 700942
rect 170312 700878 170364 700884
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 218992 700262 219020 703520
rect 218980 700256 219032 700262
rect 218980 700198 219032 700204
rect 235184 700058 235212 703520
rect 235172 700052 235224 700058
rect 235172 699994 235224 700000
rect 267660 699990 267688 703520
rect 267648 699984 267700 699990
rect 267648 699926 267700 699932
rect 283852 699922 283880 703520
rect 283840 699916 283892 699922
rect 283840 699858 283892 699864
rect 300136 699718 300164 703520
rect 328368 700868 328420 700874
rect 328368 700810 328420 700816
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 300780 584662 300808 699654
rect 321468 696992 321520 696998
rect 321468 696934 321520 696940
rect 320088 673532 320140 673538
rect 320088 673474 320140 673480
rect 315948 650072 316000 650078
rect 315948 650014 316000 650020
rect 313188 626612 313240 626618
rect 313188 626554 313240 626560
rect 309048 603152 309100 603158
rect 309048 603094 309100 603100
rect 300768 584656 300820 584662
rect 300768 584598 300820 584604
rect 304540 583704 304592 583710
rect 304540 583646 304592 583652
rect 298192 583636 298244 583642
rect 298192 583578 298244 583584
rect 256056 583568 256108 583574
rect 4802 583536 4858 583545
rect 256056 583510 256108 583516
rect 4802 583471 4858 583480
rect 251824 583500 251876 583506
rect 4712 583364 4764 583370
rect 4712 583306 4764 583312
rect 3148 583092 3200 583098
rect 3148 583034 3200 583040
rect 3056 567384 3108 567390
rect 3054 567352 3056 567361
rect 3108 567352 3110 567361
rect 3054 567287 3110 567296
rect 2780 553104 2832 553110
rect 2778 553072 2780 553081
rect 2832 553072 2834 553081
rect 2778 553007 2834 553016
rect 3056 538688 3108 538694
rect 3054 538656 3056 538665
rect 3108 538656 3110 538665
rect 3054 538591 3110 538600
rect 3056 510264 3108 510270
rect 3056 510206 3108 510212
rect 3068 509969 3096 510206
rect 3054 509960 3110 509969
rect 3054 509895 3110 509904
rect 2780 496732 2832 496738
rect 2780 496674 2832 496680
rect 2792 495553 2820 496674
rect 2778 495544 2834 495553
rect 2778 495479 2834 495488
rect 2964 481160 3016 481166
rect 2962 481128 2964 481137
rect 3016 481128 3018 481137
rect 2962 481063 3018 481072
rect 3160 452441 3188 583034
rect 3240 582888 3292 582894
rect 3240 582830 3292 582836
rect 3146 452432 3202 452441
rect 3146 452367 3202 452376
rect 3148 438864 3200 438870
rect 3148 438806 3200 438812
rect 3160 438025 3188 438806
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 3148 424108 3200 424114
rect 3148 424050 3200 424056
rect 3160 423745 3188 424050
rect 3146 423736 3202 423745
rect 3146 423671 3202 423680
rect 3252 395049 3280 582830
rect 4068 582684 4120 582690
rect 4068 582626 4120 582632
rect 3884 582548 3936 582554
rect 3884 582490 3936 582496
rect 3700 582412 3752 582418
rect 3700 582354 3752 582360
rect 3332 578536 3384 578542
rect 3332 578478 3384 578484
rect 3238 395040 3294 395049
rect 3238 394975 3294 394984
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 3344 366217 3372 578478
rect 3608 578400 3660 578406
rect 3608 578342 3660 578348
rect 3424 578332 3476 578338
rect 3424 578274 3476 578280
rect 3330 366208 3386 366217
rect 3330 366143 3386 366152
rect 3332 324284 3384 324290
rect 3332 324226 3384 324232
rect 3344 323105 3372 324226
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 2780 308848 2832 308854
rect 2778 308816 2780 308825
rect 2832 308816 2834 308825
rect 2778 308751 2834 308760
rect 2962 295216 3018 295225
rect 2962 295151 3018 295160
rect 2976 294409 3004 295151
rect 2962 294400 3018 294409
rect 2962 294335 3018 294344
rect 2780 252544 2832 252550
rect 2780 252486 2832 252492
rect 2792 251297 2820 252486
rect 2778 251288 2834 251297
rect 2778 251223 2834 251232
rect 3056 237380 3108 237386
rect 3056 237322 3108 237328
rect 3068 237017 3096 237322
rect 3054 237008 3110 237017
rect 3054 236943 3110 236952
rect 2780 165504 2832 165510
rect 2780 165446 2832 165452
rect 2792 165073 2820 165446
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 3332 151768 3384 151774
rect 3332 151710 3384 151716
rect 3344 150793 3372 151710
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2780 136536 2832 136542
rect 2780 136478 2832 136484
rect 2792 136377 2820 136478
rect 2778 136368 2834 136377
rect 2778 136303 2834 136312
rect 2780 122324 2832 122330
rect 2780 122266 2832 122272
rect 2792 122097 2820 122266
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3436 93265 3464 578274
rect 3516 578264 3568 578270
rect 3516 578206 3568 578212
rect 3528 107681 3556 578206
rect 3620 179489 3648 578342
rect 3712 193905 3740 582354
rect 3792 579896 3844 579902
rect 3792 579838 3844 579844
rect 3804 208185 3832 579838
rect 3896 222601 3924 582490
rect 3976 578468 4028 578474
rect 3976 578410 4028 578416
rect 3988 265713 4016 578410
rect 4080 280129 4108 582626
rect 4724 553110 4752 583306
rect 4712 553104 4764 553110
rect 4712 553046 4764 553052
rect 4066 280120 4122 280129
rect 4066 280055 4122 280064
rect 3974 265704 4030 265713
rect 3974 265639 4030 265648
rect 3882 222592 3938 222601
rect 3882 222527 3938 222536
rect 3790 208176 3846 208185
rect 3790 208111 3846 208120
rect 3698 193896 3754 193905
rect 3698 193831 3754 193840
rect 3606 179480 3662 179489
rect 3606 179415 3662 179424
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 2780 79824 2832 79830
rect 2780 79766 2832 79772
rect 2792 78985 2820 79766
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 4816 50522 4844 583471
rect 251824 583442 251876 583448
rect 245568 583432 245620 583438
rect 245568 583374 245620 583380
rect 5448 583296 5500 583302
rect 5448 583238 5500 583244
rect 5356 582820 5408 582826
rect 5356 582762 5408 582768
rect 5264 582616 5316 582622
rect 5078 582584 5134 582593
rect 5264 582558 5316 582564
rect 5078 582519 5134 582528
rect 4988 579828 5040 579834
rect 4988 579770 5040 579776
rect 4896 579760 4948 579766
rect 4896 579702 4948 579708
rect 4908 79830 4936 579702
rect 5000 122330 5028 579770
rect 5092 136542 5120 582519
rect 5172 582480 5224 582486
rect 5172 582422 5224 582428
rect 5184 165510 5212 582422
rect 5276 252550 5304 582558
rect 5368 308854 5396 582762
rect 5460 496738 5488 583238
rect 10324 583228 10376 583234
rect 10324 583170 10376 583176
rect 6276 583160 6328 583166
rect 6276 583102 6328 583108
rect 6184 579692 6236 579698
rect 6184 579634 6236 579640
rect 5448 496732 5500 496738
rect 5448 496674 5500 496680
rect 5356 308848 5408 308854
rect 5356 308790 5408 308796
rect 5264 252544 5316 252550
rect 5264 252486 5316 252492
rect 5172 165504 5224 165510
rect 5172 165446 5224 165452
rect 5080 136536 5132 136542
rect 5080 136478 5132 136484
rect 4988 122324 5040 122330
rect 4988 122266 5040 122272
rect 4896 79824 4948 79830
rect 4896 79766 4948 79772
rect 2780 50516 2832 50522
rect 2780 50458 2832 50464
rect 4804 50516 4856 50522
rect 4804 50458 4856 50464
rect 2792 50153 2820 50458
rect 2778 50144 2834 50153
rect 2778 50079 2834 50088
rect 6196 35902 6224 579634
rect 6288 424114 6316 583102
rect 6644 580168 6696 580174
rect 6644 580110 6696 580116
rect 6552 580100 6604 580106
rect 6552 580042 6604 580048
rect 6460 580032 6512 580038
rect 6460 579974 6512 579980
rect 6368 579964 6420 579970
rect 6368 579906 6420 579912
rect 6380 481166 6408 579906
rect 6472 510270 6500 579974
rect 6564 538694 6592 580042
rect 6656 567390 6684 580110
rect 6644 567384 6696 567390
rect 6644 567326 6696 567332
rect 6552 538688 6604 538694
rect 6552 538630 6604 538636
rect 6460 510264 6512 510270
rect 6460 510206 6512 510212
rect 6368 481160 6420 481166
rect 6368 481102 6420 481108
rect 10336 438870 10364 583170
rect 13084 583024 13136 583030
rect 13084 582966 13136 582972
rect 10324 438864 10376 438870
rect 10324 438806 10376 438812
rect 6276 424108 6328 424114
rect 6276 424050 6328 424056
rect 13096 380866 13124 582966
rect 14464 582956 14516 582962
rect 14464 582898 14516 582904
rect 13084 380860 13136 380866
rect 13084 380802 13136 380808
rect 13084 337408 13136 337414
rect 10322 337376 10378 337385
rect 13084 337350 13136 337356
rect 10322 337311 10378 337320
rect 3148 35896 3200 35902
rect 3146 35864 3148 35873
rect 6184 35896 6236 35902
rect 3200 35864 3202 35873
rect 6184 35838 6236 35844
rect 3146 35799 3202 35808
rect 3146 11656 3202 11665
rect 3146 11591 3202 11600
rect 3160 7177 3188 11591
rect 8852 7676 8904 7682
rect 8852 7618 8904 7624
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 3146 7168 3202 7177
rect 3146 7103 3202 7112
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8864 480 8892 7618
rect 10336 3466 10364 337311
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10048 3324 10100 3330
rect 10048 3266 10100 3272
rect 10060 480 10088 3266
rect 11256 480 11284 3538
rect 12452 480 12480 5034
rect 13096 3330 13124 337350
rect 14476 324290 14504 582898
rect 17222 582856 17278 582865
rect 17222 582791 17278 582800
rect 15844 582752 15896 582758
rect 15844 582694 15896 582700
rect 14464 324284 14516 324290
rect 14464 324226 14516 324232
rect 15856 237386 15884 582694
rect 15844 237380 15896 237386
rect 15844 237322 15896 237328
rect 17236 151774 17264 582791
rect 24122 582720 24178 582729
rect 24122 582655 24178 582664
rect 19984 337476 20036 337482
rect 19984 337418 20036 337424
rect 17224 151768 17276 151774
rect 17224 151710 17276 151716
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13084 3324 13136 3330
rect 13084 3266 13136 3272
rect 13648 480 13676 8910
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 480 14872 3402
rect 16040 480 16068 3470
rect 17236 480 17264 5102
rect 18340 480 18368 8978
rect 19524 3800 19576 3806
rect 19524 3742 19576 3748
rect 19536 480 19564 3742
rect 19996 3602 20024 337418
rect 24136 64870 24164 582655
rect 245580 579972 245608 583374
rect 251836 579972 251864 583442
rect 256068 579972 256096 583510
rect 293958 583264 294014 583273
rect 293958 583199 294014 583208
rect 289728 581392 289780 581398
rect 289728 581334 289780 581340
rect 287612 581324 287664 581330
rect 287612 581266 287664 581272
rect 283472 581256 283524 581262
rect 283472 581198 283524 581204
rect 281356 581188 281408 581194
rect 281356 581130 281408 581136
rect 275008 581120 275060 581126
rect 275008 581062 275060 581068
rect 264520 581052 264572 581058
rect 264520 580994 264572 581000
rect 262404 580304 262456 580310
rect 262404 580246 262456 580252
rect 262416 579972 262444 580246
rect 264532 579972 264560 580994
rect 268660 580372 268712 580378
rect 268660 580314 268712 580320
rect 268672 579972 268700 580314
rect 275020 579972 275048 581062
rect 281368 579972 281396 581130
rect 283484 579972 283512 581198
rect 287624 579972 287652 581266
rect 289740 579972 289768 581334
rect 293972 579972 294000 583199
rect 296076 581460 296128 581466
rect 296076 581402 296128 581408
rect 296088 579972 296116 581402
rect 298204 579972 298232 583578
rect 300306 583400 300362 583409
rect 300306 583335 300362 583344
rect 300320 579972 300348 583335
rect 302424 581528 302476 581534
rect 302424 581470 302476 581476
rect 302436 579972 302464 581470
rect 304552 579972 304580 583646
rect 306564 580236 306616 580242
rect 306564 580178 306616 580184
rect 306576 579972 306604 580178
rect 309060 579986 309088 603094
rect 311808 592068 311860 592074
rect 311808 592010 311860 592016
rect 311820 580122 311848 592010
rect 308706 579958 309088 579986
rect 311268 580094 311848 580122
rect 311268 579850 311296 580094
rect 313200 579986 313228 626554
rect 312938 579958 313228 579986
rect 315960 579850 315988 650014
rect 317328 638988 317380 638994
rect 317328 638930 317380 638936
rect 317340 579986 317368 638930
rect 320100 580122 320128 673474
rect 317170 579958 317368 579986
rect 319732 580094 320128 580122
rect 319732 579850 319760 580094
rect 321480 579986 321508 696934
rect 324228 685908 324280 685914
rect 324228 685850 324280 685856
rect 321402 579958 321508 579986
rect 324240 579850 324268 685850
rect 325516 584452 325568 584458
rect 325516 584394 325568 584400
rect 325528 579972 325556 584394
rect 328380 579850 328408 700810
rect 329748 700800 329800 700806
rect 329748 700742 329800 700748
rect 329760 579972 329788 700742
rect 332520 699718 332548 703520
rect 336648 700188 336700 700194
rect 336648 700130 336700 700136
rect 335268 700120 335320 700126
rect 335268 700062 335320 700068
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 331864 584520 331916 584526
rect 331864 584462 331916 584468
rect 331876 579972 331904 584462
rect 335280 580122 335308 700062
rect 334452 580094 335308 580122
rect 334452 579850 334480 580094
rect 336660 579850 336688 700130
rect 343548 699848 343600 699854
rect 343548 699790 343600 699796
rect 340788 699780 340840 699786
rect 340788 699722 340840 699728
rect 338212 584588 338264 584594
rect 338212 584530 338264 584536
rect 338224 579972 338252 584530
rect 340800 579986 340828 699722
rect 340354 579958 340828 579986
rect 343560 579850 343588 699790
rect 348804 699718 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365208 703474
rect 358820 701004 358872 701010
rect 358820 700946 358872 700952
rect 356060 700052 356112 700058
rect 356060 699994 356112 700000
rect 351920 699984 351972 699990
rect 351920 699926 351972 699932
rect 346400 699712 346452 699718
rect 346400 699654 346452 699660
rect 347780 699712 347832 699718
rect 347780 699654 347832 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 344468 584724 344520 584730
rect 344468 584666 344520 584672
rect 344480 579972 344508 584666
rect 346412 579986 346440 699654
rect 346412 579958 346610 579986
rect 310822 579822 311296 579850
rect 315054 579822 315988 579850
rect 319286 579822 319760 579850
rect 323426 579822 324268 579850
rect 327658 579822 328408 579850
rect 334006 579822 334480 579850
rect 336122 579822 336688 579850
rect 342378 579822 343588 579850
rect 347792 579850 347820 699654
rect 350816 584656 350868 584662
rect 350816 584598 350868 584604
rect 350828 579972 350856 584598
rect 351932 579850 351960 699926
rect 354680 699916 354732 699922
rect 354680 699858 354732 699864
rect 354692 579986 354720 699858
rect 354692 579958 355074 579986
rect 356072 579850 356100 699994
rect 358832 579850 358860 700946
rect 362960 700936 363012 700942
rect 362960 700878 363012 700884
rect 360200 700256 360252 700262
rect 360200 700198 360252 700204
rect 360212 580122 360240 700198
rect 360212 580094 360884 580122
rect 360856 579850 360884 580094
rect 362972 579986 363000 700878
rect 364340 700664 364392 700670
rect 364340 700606 364392 700612
rect 364352 580122 364380 700606
rect 365180 687818 365208 703446
rect 367100 700732 367152 700738
rect 367100 700674 367152 700680
rect 364616 687812 364668 687818
rect 364616 687754 364668 687760
rect 365168 687812 365220 687818
rect 365168 687754 365220 687760
rect 364628 685846 364656 687754
rect 364616 685840 364668 685846
rect 364616 685782 364668 685788
rect 364524 676252 364576 676258
rect 364524 676194 364576 676200
rect 364536 669338 364564 676194
rect 364536 669310 364748 669338
rect 364720 650026 364748 669310
rect 364536 649998 364748 650026
rect 364536 630714 364564 649998
rect 364536 630686 364656 630714
rect 364628 618254 364656 630686
rect 364616 618248 364668 618254
rect 364616 618190 364668 618196
rect 364524 608660 364576 608666
rect 364524 608602 364576 608608
rect 364536 601746 364564 608602
rect 364536 601718 364656 601746
rect 364628 598942 364656 601718
rect 364616 598936 364668 598942
rect 364616 598878 364668 598884
rect 364708 589348 364760 589354
rect 364708 589290 364760 589296
rect 364720 584730 364748 589290
rect 364708 584724 364760 584730
rect 364708 584666 364760 584672
rect 364352 580094 365208 580122
rect 365180 579986 365208 580094
rect 362972 579958 363446 579986
rect 365180 579958 365562 579986
rect 367112 579850 367140 700674
rect 368480 700596 368532 700602
rect 368480 700538 368532 700544
rect 368492 580122 368520 700538
rect 374000 700528 374052 700534
rect 374000 700470 374052 700476
rect 371240 700460 371292 700466
rect 371240 700402 371292 700408
rect 368492 580094 369348 580122
rect 369320 579850 369348 580094
rect 371252 579850 371280 700402
rect 374012 579972 374040 700470
rect 375380 700392 375432 700398
rect 375380 700334 375432 700340
rect 378138 700360 378194 700369
rect 375392 579850 375420 700334
rect 378138 700295 378194 700304
rect 379520 700324 379572 700330
rect 378152 579986 378180 700295
rect 379520 700266 379572 700272
rect 378152 579958 378258 579986
rect 379532 579850 379560 700266
rect 397472 699786 397500 703520
rect 413664 699854 413692 703520
rect 413652 699848 413704 699854
rect 413652 699790 413704 699796
rect 397460 699780 397512 699786
rect 397460 699722 397512 699728
rect 429856 688634 429884 703520
rect 462332 700126 462360 703520
rect 478524 700194 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 462320 700120 462372 700126
rect 462320 700062 462372 700068
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700874 527220 703520
rect 527180 700868 527232 700874
rect 527180 700810 527232 700816
rect 543476 700806 543504 703520
rect 543464 700800 543516 700806
rect 543464 700742 543516 700748
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 382280 681760 382332 681766
rect 382280 681702 382332 681708
rect 382292 579986 382320 681702
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 386420 667956 386472 667962
rect 386420 667898 386472 667904
rect 383660 652792 383712 652798
rect 383660 652734 383712 652740
rect 382292 579958 382398 579986
rect 383672 579850 383700 652734
rect 386432 579986 386460 667898
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 429672 659682 429700 666538
rect 429488 659654 429700 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 429488 647290 429516 659654
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 494072 644450 494100 654094
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 387800 623824 387852 623830
rect 387800 623766 387852 623772
rect 386432 579958 386630 579986
rect 387812 579850 387840 623766
rect 429396 621058 429424 630550
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 429396 621030 429516 621058
rect 429488 611386 429516 621030
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 391940 610020 391992 610026
rect 391940 609962 391992 609968
rect 390560 594856 390612 594862
rect 390560 594798 390612 594804
rect 390572 579986 390600 594798
rect 391952 580122 391980 609962
rect 429396 608598 429424 611238
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 494256 596222 494284 605798
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 429672 584594 429700 589290
rect 429660 584588 429712 584594
rect 429660 584530 429712 584536
rect 494256 584526 494284 596006
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 494244 584520 494296 584526
rect 494244 584462 494296 584468
rect 559392 584458 559420 589290
rect 559380 584452 559432 584458
rect 559380 584394 559432 584400
rect 471336 583704 471388 583710
rect 471336 583646 471388 583652
rect 471244 583636 471296 583642
rect 471244 583578 471296 583584
rect 460294 583536 460350 583545
rect 460294 583471 460350 583480
rect 399208 583364 399260 583370
rect 399208 583306 399260 583312
rect 395068 580168 395120 580174
rect 391952 580094 392532 580122
rect 395068 580110 395120 580116
rect 390572 579958 390862 579986
rect 392504 579850 392532 580094
rect 395080 579972 395108 580110
rect 397092 580100 397144 580106
rect 397092 580042 397144 580048
rect 397104 579972 397132 580042
rect 399220 579972 399248 583306
rect 405556 583296 405608 583302
rect 405556 583238 405608 583244
rect 400956 580032 401008 580038
rect 401008 579980 401350 579986
rect 400956 579974 401350 579980
rect 400968 579958 401350 579974
rect 403176 579970 403466 579986
rect 405568 579972 405596 583238
rect 411904 583228 411956 583234
rect 411904 583170 411956 583176
rect 409788 583160 409840 583166
rect 409788 583102 409840 583108
rect 407672 583092 407724 583098
rect 407672 583034 407724 583040
rect 407684 579972 407712 583034
rect 409800 579972 409828 583102
rect 411916 579972 411944 583170
rect 420274 583128 420330 583137
rect 420274 583063 420330 583072
rect 418160 583024 418212 583030
rect 418160 582966 418212 582972
rect 414020 582888 414072 582894
rect 414020 582830 414072 582836
rect 414032 579972 414060 582830
rect 418172 579972 418200 582966
rect 420288 579972 420316 583063
rect 426622 582992 426678 583001
rect 424508 582956 424560 582962
rect 426622 582927 426678 582936
rect 424508 582898 424560 582904
rect 422392 582820 422444 582826
rect 422392 582762 422444 582768
rect 422404 579972 422432 582762
rect 424520 579972 424548 582898
rect 426636 579972 426664 582927
rect 449806 582856 449862 582865
rect 449806 582791 449862 582800
rect 437112 582752 437164 582758
rect 437112 582694 437164 582700
rect 430856 582684 430908 582690
rect 430856 582626 430908 582632
rect 430868 579972 430896 582626
rect 432972 582616 433024 582622
rect 432972 582558 433024 582564
rect 432984 579972 433012 582558
rect 434996 582548 435048 582554
rect 434996 582490 435048 582496
rect 435008 579972 435036 582490
rect 437124 579972 437152 582694
rect 447690 582584 447746 582593
rect 447690 582519 447746 582528
rect 445576 582480 445628 582486
rect 445576 582422 445628 582428
rect 443460 582412 443512 582418
rect 443460 582354 443512 582360
rect 443472 579972 443500 582354
rect 445588 579972 445616 582422
rect 447704 579972 447732 582519
rect 449820 579972 449848 582791
rect 460308 579972 460336 583471
rect 462410 582720 462466 582729
rect 462410 582655 462466 582664
rect 462424 579972 462452 582655
rect 469588 581528 469640 581534
rect 469588 581470 469640 581476
rect 403164 579964 403466 579970
rect 403216 579958 403466 579964
rect 403164 579906 403216 579912
rect 438860 579896 438912 579902
rect 347792 579822 348726 579850
rect 351932 579822 352958 579850
rect 356072 579822 357190 579850
rect 358832 579822 359306 579850
rect 360856 579822 361330 579850
rect 367112 579822 367678 579850
rect 369320 579822 369794 579850
rect 371252 579822 371910 579850
rect 375392 579822 376142 579850
rect 379532 579822 380282 579850
rect 383672 579822 384514 579850
rect 387812 579822 388746 579850
rect 392504 579822 392978 579850
rect 438912 579844 439254 579850
rect 438860 579838 439254 579844
rect 438872 579822 439254 579838
rect 451568 579834 451950 579850
rect 451556 579828 451950 579834
rect 451608 579822 451950 579828
rect 451556 579770 451608 579776
rect 458272 579760 458324 579766
rect 458206 579708 458272 579714
rect 468482 579728 468538 579737
rect 458206 579702 458324 579708
rect 458206 579686 458312 579702
rect 464264 579698 464554 579714
rect 464252 579692 464554 579698
rect 464304 579686 464554 579692
rect 468538 579686 468786 579714
rect 468482 579663 468538 579672
rect 464252 579634 464304 579640
rect 270802 579426 271184 579442
rect 270802 579420 271196 579426
rect 270802 579414 271144 579420
rect 271144 579362 271196 579368
rect 247960 579352 248012 579358
rect 231122 579320 231178 579329
rect 230874 579278 231122 579306
rect 232962 579320 233018 579329
rect 232898 579278 232962 579306
rect 231122 579255 231178 579264
rect 235262 579320 235318 579329
rect 235014 579278 235262 579306
rect 232962 579255 233018 579264
rect 237194 579320 237250 579329
rect 237130 579278 237194 579306
rect 235262 579255 235318 579264
rect 239402 579320 239458 579329
rect 239246 579278 239402 579306
rect 237194 579255 237250 579264
rect 241426 579320 241482 579329
rect 241362 579278 241426 579306
rect 239402 579255 239458 579264
rect 243634 579320 243690 579329
rect 243478 579278 243634 579306
rect 241426 579255 241482 579264
rect 247710 579300 247960 579306
rect 254216 579352 254268 579358
rect 247710 579294 248012 579300
rect 249522 579320 249578 579329
rect 247710 579278 248000 579294
rect 243634 579255 243690 579264
rect 249578 579278 249734 579306
rect 253966 579300 254216 579306
rect 258448 579352 258500 579358
rect 253966 579294 254268 579300
rect 258198 579300 258448 579306
rect 260656 579352 260708 579358
rect 258198 579294 258500 579300
rect 260314 579300 260656 579306
rect 266912 579352 266964 579358
rect 260314 579294 260708 579300
rect 266662 579300 266912 579306
rect 273168 579352 273220 579358
rect 266662 579294 266964 579300
rect 272918 579300 273168 579306
rect 277308 579352 277360 579358
rect 272918 579294 273220 579300
rect 277150 579300 277308 579306
rect 279608 579352 279660 579358
rect 277150 579294 277360 579300
rect 279266 579300 279608 579306
rect 285772 579352 285824 579358
rect 279266 579294 279660 579300
rect 285614 579300 285772 579306
rect 292120 579352 292172 579358
rect 285614 579294 285824 579300
rect 291870 579300 292120 579306
rect 291870 579294 292172 579300
rect 415676 579352 415728 579358
rect 428372 579352 428424 579358
rect 415728 579300 416070 579306
rect 415676 579294 416070 579300
rect 441068 579352 441120 579358
rect 428424 579300 428766 579306
rect 428372 579294 428766 579300
rect 453580 579352 453632 579358
rect 441120 579300 441370 579306
rect 441068 579294 441370 579300
rect 455788 579352 455840 579358
rect 453632 579300 453974 579306
rect 453580 579294 453974 579300
rect 466458 579320 466514 579329
rect 455840 579300 456090 579306
rect 455788 579294 456090 579300
rect 253966 579278 254256 579294
rect 258198 579278 258488 579294
rect 260314 579278 260696 579294
rect 266662 579278 266952 579294
rect 272918 579278 273208 579294
rect 277150 579278 277348 579294
rect 279266 579278 279648 579294
rect 285614 579278 285812 579294
rect 291870 579278 292160 579294
rect 415688 579278 416070 579294
rect 428384 579278 428766 579294
rect 441080 579278 441370 579294
rect 453592 579278 453974 579294
rect 455800 579278 456090 579294
rect 249522 579255 249578 579264
rect 466514 579278 466670 579306
rect 466458 579255 466514 579264
rect 469600 557530 469628 581470
rect 469680 581460 469732 581466
rect 469680 581402 469732 581408
rect 469588 557524 469640 557530
rect 469588 557466 469640 557472
rect 469692 510610 469720 581402
rect 469772 581392 469824 581398
rect 469772 581334 469824 581340
rect 469680 510604 469732 510610
rect 469680 510546 469732 510552
rect 469784 463690 469812 581334
rect 470508 581324 470560 581330
rect 470508 581266 470560 581272
rect 470416 581256 470468 581262
rect 470416 581198 470468 581204
rect 470232 581188 470284 581194
rect 470232 581130 470284 581136
rect 470140 581120 470192 581126
rect 470140 581062 470192 581068
rect 469956 580372 470008 580378
rect 469956 580314 470008 580320
rect 469864 580304 469916 580310
rect 469864 580246 469916 580252
rect 469772 463684 469824 463690
rect 469772 463626 469824 463632
rect 232516 340190 232898 340218
rect 244752 340190 245226 340218
rect 246224 340190 246698 340218
rect 290292 340190 290766 340218
rect 291764 340190 292238 340218
rect 294708 340190 295182 340218
rect 326540 340190 327014 340218
rect 330496 340190 330878 340218
rect 386800 340190 387274 340218
rect 389744 340190 390218 340218
rect 392610 340190 393084 340218
rect 422970 340190 423444 340218
rect 438150 340190 438624 340218
rect 229112 340054 230046 340082
rect 230506 340054 230612 340082
rect 71044 338088 71096 338094
rect 71044 338030 71096 338036
rect 66904 338020 66956 338026
rect 66904 337962 66956 337968
rect 61384 337952 61436 337958
rect 61384 337894 61436 337900
rect 57244 337884 57296 337890
rect 57244 337826 57296 337832
rect 50344 337816 50396 337822
rect 50344 337758 50396 337764
rect 39304 337748 39356 337754
rect 39304 337690 39356 337696
rect 32404 337680 32456 337686
rect 32404 337622 32456 337628
rect 28264 337544 28316 337550
rect 28264 337486 28316 337492
rect 24124 64864 24176 64870
rect 24124 64806 24176 64812
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20732 480 20760 4014
rect 21928 480 21956 7686
rect 23400 610 23428 11698
rect 27896 9104 27948 9110
rect 27896 9046 27948 9052
rect 26700 7812 26752 7818
rect 26700 7754 26752 7760
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3606
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25516 480 25544 3538
rect 26712 480 26740 7754
rect 27908 480 27936 9046
rect 28276 4078 28304 337486
rect 31668 13116 31720 13122
rect 31668 13058 31720 13064
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 480 29132 3334
rect 30300 480 30328 7822
rect 31680 626 31708 13058
rect 32416 3806 32444 337622
rect 35164 337612 35216 337618
rect 35164 337554 35216 337560
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3674
rect 33888 480 33916 7890
rect 34980 4140 35032 4146
rect 34980 4082 35032 4088
rect 34992 480 35020 4082
rect 35176 3398 35204 337554
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36188 480 36216 3334
rect 37384 480 37412 7958
rect 38568 3800 38620 3806
rect 38568 3742 38620 3748
rect 38580 480 38608 3742
rect 39316 3398 39344 337690
rect 49332 9240 49384 9246
rect 49332 9182 49384 9188
rect 44548 9172 44600 9178
rect 44548 9114 44600 9120
rect 40960 8084 41012 8090
rect 40960 8026 41012 8032
rect 39764 3868 39816 3874
rect 39764 3810 39816 3816
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39776 480 39804 3810
rect 40972 480 41000 8026
rect 42156 3324 42208 3330
rect 42156 3266 42208 3272
rect 42168 480 42196 3266
rect 43352 3188 43404 3194
rect 43352 3130 43404 3136
rect 43364 480 43392 3130
rect 44560 480 44588 9114
rect 48136 5228 48188 5234
rect 48136 5170 48188 5176
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45756 480 45784 3878
rect 46952 480 46980 3946
rect 48148 480 48176 5170
rect 49344 480 49372 9182
rect 50356 4146 50384 337758
rect 56508 10396 56560 10402
rect 56508 10338 56560 10344
rect 53748 10328 53800 10334
rect 53748 10270 53800 10276
rect 51630 6216 51686 6225
rect 51630 6151 51686 6160
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50540 480 50568 4014
rect 51644 480 51672 6151
rect 53760 3262 53788 10270
rect 55220 6180 55272 6186
rect 55220 6122 55272 6128
rect 52828 3256 52880 3262
rect 52828 3198 52880 3204
rect 53748 3256 53800 3262
rect 53748 3198 53800 3204
rect 54024 3256 54076 3262
rect 54024 3198 54076 3204
rect 52840 480 52868 3198
rect 54036 480 54064 3198
rect 55232 480 55260 6122
rect 56520 3482 56548 10338
rect 56428 3454 56548 3482
rect 56428 480 56456 3454
rect 57256 3330 57284 337826
rect 57978 337784 58034 337793
rect 57978 337719 57980 337728
rect 58032 337719 58034 337728
rect 57980 337690 58032 337696
rect 60648 10464 60700 10470
rect 60648 10406 60700 10412
rect 58808 6248 58860 6254
rect 58808 6190 58860 6196
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57624 480 57652 4082
rect 58820 480 58848 6190
rect 60660 3398 60688 10406
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61396 3330 61424 337894
rect 64788 10532 64840 10538
rect 64788 10474 64840 10480
rect 62396 6316 62448 6322
rect 62396 6258 62448 6264
rect 61384 3324 61436 3330
rect 61384 3266 61436 3272
rect 61200 3188 61252 3194
rect 61200 3130 61252 3136
rect 61212 480 61240 3130
rect 62408 480 62436 6258
rect 64800 3398 64828 10474
rect 65984 6384 66036 6390
rect 65984 6326 66036 6332
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 63604 480 63632 3334
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64800 480 64828 3198
rect 65996 480 66024 6326
rect 66916 3126 66944 337962
rect 67546 337784 67602 337793
rect 67546 337719 67548 337728
rect 67600 337719 67602 337728
rect 67548 337690 67600 337696
rect 69480 6452 69532 6458
rect 69480 6394 69532 6400
rect 67180 5296 67232 5302
rect 67180 5238 67232 5244
rect 66904 3120 66956 3126
rect 66904 3062 66956 3068
rect 67192 480 67220 5238
rect 68284 3188 68336 3194
rect 68284 3130 68336 3136
rect 68296 480 68324 3130
rect 69492 480 69520 6394
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 70688 480 70716 3334
rect 71056 3126 71084 338030
rect 77298 337784 77354 337793
rect 77298 337719 77300 337728
rect 77352 337719 77354 337728
rect 86866 337784 86922 337793
rect 86866 337719 86868 337728
rect 77300 337690 77352 337696
rect 86920 337719 86922 337728
rect 95238 337784 95294 337793
rect 95238 337719 95240 337728
rect 86868 337690 86920 337696
rect 95292 337719 95294 337728
rect 104806 337784 104862 337793
rect 104806 337719 104808 337728
rect 95240 337690 95292 337696
rect 104860 337719 104862 337728
rect 114558 337784 114614 337793
rect 114558 337719 114560 337728
rect 104808 337690 104860 337696
rect 114612 337719 114614 337728
rect 124126 337784 124182 337793
rect 124126 337719 124128 337728
rect 114560 337690 114612 337696
rect 124180 337719 124182 337728
rect 133878 337784 133934 337793
rect 133878 337719 133880 337728
rect 124128 337690 124180 337696
rect 133932 337719 133934 337728
rect 143446 337784 143502 337793
rect 143446 337719 143448 337728
rect 133880 337690 133932 337696
rect 143500 337719 143502 337728
rect 153198 337784 153254 337793
rect 153198 337719 153200 337728
rect 143448 337690 143500 337696
rect 153252 337719 153254 337728
rect 162766 337784 162822 337793
rect 162766 337719 162768 337728
rect 153200 337690 153252 337696
rect 162820 337719 162822 337728
rect 172518 337784 172574 337793
rect 172518 337719 172520 337728
rect 162768 337690 162820 337696
rect 172572 337719 172574 337728
rect 182086 337784 182142 337793
rect 182086 337719 182088 337728
rect 172520 337690 172572 337696
rect 182140 337719 182142 337728
rect 191838 337784 191894 337793
rect 191838 337719 191840 337728
rect 182088 337690 182140 337696
rect 191892 337719 191894 337728
rect 201406 337784 201462 337793
rect 201406 337719 201408 337728
rect 191840 337690 191892 337696
rect 201460 337719 201462 337728
rect 211158 337784 211214 337793
rect 211158 337719 211160 337728
rect 201408 337690 201460 337696
rect 211212 337719 211214 337728
rect 220726 337784 220782 337793
rect 220726 337719 220728 337728
rect 211160 337690 211212 337696
rect 220780 337719 220782 337728
rect 220728 337690 220780 337696
rect 220832 337606 221044 337634
rect 220832 337550 220860 337606
rect 221016 337550 221044 337606
rect 220820 337544 220872 337550
rect 220820 337486 220872 337492
rect 221004 337544 221056 337550
rect 221004 337486 221056 337492
rect 220820 337408 220872 337414
rect 221004 337408 221056 337414
rect 220872 337356 221004 337362
rect 220820 337350 221056 337356
rect 79324 337340 79376 337346
rect 220832 337334 221044 337350
rect 79324 337282 79376 337288
rect 77944 337000 77996 337006
rect 77944 336942 77996 336948
rect 74448 14476 74500 14482
rect 74448 14418 74500 14424
rect 71688 13184 71740 13190
rect 71688 13126 71740 13132
rect 71700 3398 71728 13126
rect 73068 6520 73120 6526
rect 73068 6462 73120 6468
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71044 3120 71096 3126
rect 71044 3062 71096 3068
rect 71884 480 71912 3266
rect 73080 480 73108 6462
rect 74460 3380 74488 14418
rect 76656 6588 76708 6594
rect 76656 6530 76708 6536
rect 74276 3352 74488 3380
rect 74276 480 74304 3352
rect 75460 3188 75512 3194
rect 75460 3130 75512 3136
rect 75472 480 75500 3130
rect 76668 480 76696 6530
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 77864 480 77892 3198
rect 77956 3058 77984 336942
rect 78588 14544 78640 14550
rect 78588 14486 78640 14492
rect 78600 3262 78628 14486
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 79336 3194 79364 337282
rect 132500 337272 132552 337278
rect 132498 337240 132500 337249
rect 142068 337272 142120 337278
rect 132552 337240 132554 337249
rect 84844 337204 84896 337210
rect 132498 337175 132554 337184
rect 142066 337240 142068 337249
rect 151820 337272 151872 337278
rect 142120 337240 142122 337249
rect 142066 337175 142122 337184
rect 151818 337240 151820 337249
rect 161388 337272 161440 337278
rect 151872 337240 151874 337249
rect 151818 337175 151874 337184
rect 161386 337240 161388 337249
rect 171140 337272 171192 337278
rect 161440 337240 161442 337249
rect 161386 337175 161442 337184
rect 171138 337240 171140 337249
rect 180708 337272 180760 337278
rect 171192 337240 171194 337249
rect 171138 337175 171194 337184
rect 180706 337240 180708 337249
rect 190460 337272 190512 337278
rect 180760 337240 180762 337249
rect 180706 337175 180762 337184
rect 190458 337240 190460 337249
rect 200028 337272 200080 337278
rect 190512 337240 190514 337249
rect 190458 337175 190514 337184
rect 200026 337240 200028 337249
rect 209780 337272 209832 337278
rect 200080 337240 200082 337249
rect 200026 337175 200082 337184
rect 209778 337240 209780 337249
rect 219348 337272 219400 337278
rect 209832 337240 209834 337249
rect 209778 337175 209834 337184
rect 219346 337240 219348 337249
rect 221004 337272 221056 337278
rect 219400 337240 219402 337249
rect 219346 337175 219402 337184
rect 221002 337240 221004 337249
rect 221056 337240 221058 337249
rect 221002 337175 221058 337184
rect 84844 337146 84896 337152
rect 82728 14612 82780 14618
rect 82728 14554 82780 14560
rect 80244 8152 80296 8158
rect 80244 8094 80296 8100
rect 79324 3188 79376 3194
rect 79324 3130 79376 3136
rect 77944 3052 77996 3058
rect 77944 2994 77996 3000
rect 79048 2984 79100 2990
rect 79048 2926 79100 2932
rect 79060 480 79088 2926
rect 80256 480 80284 8094
rect 82740 3262 82768 14554
rect 83832 8220 83884 8226
rect 83832 8162 83884 8168
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 81452 480 81480 3198
rect 82636 3188 82688 3194
rect 82636 3130 82688 3136
rect 82648 480 82676 3130
rect 83844 480 83872 8162
rect 84856 3262 84884 337146
rect 100668 337136 100720 337142
rect 100668 337078 100720 337084
rect 95884 337068 95936 337074
rect 95884 337010 95936 337016
rect 92388 14816 92440 14822
rect 92388 14758 92440 14764
rect 89628 14748 89680 14754
rect 89628 14690 89680 14696
rect 85488 14680 85540 14686
rect 85488 14622 85540 14628
rect 85500 3262 85528 14622
rect 87328 8288 87380 8294
rect 87328 8230 87380 8236
rect 84844 3256 84896 3262
rect 84844 3198 84896 3204
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84948 480 84976 3198
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 86144 480 86172 2926
rect 87340 480 87368 8230
rect 89640 3262 89668 14690
rect 91008 10600 91060 10606
rect 91008 10542 91060 10548
rect 91020 3482 91048 10542
rect 92400 3482 92428 14758
rect 95148 10668 95200 10674
rect 95148 10610 95200 10616
rect 90928 3454 91048 3482
rect 92124 3454 92428 3482
rect 88524 3256 88576 3262
rect 88524 3198 88576 3204
rect 89628 3256 89680 3262
rect 89628 3198 89680 3204
rect 88536 480 88564 3198
rect 89720 3120 89772 3126
rect 89720 3062 89772 3068
rect 89732 480 89760 3062
rect 90928 480 90956 3454
rect 92124 480 92152 3454
rect 95160 3126 95188 10610
rect 94504 3120 94556 3126
rect 94504 3062 94556 3068
rect 95148 3120 95200 3126
rect 95148 3062 95200 3068
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 93308 3052 93360 3058
rect 93308 2994 93360 3000
rect 93320 480 93348 2994
rect 94516 480 94544 3062
rect 95712 480 95740 3062
rect 95896 2854 95924 337010
rect 99288 14952 99340 14958
rect 99288 14894 99340 14900
rect 96528 14884 96580 14890
rect 96528 14826 96580 14832
rect 96540 3126 96568 14826
rect 99196 10736 99248 10742
rect 99196 10678 99248 10684
rect 99208 3126 99236 10678
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 98092 3120 98144 3126
rect 98092 3062 98144 3068
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 96896 2984 96948 2990
rect 96896 2926 96948 2932
rect 95884 2848 95936 2854
rect 95884 2790 95936 2796
rect 96908 480 96936 2926
rect 98104 480 98132 3062
rect 99300 480 99328 14894
rect 100680 3482 100708 337078
rect 107568 337000 107620 337006
rect 107568 336942 107620 336948
rect 102784 336932 102836 336938
rect 102784 336874 102836 336880
rect 102048 10804 102100 10810
rect 102048 10746 102100 10752
rect 100496 3454 100708 3482
rect 100496 480 100524 3454
rect 102060 3126 102088 10746
rect 102796 3210 102824 336874
rect 107476 15088 107528 15094
rect 107476 15030 107528 15036
rect 103428 15020 103480 15026
rect 103428 14962 103480 14968
rect 102612 3182 102824 3210
rect 101588 3120 101640 3126
rect 101588 3062 101640 3068
rect 102048 3120 102100 3126
rect 102048 3062 102100 3068
rect 101600 480 101628 3062
rect 102612 3058 102640 3182
rect 103440 3126 103468 14962
rect 106188 10872 106240 10878
rect 106188 10814 106240 10820
rect 106200 3126 106228 10814
rect 107488 3126 107516 15030
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 105176 3120 105228 3126
rect 105176 3062 105228 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 102600 3052 102652 3058
rect 102600 2994 102652 3000
rect 102796 480 102824 3062
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 103992 480 104020 2858
rect 105188 480 105216 3062
rect 106384 480 106412 3062
rect 107580 480 107608 336942
rect 118608 336864 118660 336870
rect 118608 336806 118660 336812
rect 110328 15156 110380 15162
rect 110328 15098 110380 15104
rect 108948 10940 109000 10946
rect 108948 10882 109000 10888
rect 108960 3482 108988 10882
rect 110340 3482 110368 15098
rect 114468 14408 114520 14414
rect 114468 14350 114520 14356
rect 113088 11008 113140 11014
rect 113088 10950 113140 10956
rect 108776 3454 108988 3482
rect 109972 3454 110368 3482
rect 108776 480 108804 3454
rect 109972 480 110000 3454
rect 113100 2990 113128 10950
rect 114480 2990 114508 14350
rect 117228 14340 117280 14346
rect 117228 14282 117280 14288
rect 117136 10260 117188 10266
rect 117136 10202 117188 10208
rect 117148 3618 117176 10202
rect 116964 3590 117176 3618
rect 116964 2990 116992 3590
rect 117240 3482 117268 14282
rect 117148 3454 117268 3482
rect 112352 2984 112404 2990
rect 112352 2926 112404 2932
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 115940 2984 115992 2990
rect 115940 2926 115992 2932
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 111168 480 111196 2858
rect 112364 480 112392 2926
rect 113560 480 113588 2926
rect 114744 2848 114796 2854
rect 114744 2790 114796 2796
rect 114756 480 114784 2790
rect 115952 480 115980 2926
rect 117148 480 117176 3454
rect 118620 3346 118648 336806
rect 125508 336796 125560 336802
rect 125508 336738 125560 336744
rect 121368 14272 121420 14278
rect 121368 14214 121420 14220
rect 119988 10192 120040 10198
rect 119988 10134 120040 10140
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 120000 2990 120028 10134
rect 121380 2990 121408 14214
rect 125416 14204 125468 14210
rect 125416 14146 125468 14152
rect 124128 10124 124180 10130
rect 124128 10066 124180 10072
rect 124140 3482 124168 10066
rect 125428 4214 125456 14146
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 123036 3454 124168 3482
rect 119436 2984 119488 2990
rect 119436 2926 119488 2932
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 119448 480 119476 2926
rect 120644 480 120672 2926
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 3454
rect 124232 480 124260 4150
rect 125520 3482 125548 336738
rect 183468 13796 183520 13802
rect 183468 13738 183520 13744
rect 179328 13660 179380 13666
rect 179328 13602 179380 13608
rect 176568 13592 176620 13598
rect 176568 13534 176620 13540
rect 172428 13524 172480 13530
rect 172428 13466 172480 13472
rect 168288 13456 168340 13462
rect 168288 13398 168340 13404
rect 165528 13388 165580 13394
rect 165528 13330 165580 13336
rect 160008 13320 160060 13326
rect 160008 13262 160060 13268
rect 155868 13252 155920 13258
rect 155868 13194 155920 13200
rect 151728 12164 151780 12170
rect 151728 12106 151780 12112
rect 148968 12096 149020 12102
rect 148968 12038 149020 12044
rect 144828 12028 144880 12034
rect 144828 11970 144880 11976
rect 142068 11960 142120 11966
rect 142068 11902 142120 11908
rect 128268 11892 128320 11898
rect 128268 11834 128320 11840
rect 126888 11824 126940 11830
rect 126888 11766 126940 11772
rect 126900 3482 126928 11766
rect 128280 3482 128308 11834
rect 139676 9376 139728 9382
rect 139676 9318 139728 9324
rect 136088 9308 136140 9314
rect 136088 9250 136140 9256
rect 132590 8936 132646 8945
rect 132590 8871 132646 8880
rect 129002 7576 129058 7585
rect 129002 7511 129058 7520
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 7511
rect 131396 6656 131448 6662
rect 131396 6598 131448 6604
rect 130200 5364 130252 5370
rect 130200 5306 130252 5312
rect 130212 480 130240 5306
rect 131408 480 131436 6598
rect 132604 480 132632 8871
rect 134892 7540 134944 7546
rect 134892 7482 134944 7488
rect 133788 5432 133840 5438
rect 133788 5374 133840 5380
rect 133800 480 133828 5374
rect 134904 480 134932 7482
rect 136100 480 136128 9250
rect 138480 7472 138532 7478
rect 138480 7414 138532 7420
rect 137284 5500 137336 5506
rect 137284 5442 137336 5448
rect 137296 480 137324 5442
rect 138492 480 138520 7414
rect 139688 480 139716 9318
rect 141976 7404 142028 7410
rect 141976 7346 142028 7352
rect 140872 4208 140924 4214
rect 140872 4150 140924 4156
rect 140884 480 140912 4150
rect 141988 3482 142016 7346
rect 142080 4214 142108 11902
rect 143448 10056 143500 10062
rect 143448 9998 143500 10004
rect 142068 4208 142120 4214
rect 142068 4150 142120 4156
rect 143460 3482 143488 9998
rect 144840 3482 144868 11970
rect 147588 9988 147640 9994
rect 147588 9930 147640 9936
rect 145656 7336 145708 7342
rect 145656 7278 145708 7284
rect 141988 3454 142108 3482
rect 142080 480 142108 3454
rect 143276 3454 143488 3482
rect 144472 3454 144868 3482
rect 143276 480 143304 3454
rect 144472 480 144500 3454
rect 145668 480 145696 7278
rect 147600 3482 147628 9930
rect 148980 3482 149008 12038
rect 151636 9920 151688 9926
rect 151636 9862 151688 9868
rect 149244 7268 149296 7274
rect 149244 7210 149296 7216
rect 146864 3454 147628 3482
rect 148060 3454 149008 3482
rect 146864 480 146892 3454
rect 148060 480 148088 3454
rect 149256 480 149284 7210
rect 151648 4214 151676 9862
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 150452 480 150480 4150
rect 151740 3482 151768 12106
rect 154488 9852 154540 9858
rect 154488 9794 154540 9800
rect 152740 7200 152792 7206
rect 152740 7142 152792 7148
rect 151556 3454 151768 3482
rect 151556 480 151584 3454
rect 152752 480 152780 7142
rect 154500 3482 154528 9794
rect 155880 3482 155908 13194
rect 158628 9784 158680 9790
rect 158628 9726 158680 9732
rect 156328 7132 156380 7138
rect 156328 7074 156380 7080
rect 153948 3454 154528 3482
rect 155144 3454 155908 3482
rect 153948 480 153976 3454
rect 155144 480 155172 3454
rect 156340 480 156368 7074
rect 158640 3482 158668 9726
rect 159916 7064 159968 7070
rect 159916 7006 159968 7012
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 157536 3454 158668 3482
rect 157536 480 157564 3454
rect 158732 480 158760 4150
rect 159928 480 159956 7006
rect 160020 4214 160048 13262
rect 162768 12232 162820 12238
rect 162768 12174 162820 12180
rect 161388 9716 161440 9722
rect 161388 9658 161440 9664
rect 160008 4208 160060 4214
rect 160008 4150 160060 4156
rect 161400 3482 161428 9658
rect 161124 3454 161428 3482
rect 161124 480 161152 3454
rect 162780 626 162808 12174
rect 163504 6724 163556 6730
rect 163504 6666 163556 6672
rect 162320 598 162808 626
rect 162320 480 162348 598
rect 163516 480 163544 6666
rect 165540 610 165568 13330
rect 166908 12300 166960 12306
rect 166908 12242 166960 12248
rect 166920 610 166948 12242
rect 167092 6792 167144 6798
rect 167092 6734 167144 6740
rect 164700 604 164752 610
rect 164700 546 164752 552
rect 165528 604 165580 610
rect 165528 546 165580 552
rect 165896 604 165948 610
rect 165896 546 165948 552
rect 166908 604 166960 610
rect 166908 546 166960 552
rect 164712 480 164740 546
rect 165908 480 165936 546
rect 167104 480 167132 6734
rect 168300 626 168328 13398
rect 169668 12368 169720 12374
rect 169668 12310 169720 12316
rect 168208 598 168328 626
rect 169680 610 169708 12310
rect 170588 6860 170640 6866
rect 170588 6802 170640 6808
rect 169392 604 169444 610
rect 168208 480 168236 598
rect 169392 546 169444 552
rect 169668 604 169720 610
rect 169668 546 169720 552
rect 169404 480 169432 546
rect 170600 480 170628 6802
rect 172440 3346 172468 13466
rect 173808 12436 173860 12442
rect 173808 12378 173860 12384
rect 173820 3346 173848 12378
rect 176476 11688 176528 11694
rect 176476 11630 176528 11636
rect 174176 6112 174228 6118
rect 174176 6054 174228 6060
rect 171796 3318 172468 3346
rect 172992 3318 173848 3346
rect 171796 480 171824 3318
rect 172992 480 173020 3318
rect 174188 480 174216 6054
rect 175372 4208 175424 4214
rect 175372 4150 175424 4156
rect 175384 480 175412 4150
rect 176488 3482 176516 11630
rect 176580 4214 176608 13534
rect 177764 6044 177816 6050
rect 177764 5986 177816 5992
rect 176568 4208 176620 4214
rect 176568 4150 176620 4156
rect 176488 3454 176608 3482
rect 176580 480 176608 3454
rect 177776 480 177804 5986
rect 179340 3346 179368 13602
rect 180708 11620 180760 11626
rect 180708 11562 180760 11568
rect 180720 3346 180748 11562
rect 181352 5976 181404 5982
rect 181352 5918 181404 5924
rect 178972 3318 179368 3346
rect 180168 3318 180748 3346
rect 178972 480 179000 3318
rect 180168 480 180196 3318
rect 181364 480 181392 5918
rect 183480 610 183508 13738
rect 186228 13728 186280 13734
rect 186228 13670 186280 13676
rect 184848 11552 184900 11558
rect 184848 11494 184900 11500
rect 184860 6066 184888 11494
rect 184768 6038 184888 6066
rect 184768 610 184796 6038
rect 184848 5908 184900 5914
rect 184848 5850 184900 5856
rect 182548 604 182600 610
rect 182548 546 182600 552
rect 183468 604 183520 610
rect 183468 546 183520 552
rect 183744 604 183796 610
rect 183744 546 183796 552
rect 184756 604 184808 610
rect 184756 546 184808 552
rect 182560 480 182588 546
rect 183756 480 183784 546
rect 184860 480 184888 5850
rect 186240 626 186268 13670
rect 190368 13048 190420 13054
rect 190368 12990 190420 12996
rect 187608 11484 187660 11490
rect 187608 11426 187660 11432
rect 186056 598 186268 626
rect 187620 610 187648 11426
rect 188436 5840 188488 5846
rect 188436 5782 188488 5788
rect 187240 604 187292 610
rect 186056 480 186084 598
rect 187240 546 187292 552
rect 187608 604 187660 610
rect 187608 546 187660 552
rect 187252 480 187280 546
rect 188448 480 188476 5782
rect 190380 610 190408 12990
rect 206928 12980 206980 12986
rect 206928 12922 206980 12928
rect 191748 11416 191800 11422
rect 191748 11358 191800 11364
rect 191760 3346 191788 11358
rect 194508 11348 194560 11354
rect 194508 11290 194560 11296
rect 193220 9444 193272 9450
rect 193220 9386 193272 9392
rect 192024 5772 192076 5778
rect 192024 5714 192076 5720
rect 190840 3318 191788 3346
rect 189632 604 189684 610
rect 189632 546 189684 552
rect 190368 604 190420 610
rect 190368 546 190420 552
rect 189644 480 189672 546
rect 190840 480 190868 3318
rect 192036 480 192064 5714
rect 193232 480 193260 9386
rect 194520 3482 194548 11290
rect 198648 11280 198700 11286
rect 198648 11222 198700 11228
rect 196808 9512 196860 9518
rect 196808 9454 196860 9460
rect 195612 5704 195664 5710
rect 195612 5646 195664 5652
rect 194428 3454 194548 3482
rect 194428 480 194456 3454
rect 195624 480 195652 5646
rect 196820 480 196848 9454
rect 198660 3346 198688 11222
rect 203892 9648 203944 9654
rect 203892 9590 203944 9596
rect 200396 9580 200448 9586
rect 200396 9522 200448 9528
rect 199200 5636 199252 5642
rect 199200 5578 199252 5584
rect 198016 3318 198688 3346
rect 198016 480 198044 3318
rect 199212 480 199240 5578
rect 200408 480 200436 9522
rect 202696 5568 202748 5574
rect 202696 5510 202748 5516
rect 201500 4412 201552 4418
rect 201500 4354 201552 4360
rect 201512 480 201540 4354
rect 202708 480 202736 5510
rect 203904 480 203932 9590
rect 205088 4344 205140 4350
rect 205088 4286 205140 4292
rect 205100 480 205128 4286
rect 206940 3346 206968 12922
rect 211068 12912 211120 12918
rect 211068 12854 211120 12860
rect 207480 8900 207532 8906
rect 207480 8842 207532 8848
rect 206296 3318 206968 3346
rect 206296 480 206324 3318
rect 207492 480 207520 8842
rect 210976 8832 211028 8838
rect 210976 8774 211028 8780
rect 208674 4856 208730 4865
rect 208674 4791 208730 4800
rect 208688 480 208716 4791
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 209884 480 209912 4150
rect 210988 3482 211016 8774
rect 211080 4214 211108 12854
rect 213828 12844 213880 12850
rect 213828 12786 213880 12792
rect 212264 4752 212316 4758
rect 212264 4694 212316 4700
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 4694
rect 213840 3346 213868 12786
rect 217968 12776 218020 12782
rect 217968 12718 218020 12724
rect 214656 8764 214708 8770
rect 214656 8706 214708 8712
rect 213472 3318 213868 3346
rect 213472 480 213500 3318
rect 214668 480 214696 8706
rect 215852 4684 215904 4690
rect 215852 4626 215904 4632
rect 215864 480 215892 4626
rect 217980 3346 218008 12718
rect 220728 12708 220780 12714
rect 220728 12650 220780 12656
rect 218152 8696 218204 8702
rect 218152 8638 218204 8644
rect 217060 3318 218008 3346
rect 217060 480 217088 3318
rect 218164 480 218192 8638
rect 219348 4616 219400 4622
rect 219348 4558 219400 4564
rect 219360 480 219388 4558
rect 220740 3346 220768 12650
rect 224868 12640 224920 12646
rect 224868 12582 224920 12588
rect 221740 8628 221792 8634
rect 221740 8570 221792 8576
rect 220556 3318 220768 3346
rect 220556 480 220584 3318
rect 221752 480 221780 8570
rect 222936 4548 222988 4554
rect 222936 4490 222988 4496
rect 222948 480 222976 4490
rect 224880 3346 224908 12582
rect 229008 12572 229060 12578
rect 229008 12514 229060 12520
rect 225328 8560 225380 8566
rect 225328 8502 225380 8508
rect 224144 3318 224908 3346
rect 224144 480 224172 3318
rect 225340 480 225368 8502
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 227720 7608 227772 7614
rect 227720 7550 227772 7556
rect 226524 4480 226576 4486
rect 226524 4422 226576 4428
rect 226536 480 226564 4422
rect 227732 480 227760 7550
rect 228928 480 228956 8434
rect 229020 7614 229048 12514
rect 229008 7608 229060 7614
rect 229008 7550 229060 7556
rect 229112 4962 229140 340054
rect 229100 4956 229152 4962
rect 229100 4898 229152 4904
rect 230112 4888 230164 4894
rect 230112 4830 230164 4836
rect 230124 480 230152 4830
rect 230584 4282 230612 340054
rect 230768 340054 230966 340082
rect 231136 340054 231426 340082
rect 230664 337680 230716 337686
rect 230664 337622 230716 337628
rect 230676 7682 230704 337622
rect 230664 7676 230716 7682
rect 230664 7618 230716 7624
rect 230768 4826 230796 340054
rect 231136 337686 231164 340054
rect 231124 337680 231176 337686
rect 231124 337622 231176 337628
rect 231964 337385 231992 340068
rect 232056 340054 232438 340082
rect 231950 337376 232006 337385
rect 231950 337311 232006 337320
rect 231308 7608 231360 7614
rect 231308 7550 231360 7556
rect 230756 4820 230808 4826
rect 230756 4762 230808 4768
rect 230572 4276 230624 4282
rect 230572 4218 230624 4224
rect 231320 480 231348 7550
rect 232056 3369 232084 340054
rect 232516 337770 232544 340190
rect 232240 337742 232544 337770
rect 232240 318889 232268 337742
rect 232226 318880 232282 318889
rect 232226 318815 232282 318824
rect 232410 318880 232466 318889
rect 232410 318815 232466 318824
rect 232424 312610 232452 318815
rect 232332 312582 232452 312610
rect 232332 307766 232360 312582
rect 232320 307760 232372 307766
rect 232320 307702 232372 307708
rect 232320 298172 232372 298178
rect 232320 298114 232372 298120
rect 232332 298042 232360 298114
rect 232320 298036 232372 298042
rect 232320 297978 232372 297984
rect 232228 288448 232280 288454
rect 232228 288390 232280 288396
rect 232240 280226 232268 288390
rect 232228 280220 232280 280226
rect 232228 280162 232280 280168
rect 232320 280220 232372 280226
rect 232320 280162 232372 280168
rect 232332 278746 232360 280162
rect 232240 278718 232360 278746
rect 232240 270570 232268 278718
rect 232228 270564 232280 270570
rect 232228 270506 232280 270512
rect 232228 269136 232280 269142
rect 232228 269078 232280 269084
rect 232240 260914 232268 269078
rect 232228 260908 232280 260914
rect 232228 260850 232280 260856
rect 232320 260908 232372 260914
rect 232320 260850 232372 260856
rect 232332 251326 232360 260850
rect 232320 251320 232372 251326
rect 232320 251262 232372 251268
rect 232228 251116 232280 251122
rect 232228 251058 232280 251064
rect 232240 249801 232268 251058
rect 232226 249792 232282 249801
rect 232226 249727 232282 249736
rect 232502 249792 232558 249801
rect 232502 249727 232558 249736
rect 232516 240174 232544 249727
rect 232320 240168 232372 240174
rect 232320 240110 232372 240116
rect 232504 240168 232556 240174
rect 232504 240110 232556 240116
rect 232332 235362 232360 240110
rect 232240 235334 232360 235362
rect 232240 230489 232268 235334
rect 232226 230480 232282 230489
rect 232226 230415 232282 230424
rect 232502 230480 232558 230489
rect 232502 230415 232558 230424
rect 232516 220862 232544 230415
rect 232320 220856 232372 220862
rect 232320 220798 232372 220804
rect 232504 220856 232556 220862
rect 232504 220798 232556 220804
rect 232332 211274 232360 220798
rect 232320 211268 232372 211274
rect 232320 211210 232372 211216
rect 232228 209840 232280 209846
rect 232228 209782 232280 209788
rect 232240 190482 232268 209782
rect 232240 190454 232360 190482
rect 232332 186266 232360 190454
rect 232240 186238 232360 186266
rect 232240 176730 232268 186238
rect 232228 176724 232280 176730
rect 232228 176666 232280 176672
rect 232320 176656 232372 176662
rect 232320 176598 232372 176604
rect 232332 166954 232360 176598
rect 232240 166926 232360 166954
rect 232240 154578 232268 166926
rect 232240 154562 232360 154578
rect 232240 154556 232372 154562
rect 232240 154550 232320 154556
rect 232320 154498 232372 154504
rect 232332 154467 232360 154498
rect 232320 144968 232372 144974
rect 232320 144910 232372 144916
rect 232332 143546 232360 144910
rect 232320 143540 232372 143546
rect 232320 143482 232372 143488
rect 232320 125724 232372 125730
rect 232320 125666 232372 125672
rect 232332 124166 232360 125666
rect 232320 124160 232372 124166
rect 232320 124102 232372 124108
rect 232320 114572 232372 114578
rect 232320 114514 232372 114520
rect 232332 104854 232360 114514
rect 232320 104848 232372 104854
rect 232320 104790 232372 104796
rect 232320 95260 232372 95266
rect 232320 95202 232372 95208
rect 232332 85542 232360 95202
rect 232320 85536 232372 85542
rect 232320 85478 232372 85484
rect 232228 75948 232280 75954
rect 232228 75890 232280 75896
rect 232240 67674 232268 75890
rect 232240 67646 232360 67674
rect 232332 66230 232360 67646
rect 232320 66224 232372 66230
rect 232320 66166 232372 66172
rect 232228 48340 232280 48346
rect 232228 48282 232280 48288
rect 232240 48226 232268 48282
rect 232240 48198 232452 48226
rect 232424 38758 232452 48198
rect 232320 38752 232372 38758
rect 232320 38694 232372 38700
rect 232412 38752 232464 38758
rect 232412 38694 232464 38700
rect 232332 36122 232360 38694
rect 232240 36094 232360 36122
rect 232240 29034 232268 36094
rect 232228 29028 232280 29034
rect 232228 28970 232280 28976
rect 232412 29028 232464 29034
rect 232412 28970 232464 28976
rect 232424 19378 232452 28970
rect 232412 19372 232464 19378
rect 232412 19314 232464 19320
rect 232504 19236 232556 19242
rect 232504 19178 232556 19184
rect 232516 14142 232544 19178
rect 232136 14136 232188 14142
rect 232136 14078 232188 14084
rect 232504 14136 232556 14142
rect 232504 14078 232556 14084
rect 232148 5030 232176 14078
rect 232504 8424 232556 8430
rect 232504 8366 232556 8372
rect 232136 5024 232188 5030
rect 232136 4966 232188 4972
rect 232042 3360 232098 3369
rect 232042 3295 232098 3304
rect 232516 480 232544 8366
rect 233436 7002 233464 340068
rect 233528 340054 233910 340082
rect 233528 337414 233556 340054
rect 234356 337482 234384 340068
rect 234724 340054 234922 340082
rect 235000 340054 235382 340082
rect 235644 340054 235842 340082
rect 236394 340054 236500 340082
rect 234344 337476 234396 337482
rect 234344 337418 234396 337424
rect 233516 337408 233568 337414
rect 233516 337350 233568 337356
rect 233884 337408 233936 337414
rect 233884 337350 233936 337356
rect 233896 9110 233924 337350
rect 234620 337272 234672 337278
rect 234618 337240 234620 337249
rect 234672 337240 234674 337249
rect 234618 337175 234674 337184
rect 233884 9104 233936 9110
rect 233884 9046 233936 9052
rect 233424 6996 233476 7002
rect 233424 6938 233476 6944
rect 234724 5098 234752 340054
rect 235000 334642 235028 340054
rect 234816 334614 235028 334642
rect 234816 8974 234844 334614
rect 235644 334558 235672 340054
rect 236184 335708 236236 335714
rect 236184 335650 236236 335656
rect 236092 335640 236144 335646
rect 236092 335582 236144 335588
rect 234988 334552 235040 334558
rect 234988 334494 235040 334500
rect 235632 334552 235684 334558
rect 235632 334494 235684 334500
rect 235000 46918 235028 334494
rect 234988 46912 235040 46918
rect 234988 46854 235040 46860
rect 235080 37324 235132 37330
rect 235080 37266 235132 37272
rect 234804 8968 234856 8974
rect 234804 8910 234856 8916
rect 235092 8362 235120 37266
rect 236000 8968 236052 8974
rect 236000 8910 236052 8916
rect 234896 8356 234948 8362
rect 234896 8298 234948 8304
rect 235080 8356 235132 8362
rect 235080 8298 235132 8304
rect 234908 8242 234936 8298
rect 234908 8214 235028 8242
rect 234804 7676 234856 7682
rect 234804 7618 234856 7624
rect 234712 5092 234764 5098
rect 234712 5034 234764 5040
rect 233700 4820 233752 4826
rect 233700 4762 233752 4768
rect 233712 480 233740 4762
rect 234816 480 234844 7618
rect 235000 3466 235028 8214
rect 234988 3460 235040 3466
rect 234988 3402 235040 3408
rect 236012 480 236040 8910
rect 236104 5166 236132 335582
rect 236196 9042 236224 335650
rect 236472 321706 236500 340054
rect 236564 340054 236854 340082
rect 237024 340054 237314 340082
rect 236564 335646 236592 340054
rect 237024 335714 237052 340054
rect 237852 337550 237880 340068
rect 237840 337544 237892 337550
rect 237840 337486 237892 337492
rect 238312 337482 238340 340068
rect 238786 340054 238892 340082
rect 238300 337476 238352 337482
rect 238300 337418 238352 337424
rect 237012 335708 237064 335714
rect 237012 335650 237064 335656
rect 236552 335640 236604 335646
rect 236552 335582 236604 335588
rect 236460 321700 236512 321706
rect 236460 321642 236512 321648
rect 236460 318844 236512 318850
rect 236460 318786 236512 318792
rect 236472 317422 236500 318786
rect 236276 317416 236328 317422
rect 236276 317358 236328 317364
rect 236460 317416 236512 317422
rect 236460 317358 236512 317364
rect 236288 298110 236316 317358
rect 236276 298104 236328 298110
rect 236276 298046 236328 298052
rect 236276 288448 236328 288454
rect 236276 288390 236328 288396
rect 236288 282946 236316 288390
rect 236276 282940 236328 282946
rect 236276 282882 236328 282888
rect 236460 282804 236512 282810
rect 236460 282746 236512 282752
rect 236472 273290 236500 282746
rect 236276 273284 236328 273290
rect 236276 273226 236328 273232
rect 236460 273284 236512 273290
rect 236460 273226 236512 273232
rect 236288 263634 236316 273226
rect 236276 263628 236328 263634
rect 236276 263570 236328 263576
rect 236460 263492 236512 263498
rect 236460 263434 236512 263440
rect 236472 253978 236500 263434
rect 236276 253972 236328 253978
rect 236276 253914 236328 253920
rect 236460 253972 236512 253978
rect 236460 253914 236512 253920
rect 236288 244322 236316 253914
rect 236276 244316 236328 244322
rect 236276 244258 236328 244264
rect 236460 244180 236512 244186
rect 236460 244122 236512 244128
rect 236472 241482 236500 244122
rect 236472 241454 236592 241482
rect 236564 231946 236592 241454
rect 236276 231940 236328 231946
rect 236276 231882 236328 231888
rect 236552 231940 236604 231946
rect 236552 231882 236604 231888
rect 236288 225010 236316 231882
rect 236276 225004 236328 225010
rect 236276 224946 236328 224952
rect 236460 224868 236512 224874
rect 236460 224810 236512 224816
rect 236472 212634 236500 224810
rect 236276 212628 236328 212634
rect 236276 212570 236328 212576
rect 236460 212628 236512 212634
rect 236460 212570 236512 212576
rect 236288 193390 236316 212570
rect 236276 193384 236328 193390
rect 236276 193326 236328 193332
rect 236276 193248 236328 193254
rect 236276 193190 236328 193196
rect 236288 174010 236316 193190
rect 236276 174004 236328 174010
rect 236276 173946 236328 173952
rect 236276 173868 236328 173874
rect 236276 173810 236328 173816
rect 236288 172553 236316 173810
rect 236274 172544 236330 172553
rect 236274 172479 236330 172488
rect 236458 172544 236514 172553
rect 236458 172479 236514 172488
rect 236472 162858 236500 172479
rect 236276 162852 236328 162858
rect 236276 162794 236328 162800
rect 236460 162852 236512 162858
rect 236460 162794 236512 162800
rect 236288 147642 236316 162794
rect 236288 147614 236500 147642
rect 236472 135289 236500 147614
rect 236274 135280 236330 135289
rect 236274 135215 236330 135224
rect 236458 135280 236514 135289
rect 236458 135215 236514 135224
rect 236288 128330 236316 135215
rect 236288 128302 236500 128330
rect 236472 115977 236500 128302
rect 236274 115968 236330 115977
rect 236274 115903 236330 115912
rect 236458 115968 236514 115977
rect 236458 115903 236514 115912
rect 236288 109018 236316 115903
rect 236288 108990 236500 109018
rect 236472 106282 236500 108990
rect 236460 106276 236512 106282
rect 236460 106218 236512 106224
rect 236644 106276 236696 106282
rect 236644 106218 236696 106224
rect 236656 96665 236684 106218
rect 236274 96656 236330 96665
rect 236274 96591 236330 96600
rect 236642 96656 236698 96665
rect 236642 96591 236698 96600
rect 236288 89706 236316 96591
rect 236288 89678 236500 89706
rect 236472 77314 236500 89678
rect 236276 77308 236328 77314
rect 236276 77250 236328 77256
rect 236460 77308 236512 77314
rect 236460 77250 236512 77256
rect 236288 67590 236316 77250
rect 236276 67584 236328 67590
rect 236276 67526 236328 67532
rect 236276 57996 236328 58002
rect 236276 57938 236328 57944
rect 236288 48278 236316 57938
rect 236276 48272 236328 48278
rect 236276 48214 236328 48220
rect 236276 37324 236328 37330
rect 236276 37266 236328 37272
rect 236288 27606 236316 37266
rect 238758 29200 238814 29209
rect 238758 29135 238760 29144
rect 238812 29135 238814 29144
rect 238760 29106 238812 29112
rect 236276 27600 236328 27606
rect 236276 27542 236328 27548
rect 236276 18012 236328 18018
rect 236276 17954 236328 17960
rect 236184 9036 236236 9042
rect 236184 8978 236236 8984
rect 236092 5160 236144 5166
rect 236092 5102 236144 5108
rect 236288 3534 236316 17954
rect 238864 7750 238892 340054
rect 238956 340054 239338 340082
rect 239508 340054 239798 340082
rect 240258 340054 240364 340082
rect 238956 11762 238984 340054
rect 239508 331242 239536 340054
rect 239140 331214 239536 331242
rect 239140 321450 239168 331214
rect 239140 321422 239260 321450
rect 239232 311914 239260 321422
rect 239036 311908 239088 311914
rect 239036 311850 239088 311856
rect 239220 311908 239272 311914
rect 239220 311850 239272 311856
rect 239048 311794 239076 311850
rect 239048 311766 239168 311794
rect 239140 309126 239168 311766
rect 239128 309120 239180 309126
rect 239128 309062 239180 309068
rect 239220 299532 239272 299538
rect 239220 299474 239272 299480
rect 239232 292602 239260 299474
rect 239036 292596 239088 292602
rect 239036 292538 239088 292544
rect 239220 292596 239272 292602
rect 239220 292538 239272 292544
rect 239048 292482 239076 292538
rect 239048 292454 239168 292482
rect 239140 282946 239168 292454
rect 239128 282940 239180 282946
rect 239128 282882 239180 282888
rect 239220 282804 239272 282810
rect 239220 282746 239272 282752
rect 239232 273290 239260 282746
rect 239036 273284 239088 273290
rect 239036 273226 239088 273232
rect 239220 273284 239272 273290
rect 239220 273226 239272 273232
rect 239048 273170 239076 273226
rect 239048 273142 239168 273170
rect 239140 263634 239168 273142
rect 239128 263628 239180 263634
rect 239128 263570 239180 263576
rect 239220 263492 239272 263498
rect 239220 263434 239272 263440
rect 239232 253978 239260 263434
rect 239036 253972 239088 253978
rect 239036 253914 239088 253920
rect 239220 253972 239272 253978
rect 239220 253914 239272 253920
rect 239048 253858 239076 253914
rect 239048 253830 239168 253858
rect 239140 251190 239168 253830
rect 239128 251184 239180 251190
rect 239128 251126 239180 251132
rect 239220 251184 239272 251190
rect 239220 251126 239272 251132
rect 239232 246242 239260 251126
rect 239232 246214 239352 246242
rect 239324 240145 239352 246214
rect 239310 240136 239366 240145
rect 239310 240071 239366 240080
rect 239494 240136 239550 240145
rect 239494 240071 239550 240080
rect 239508 231554 239536 240071
rect 239324 231526 239536 231554
rect 239324 227338 239352 231526
rect 239324 227310 239444 227338
rect 239416 212634 239444 227310
rect 239128 212628 239180 212634
rect 239128 212570 239180 212576
rect 239404 212628 239456 212634
rect 239404 212570 239456 212576
rect 239140 212537 239168 212570
rect 239126 212528 239182 212537
rect 239126 212463 239182 212472
rect 239310 212528 239366 212537
rect 239310 212463 239366 212472
rect 239324 211138 239352 212463
rect 239036 211132 239088 211138
rect 239036 211074 239088 211080
rect 239312 211132 239364 211138
rect 239312 211074 239364 211080
rect 239048 201521 239076 211074
rect 239034 201512 239090 201521
rect 239034 201447 239090 201456
rect 239218 201512 239274 201521
rect 239218 201447 239274 201456
rect 239232 193254 239260 201447
rect 239128 193248 239180 193254
rect 239128 193190 239180 193196
rect 239220 193248 239272 193254
rect 239220 193190 239272 193196
rect 239140 191826 239168 193190
rect 239128 191820 239180 191826
rect 239128 191762 239180 191768
rect 239404 191820 239456 191826
rect 239404 191762 239456 191768
rect 239416 172650 239444 191762
rect 239128 172644 239180 172650
rect 239128 172586 239180 172592
rect 239404 172644 239456 172650
rect 239404 172586 239456 172592
rect 239140 164286 239168 172586
rect 239128 164280 239180 164286
rect 239128 164222 239180 164228
rect 239312 164144 239364 164150
rect 239312 164086 239364 164092
rect 239324 162790 239352 164086
rect 239036 162784 239088 162790
rect 239036 162726 239088 162732
rect 239312 162784 239364 162790
rect 239312 162726 239364 162732
rect 239048 147642 239076 162726
rect 239048 147614 239168 147642
rect 239140 138145 239168 147614
rect 239126 138136 239182 138145
rect 239126 138071 239182 138080
rect 239126 135280 239182 135289
rect 239126 135215 239128 135224
rect 239180 135215 239182 135224
rect 239312 135244 239364 135250
rect 239128 135186 239180 135192
rect 239312 135186 239364 135192
rect 239324 115977 239352 135186
rect 239126 115968 239182 115977
rect 239126 115903 239182 115912
rect 239310 115968 239366 115977
rect 239310 115903 239366 115912
rect 239140 106282 239168 115903
rect 239128 106276 239180 106282
rect 239128 106218 239180 106224
rect 239312 106276 239364 106282
rect 239312 106218 239364 106224
rect 239324 96665 239352 106218
rect 239126 96656 239182 96665
rect 239126 96591 239182 96600
rect 239310 96656 239366 96665
rect 239310 96591 239366 96600
rect 239140 60738 239168 96591
rect 239048 60710 239168 60738
rect 239048 60602 239076 60710
rect 239048 60574 239168 60602
rect 239140 41342 239168 60574
rect 239128 41336 239180 41342
rect 239128 41278 239180 41284
rect 239128 37324 239180 37330
rect 239128 37266 239180 37272
rect 238944 11756 238996 11762
rect 238944 11698 238996 11704
rect 239140 9738 239168 37266
rect 239048 9710 239168 9738
rect 238852 7744 238904 7750
rect 238852 7686 238904 7692
rect 238392 6996 238444 7002
rect 238392 6938 238444 6944
rect 237196 4956 237248 4962
rect 237196 4898 237248 4904
rect 236276 3528 236328 3534
rect 236276 3470 236328 3476
rect 237208 480 237236 4898
rect 238404 480 238432 6938
rect 239048 3670 239076 9710
rect 239588 9036 239640 9042
rect 239588 8978 239640 8984
rect 239036 3664 239088 3670
rect 239036 3606 239088 3612
rect 239600 480 239628 8978
rect 240336 3602 240364 340054
rect 240428 340054 240810 340082
rect 240428 7818 240456 340054
rect 241256 337414 241284 340068
rect 241716 337618 241744 340068
rect 241808 340054 242282 340082
rect 242360 340054 242742 340082
rect 243096 340054 243202 340082
rect 243464 340054 243754 340082
rect 241704 337612 241756 337618
rect 241704 337554 241756 337560
rect 241244 337408 241296 337414
rect 241244 337350 241296 337356
rect 241612 335640 241664 335646
rect 241612 335582 241664 335588
rect 241624 13122 241652 335582
rect 241612 13116 241664 13122
rect 241612 13058 241664 13064
rect 241808 7886 241836 340054
rect 242360 335646 242388 340054
rect 242348 335640 242400 335646
rect 242348 335582 242400 335588
rect 242992 332104 243044 332110
rect 242992 332046 243044 332052
rect 243004 7954 243032 332046
rect 242992 7948 243044 7954
rect 242992 7890 243044 7896
rect 241796 7880 241848 7886
rect 241796 7822 241848 7828
rect 240416 7812 240468 7818
rect 240416 7754 240468 7760
rect 241980 7744 242032 7750
rect 241980 7686 242032 7692
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 240324 3596 240376 3602
rect 240324 3538 240376 3544
rect 240796 480 240824 4966
rect 241992 480 242020 7686
rect 243096 3738 243124 340054
rect 243464 332110 243492 340054
rect 244200 337822 244228 340068
rect 244660 338706 244688 340068
rect 244648 338700 244700 338706
rect 244648 338642 244700 338648
rect 244188 337816 244240 337822
rect 244188 337758 244240 337764
rect 243452 332104 243504 332110
rect 243452 332046 243504 332052
rect 244752 331242 244780 340190
rect 244476 331214 244780 331242
rect 244476 321638 244504 331214
rect 244464 321632 244516 321638
rect 244464 321574 244516 321580
rect 244372 321564 244424 321570
rect 244372 321506 244424 321512
rect 244384 315994 244412 321506
rect 244372 315988 244424 315994
rect 244372 315930 244424 315936
rect 244556 315852 244608 315858
rect 244556 315794 244608 315800
rect 244568 270552 244596 315794
rect 244476 270524 244596 270552
rect 244476 267753 244504 270524
rect 244462 267744 244518 267753
rect 244462 267679 244518 267688
rect 244646 267744 244702 267753
rect 244646 267679 244702 267688
rect 244660 260658 244688 267679
rect 244476 260630 244688 260658
rect 244476 240174 244504 260630
rect 244372 240168 244424 240174
rect 244372 240110 244424 240116
rect 244464 240168 244516 240174
rect 244464 240110 244516 240116
rect 244384 234870 244412 240110
rect 244372 234864 244424 234870
rect 244372 234806 244424 234812
rect 244372 230512 244424 230518
rect 244372 230454 244424 230460
rect 244384 229090 244412 230454
rect 244280 229084 244332 229090
rect 244280 229026 244332 229032
rect 244372 229084 244424 229090
rect 244372 229026 244424 229032
rect 244292 219473 244320 229026
rect 244278 219464 244334 219473
rect 244554 219464 244610 219473
rect 244278 219399 244334 219408
rect 244464 219428 244516 219434
rect 244554 219399 244556 219408
rect 244464 219370 244516 219376
rect 244608 219399 244610 219408
rect 244556 219370 244608 219376
rect 244476 218006 244504 219370
rect 244464 218000 244516 218006
rect 244464 217942 244516 217948
rect 244464 200184 244516 200190
rect 244464 200126 244516 200132
rect 244476 186998 244504 200126
rect 244464 186992 244516 186998
rect 244464 186934 244516 186940
rect 244372 180872 244424 180878
rect 244372 180814 244424 180820
rect 244384 173942 244412 180814
rect 244372 173936 244424 173942
rect 244372 173878 244424 173884
rect 244464 173936 244516 173942
rect 244464 173878 244516 173884
rect 244476 169130 244504 173878
rect 244384 169102 244504 169130
rect 244384 164218 244412 169102
rect 244372 164212 244424 164218
rect 244372 164154 244424 164160
rect 244556 164212 244608 164218
rect 244556 164154 244608 164160
rect 244568 159202 244596 164154
rect 244476 159174 244596 159202
rect 244476 145081 244504 159174
rect 244462 145072 244518 145081
rect 244462 145007 244518 145016
rect 244462 144936 244518 144945
rect 244462 144871 244518 144880
rect 244476 143546 244504 144871
rect 244464 143540 244516 143546
rect 244464 143482 244516 143488
rect 244464 137964 244516 137970
rect 244464 137906 244516 137912
rect 244476 116090 244504 137906
rect 244384 116062 244504 116090
rect 244384 115954 244412 116062
rect 244384 115926 244504 115954
rect 244476 99482 244504 115926
rect 244464 99476 244516 99482
rect 244464 99418 244516 99424
rect 244464 99340 244516 99346
rect 244464 99282 244516 99288
rect 244476 60738 244504 99282
rect 244384 60710 244504 60738
rect 244384 60602 244412 60710
rect 244384 60574 244504 60602
rect 244476 51134 244504 60574
rect 245568 57928 245620 57934
rect 245568 57870 245620 57876
rect 244464 51128 244516 51134
rect 244464 51070 244516 51076
rect 244372 51060 244424 51066
rect 244372 51002 244424 51008
rect 244384 38758 244412 51002
rect 245580 48385 245608 57870
rect 245566 48376 245622 48385
rect 245566 48311 245622 48320
rect 245566 48240 245622 48249
rect 245566 48175 245622 48184
rect 244372 38752 244424 38758
rect 244372 38694 244424 38700
rect 245580 38690 245608 48175
rect 244464 38684 244516 38690
rect 244464 38626 244516 38632
rect 245568 38684 245620 38690
rect 245568 38626 245620 38632
rect 244476 37262 244504 38626
rect 244464 37256 244516 37262
rect 244464 37198 244516 37204
rect 244372 28076 244424 28082
rect 244372 28018 244424 28024
rect 244384 26246 244412 28018
rect 244372 26240 244424 26246
rect 244372 26182 244424 26188
rect 244188 16652 244240 16658
rect 244188 16594 244240 16600
rect 243176 9104 243228 9110
rect 243176 9046 243228 9052
rect 243084 3732 243136 3738
rect 243084 3674 243136 3680
rect 243188 480 243216 9046
rect 244200 8022 244228 16594
rect 244188 8016 244240 8022
rect 244188 7958 244240 7964
rect 245568 7812 245620 7818
rect 245568 7754 245620 7760
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 244384 480 244412 5034
rect 245580 480 245608 7754
rect 245672 3806 245700 340068
rect 245764 340054 246146 340082
rect 245764 3874 245792 340054
rect 246224 334642 246252 340190
rect 247144 337890 247172 340068
rect 247604 337958 247632 340068
rect 247592 337952 247644 337958
rect 247592 337894 247644 337900
rect 247132 337884 247184 337890
rect 247132 337826 247184 337832
rect 248156 336462 248184 340068
rect 247224 336456 247276 336462
rect 247224 336398 247276 336404
rect 248144 336456 248196 336462
rect 248144 336398 248196 336404
rect 245948 334614 246252 334642
rect 245948 325689 245976 334614
rect 245934 325680 245990 325689
rect 245934 325615 245990 325624
rect 246118 325680 246174 325689
rect 246118 325615 246174 325624
rect 246132 316062 246160 325615
rect 245844 316056 245896 316062
rect 245842 316024 245844 316033
rect 246120 316056 246172 316062
rect 245896 316024 245898 316033
rect 246120 315998 246172 316004
rect 245842 315959 245898 315968
rect 245934 315888 245990 315897
rect 245934 315823 245990 315832
rect 245948 302462 245976 315823
rect 245936 302456 245988 302462
rect 245936 302398 245988 302404
rect 246028 298036 246080 298042
rect 246028 297978 246080 297984
rect 246040 270552 246068 297978
rect 245948 270524 246068 270552
rect 245948 267753 245976 270524
rect 245934 267744 245990 267753
rect 245934 267679 245990 267688
rect 246118 267744 246174 267753
rect 246118 267679 246174 267688
rect 246132 258097 246160 267679
rect 245842 258088 245898 258097
rect 245842 258023 245898 258032
rect 246118 258088 246174 258097
rect 246118 258023 246174 258032
rect 245856 257990 245884 258023
rect 245844 257984 245896 257990
rect 245844 257926 245896 257932
rect 245936 257984 245988 257990
rect 245936 257926 245988 257932
rect 245948 240174 245976 257926
rect 245844 240168 245896 240174
rect 245842 240136 245844 240145
rect 245936 240168 245988 240174
rect 245896 240136 245898 240145
rect 245936 240110 245988 240116
rect 246118 240136 246174 240145
rect 245842 240071 245898 240080
rect 246118 240071 246174 240080
rect 246132 230518 246160 240071
rect 245936 230512 245988 230518
rect 245936 230454 245988 230460
rect 246120 230512 246172 230518
rect 246120 230454 246172 230460
rect 245948 227202 245976 230454
rect 245948 227174 246068 227202
rect 246040 222222 246068 227174
rect 245844 222216 245896 222222
rect 245844 222158 245896 222164
rect 246028 222216 246080 222222
rect 246028 222158 246080 222164
rect 245856 212566 245884 222158
rect 245844 212560 245896 212566
rect 245844 212502 245896 212508
rect 245936 212560 245988 212566
rect 245936 212502 245988 212508
rect 245948 202910 245976 212502
rect 245844 202904 245896 202910
rect 245844 202846 245896 202852
rect 245936 202904 245988 202910
rect 245936 202846 245988 202852
rect 245856 193390 245884 202846
rect 245844 193384 245896 193390
rect 245844 193326 245896 193332
rect 245844 193180 245896 193186
rect 245844 193122 245896 193128
rect 245856 173942 245884 193122
rect 245844 173936 245896 173942
rect 245844 173878 245896 173884
rect 245936 173936 245988 173942
rect 245936 173878 245988 173884
rect 245948 164257 245976 173878
rect 245934 164248 245990 164257
rect 245934 164183 245990 164192
rect 245842 164112 245898 164121
rect 245842 164047 245898 164056
rect 245856 162858 245884 164047
rect 245844 162852 245896 162858
rect 245844 162794 245896 162800
rect 245936 154488 245988 154494
rect 245936 154430 245988 154436
rect 245948 153202 245976 154430
rect 245936 153196 245988 153202
rect 245936 153138 245988 153144
rect 245936 143608 245988 143614
rect 245936 143550 245988 143556
rect 245948 143426 245976 143550
rect 245856 143398 245976 143426
rect 245856 133929 245884 143398
rect 245842 133920 245898 133929
rect 245842 133855 245898 133864
rect 246118 133920 246174 133929
rect 246118 133855 246174 133864
rect 246132 125633 246160 133855
rect 245934 125624 245990 125633
rect 245934 125559 245990 125568
rect 246118 125624 246174 125633
rect 246118 125559 246174 125568
rect 245948 99482 245976 125559
rect 245936 99476 245988 99482
rect 245936 99418 245988 99424
rect 245936 99340 245988 99346
rect 245936 99282 245988 99288
rect 245948 60738 245976 99282
rect 245856 60710 245976 60738
rect 245856 60602 245884 60710
rect 245856 60574 245976 60602
rect 245948 57934 245976 60574
rect 245936 57928 245988 57934
rect 245936 57870 245988 57876
rect 245936 38684 245988 38690
rect 245936 38626 245988 38632
rect 245948 37262 245976 38626
rect 245936 37256 245988 37262
rect 245936 37198 245988 37204
rect 245844 27668 245896 27674
rect 245844 27610 245896 27616
rect 245856 26246 245884 27610
rect 245844 26240 245896 26246
rect 245844 26182 245896 26188
rect 246028 16652 246080 16658
rect 246028 16594 246080 16600
rect 246040 13122 246068 16594
rect 245844 13116 245896 13122
rect 245844 13058 245896 13064
rect 246028 13116 246080 13122
rect 246028 13058 246080 13064
rect 245856 8242 245884 13058
rect 247236 9178 247264 336398
rect 248512 334960 248564 334966
rect 248512 334902 248564 334908
rect 247868 334008 247920 334014
rect 247868 333950 247920 333956
rect 247880 331242 247908 333950
rect 247696 331214 247908 331242
rect 247224 9172 247276 9178
rect 247224 9114 247276 9120
rect 246764 8356 246816 8362
rect 246764 8298 246816 8304
rect 245856 8214 245976 8242
rect 245948 8090 245976 8214
rect 245936 8084 245988 8090
rect 245936 8026 245988 8032
rect 245752 3868 245804 3874
rect 245752 3810 245804 3816
rect 245660 3800 245712 3806
rect 245660 3742 245712 3748
rect 246776 480 246804 8298
rect 247696 3942 247724 331214
rect 248524 5234 248552 334902
rect 248616 334014 248644 340068
rect 248708 340054 249090 340082
rect 248604 334008 248656 334014
rect 248604 333950 248656 333956
rect 248512 5228 248564 5234
rect 248512 5170 248564 5176
rect 247960 5160 248012 5166
rect 247960 5102 248012 5108
rect 247684 3936 247736 3942
rect 247684 3878 247736 3884
rect 247972 480 248000 5102
rect 248708 4010 248736 340054
rect 249064 336728 249116 336734
rect 249064 336670 249116 336676
rect 249246 336696 249302 336705
rect 249076 4078 249104 336670
rect 249246 336631 249302 336640
rect 249260 316305 249288 336631
rect 249536 334966 249564 340068
rect 249904 340054 250102 340082
rect 249524 334960 249576 334966
rect 249524 334902 249576 334908
rect 249246 316296 249302 316305
rect 249246 316231 249302 316240
rect 249246 306368 249302 306377
rect 249246 306303 249302 306312
rect 249260 296993 249288 306303
rect 249246 296984 249302 296993
rect 249246 296919 249302 296928
rect 249430 275088 249486 275097
rect 249430 275023 249486 275032
rect 249444 267889 249472 275023
rect 249430 267880 249486 267889
rect 249430 267815 249486 267824
rect 249246 257952 249302 257961
rect 249246 257887 249302 257896
rect 249260 248441 249288 257887
rect 249246 248432 249302 248441
rect 249246 248367 249302 248376
rect 249614 209672 249670 209681
rect 249614 209607 249670 209616
rect 249628 200161 249656 209607
rect 249614 200152 249670 200161
rect 249614 200087 249670 200096
rect 249338 193216 249394 193225
rect 249338 193151 249394 193160
rect 249352 182209 249380 193151
rect 249338 182200 249394 182209
rect 249338 182135 249394 182144
rect 249904 9246 249932 340054
rect 250444 337408 250496 337414
rect 250444 337350 250496 337356
rect 250168 327140 250220 327146
rect 250168 327082 250220 327088
rect 250180 317422 250208 327082
rect 250168 317416 250220 317422
rect 250168 317358 250220 317364
rect 250168 307828 250220 307834
rect 250168 307770 250220 307776
rect 250180 298110 250208 307770
rect 250168 298104 250220 298110
rect 250168 298046 250220 298052
rect 250168 289808 250220 289814
rect 250168 289750 250220 289756
rect 250180 280158 250208 289750
rect 250076 280152 250128 280158
rect 250076 280094 250128 280100
rect 250168 280152 250220 280158
rect 250168 280094 250220 280100
rect 250088 278769 250116 280094
rect 250074 278760 250130 278769
rect 250074 278695 250130 278704
rect 250258 278760 250314 278769
rect 250258 278695 250314 278704
rect 250272 269142 250300 278695
rect 250076 269136 250128 269142
rect 250076 269078 250128 269084
rect 250260 269136 250312 269142
rect 250260 269078 250312 269084
rect 250088 260914 250116 269078
rect 250076 260908 250128 260914
rect 250076 260850 250128 260856
rect 250168 260908 250220 260914
rect 250168 260850 250220 260856
rect 250180 259434 250208 260850
rect 250088 259406 250208 259434
rect 250088 253978 250116 259406
rect 250076 253972 250128 253978
rect 250076 253914 250128 253920
rect 250076 249824 250128 249830
rect 250076 249766 250128 249772
rect 250088 241534 250116 249766
rect 250076 241528 250128 241534
rect 250076 241470 250128 241476
rect 250168 241528 250220 241534
rect 250168 241470 250220 241476
rect 250180 240122 250208 241470
rect 250088 240094 250208 240122
rect 250088 234666 250116 240094
rect 250076 234660 250128 234666
rect 250076 234602 250128 234608
rect 250168 230512 250220 230518
rect 250168 230454 250220 230460
rect 250180 217410 250208 230454
rect 250180 217382 250300 217410
rect 250272 212566 250300 217382
rect 250076 212560 250128 212566
rect 250076 212502 250128 212508
rect 250260 212560 250312 212566
rect 250260 212502 250312 212508
rect 250088 205698 250116 212502
rect 250076 205692 250128 205698
rect 250076 205634 250128 205640
rect 250168 205624 250220 205630
rect 250168 205566 250220 205572
rect 250180 198098 250208 205566
rect 250180 198070 250300 198098
rect 250272 193254 250300 198070
rect 250076 193248 250128 193254
rect 250074 193216 250076 193225
rect 250260 193248 250312 193254
rect 250128 193216 250130 193225
rect 250074 193151 250130 193160
rect 250258 193216 250260 193225
rect 250312 193216 250314 193225
rect 250258 193151 250314 193160
rect 250272 186266 250300 193151
rect 250180 186238 250300 186266
rect 250180 178786 250208 186238
rect 250180 178758 250300 178786
rect 250272 173942 250300 178758
rect 250076 173936 250128 173942
rect 250076 173878 250128 173884
rect 250260 173936 250312 173942
rect 250260 173878 250312 173884
rect 250088 162858 250116 173878
rect 250076 162852 250128 162858
rect 250076 162794 250128 162800
rect 250352 162784 250404 162790
rect 250352 162726 250404 162732
rect 250364 161430 250392 162726
rect 250352 161424 250404 161430
rect 250352 161366 250404 161372
rect 250352 151836 250404 151842
rect 250352 151778 250404 151784
rect 250364 144974 250392 151778
rect 250352 144968 250404 144974
rect 250352 144910 250404 144916
rect 250168 144900 250220 144906
rect 250168 144842 250220 144848
rect 250180 143546 250208 144842
rect 250168 143540 250220 143546
rect 250168 143482 250220 143488
rect 250260 143540 250312 143546
rect 250260 143482 250312 143488
rect 250272 142118 250300 143482
rect 250260 142112 250312 142118
rect 250260 142054 250312 142060
rect 249984 132524 250036 132530
rect 249984 132466 250036 132472
rect 249996 124166 250024 132466
rect 249984 124160 250036 124166
rect 249984 124102 250036 124108
rect 250260 114572 250312 114578
rect 250260 114514 250312 114520
rect 250272 96694 250300 114514
rect 250076 96688 250128 96694
rect 250076 96630 250128 96636
rect 250260 96688 250312 96694
rect 250260 96630 250312 96636
rect 250088 77450 250116 96630
rect 250076 77444 250128 77450
rect 250076 77386 250128 77392
rect 249984 77308 250036 77314
rect 249984 77250 250036 77256
rect 249996 67674 250024 77250
rect 249996 67646 250116 67674
rect 250088 66230 250116 67646
rect 250076 66224 250128 66230
rect 250076 66166 250128 66172
rect 250076 60716 250128 60722
rect 250076 60658 250128 60664
rect 250088 50998 250116 60658
rect 250076 50992 250128 50998
rect 250076 50934 250128 50940
rect 250076 48340 250128 48346
rect 250076 48282 250128 48288
rect 250088 31770 250116 48282
rect 250088 31742 250300 31770
rect 250272 31634 250300 31742
rect 250180 31606 250300 31634
rect 250180 26246 250208 31606
rect 249984 26240 250036 26246
rect 249984 26182 250036 26188
rect 250168 26240 250220 26246
rect 250168 26182 250220 26188
rect 249892 9240 249944 9246
rect 249892 9182 249944 9188
rect 249156 7880 249208 7886
rect 249156 7822 249208 7828
rect 249064 4072 249116 4078
rect 249064 4014 249116 4020
rect 248696 4004 248748 4010
rect 248696 3946 248748 3952
rect 249168 480 249196 7822
rect 249996 6225 250024 26182
rect 250352 9172 250404 9178
rect 250352 9114 250404 9120
rect 249982 6216 250038 6225
rect 249982 6151 250038 6160
rect 250364 480 250392 9114
rect 250456 4146 250484 337350
rect 250548 336734 250576 340068
rect 250640 340054 251022 340082
rect 251284 340054 251574 340082
rect 250536 336728 250588 336734
rect 250536 336670 250588 336676
rect 250640 334490 250668 340054
rect 250628 334484 250680 334490
rect 250628 334426 250680 334432
rect 251178 280120 251234 280129
rect 251178 280055 251234 280064
rect 251192 270570 251220 280055
rect 251180 270564 251232 270570
rect 251180 270506 251232 270512
rect 251178 260808 251234 260817
rect 251178 260743 251234 260752
rect 251192 259078 251220 260743
rect 251180 259072 251232 259078
rect 251180 259014 251232 259020
rect 251086 240136 251142 240145
rect 251086 240071 251142 240080
rect 251100 230518 251128 240071
rect 251088 230512 251140 230518
rect 251088 230454 251140 230460
rect 251180 180804 251232 180810
rect 251180 180746 251232 180752
rect 251192 162897 251220 180746
rect 251178 162888 251234 162897
rect 251178 162823 251234 162832
rect 251086 87544 251142 87553
rect 251086 87479 251142 87488
rect 251100 87281 251128 87479
rect 251086 87272 251142 87281
rect 251086 87207 251142 87216
rect 251178 87136 251234 87145
rect 251178 87071 251180 87080
rect 251232 87071 251234 87080
rect 251180 87042 251232 87048
rect 251086 76120 251142 76129
rect 251086 76055 251142 76064
rect 251100 75721 251128 76055
rect 251086 75712 251142 75721
rect 251086 75647 251142 75656
rect 251284 10334 251312 340054
rect 252020 338026 252048 340068
rect 252008 338020 252060 338026
rect 252008 337962 252060 337968
rect 251824 336728 251876 336734
rect 251824 336670 251876 336676
rect 251456 335844 251508 335850
rect 251456 335786 251508 335792
rect 251468 323626 251496 335786
rect 251468 323598 251588 323626
rect 251560 317422 251588 323598
rect 251548 317416 251600 317422
rect 251548 317358 251600 317364
rect 251548 307828 251600 307834
rect 251548 307770 251600 307776
rect 251560 307737 251588 307770
rect 251546 307728 251602 307737
rect 251546 307663 251602 307672
rect 251546 298208 251602 298217
rect 251546 298143 251602 298152
rect 251560 298110 251588 298143
rect 251548 298104 251600 298110
rect 251548 298046 251600 298052
rect 251364 288448 251416 288454
rect 251364 288390 251416 288396
rect 251376 280129 251404 288390
rect 251362 280120 251418 280129
rect 251362 280055 251418 280064
rect 251456 270564 251508 270570
rect 251456 270506 251508 270512
rect 251468 265690 251496 270506
rect 251468 265662 251588 265690
rect 251560 263514 251588 265662
rect 251376 263486 251588 263514
rect 251376 260817 251404 263486
rect 251362 260808 251418 260817
rect 251362 260743 251418 260752
rect 251364 259072 251416 259078
rect 251364 259014 251416 259020
rect 251376 241534 251404 259014
rect 251364 241528 251416 241534
rect 251364 241470 251416 241476
rect 251364 240168 251416 240174
rect 251362 240136 251364 240145
rect 251416 240136 251418 240145
rect 251362 240071 251418 240080
rect 251364 230512 251416 230518
rect 251362 230480 251364 230489
rect 251416 230480 251418 230489
rect 251362 230415 251418 230424
rect 251546 230480 251602 230489
rect 251546 230415 251602 230424
rect 251560 220862 251588 230415
rect 251548 220856 251600 220862
rect 251548 220798 251600 220804
rect 251640 220856 251692 220862
rect 251640 220798 251692 220804
rect 251652 212514 251680 220798
rect 251560 212486 251680 212514
rect 251560 205578 251588 212486
rect 251468 205550 251588 205578
rect 251468 202722 251496 205550
rect 251468 202694 251588 202722
rect 251560 191826 251588 202694
rect 251548 191820 251600 191826
rect 251548 191762 251600 191768
rect 251640 191820 251692 191826
rect 251640 191762 251692 191768
rect 251652 182186 251680 191762
rect 251652 182170 251772 182186
rect 251456 182164 251508 182170
rect 251652 182164 251784 182170
rect 251652 182158 251732 182164
rect 251456 182106 251508 182112
rect 251732 182106 251784 182112
rect 251468 180810 251496 182106
rect 251456 180804 251508 180810
rect 251456 180746 251508 180752
rect 251362 162888 251418 162897
rect 251362 162823 251418 162832
rect 251376 157162 251404 162823
rect 251376 157134 251680 157162
rect 251652 143585 251680 157134
rect 251454 143576 251510 143585
rect 251454 143511 251510 143520
rect 251638 143576 251694 143585
rect 251638 143511 251694 143520
rect 251468 138038 251496 143511
rect 251456 138032 251508 138038
rect 251456 137974 251508 137980
rect 251456 133952 251508 133958
rect 251456 133894 251508 133900
rect 251468 118794 251496 133894
rect 251456 118788 251508 118794
rect 251456 118730 251508 118736
rect 251456 118652 251508 118658
rect 251456 118594 251508 118600
rect 251468 99414 251496 118594
rect 251456 99408 251508 99414
rect 251456 99350 251508 99356
rect 251456 96688 251508 96694
rect 251456 96630 251508 96636
rect 251468 86970 251496 96630
rect 251456 86964 251508 86970
rect 251456 86906 251508 86912
rect 251456 77308 251508 77314
rect 251456 77250 251508 77256
rect 251468 60738 251496 77250
rect 251376 60710 251496 60738
rect 251376 60602 251404 60710
rect 251376 60574 251496 60602
rect 251468 48521 251496 60574
rect 251454 48512 251510 48521
rect 251454 48447 251510 48456
rect 251362 48376 251418 48385
rect 251362 48311 251418 48320
rect 251376 44146 251404 48311
rect 251376 44118 251496 44146
rect 251468 41478 251496 44118
rect 251456 41472 251508 41478
rect 251456 41414 251508 41420
rect 251364 41404 251416 41410
rect 251364 41346 251416 41352
rect 251376 26353 251404 41346
rect 251362 26344 251418 26353
rect 251362 26279 251418 26288
rect 251638 26208 251694 26217
rect 251638 26143 251694 26152
rect 251652 21434 251680 26143
rect 251376 21406 251680 21434
rect 251272 10328 251324 10334
rect 251272 10270 251324 10276
rect 251376 6186 251404 21406
rect 251364 6180 251416 6186
rect 251364 6122 251416 6128
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 250444 4140 250496 4146
rect 250444 4082 250496 4088
rect 251468 480 251496 5170
rect 251836 3398 251864 336670
rect 252480 335850 252508 340068
rect 252664 340054 253046 340082
rect 252468 335844 252520 335850
rect 252468 335786 252520 335792
rect 252664 10402 252692 340054
rect 253204 337544 253256 337550
rect 253204 337486 253256 337492
rect 252652 10396 252704 10402
rect 252652 10338 252704 10344
rect 252652 7948 252704 7954
rect 252652 7890 252704 7896
rect 251824 3392 251876 3398
rect 251824 3334 251876 3340
rect 252664 480 252692 7890
rect 253216 3330 253244 337486
rect 253492 337414 253520 340068
rect 253480 337408 253532 337414
rect 253480 337350 253532 337356
rect 253848 9240 253900 9246
rect 253848 9182 253900 9188
rect 253204 3324 253256 3330
rect 253204 3266 253256 3272
rect 253860 480 253888 9182
rect 253952 6254 253980 340068
rect 254044 340054 254518 340082
rect 254044 10470 254072 340054
rect 254964 338094 254992 340068
rect 255438 340054 255544 340082
rect 254952 338088 255004 338094
rect 254952 338030 255004 338036
rect 254584 337748 254636 337754
rect 254584 337690 254636 337696
rect 254032 10464 254084 10470
rect 254032 10406 254084 10412
rect 253940 6248 253992 6254
rect 253940 6190 253992 6196
rect 254596 3262 254624 337690
rect 255516 6322 255544 340054
rect 255608 340054 255990 340082
rect 255608 10538 255636 340054
rect 255964 337680 256016 337686
rect 255964 337622 256016 337628
rect 255596 10532 255648 10538
rect 255596 10474 255648 10480
rect 255504 6316 255556 6322
rect 255504 6258 255556 6264
rect 255044 3460 255096 3466
rect 255044 3402 255096 3408
rect 254584 3256 254636 3262
rect 254584 3198 254636 3204
rect 255056 480 255084 3402
rect 255976 3194 256004 337622
rect 256436 336734 256464 340068
rect 256804 340054 256910 340082
rect 256988 340054 257462 340082
rect 256424 336728 256476 336734
rect 256424 336670 256476 336676
rect 256608 29164 256660 29170
rect 256608 29106 256660 29112
rect 256620 29073 256648 29106
rect 256606 29064 256662 29073
rect 256606 28999 256662 29008
rect 256240 8016 256292 8022
rect 256240 7958 256292 7964
rect 255964 3188 256016 3194
rect 255964 3130 256016 3136
rect 256252 480 256280 7958
rect 256804 6390 256832 340054
rect 256792 6384 256844 6390
rect 256792 6326 256844 6332
rect 256988 5302 257016 340054
rect 257344 337408 257396 337414
rect 257344 337350 257396 337356
rect 256976 5296 257028 5302
rect 256976 5238 257028 5244
rect 257356 3126 257384 337350
rect 257908 337278 257936 340068
rect 258276 340054 258382 340082
rect 258552 340054 258934 340082
rect 257896 337272 257948 337278
rect 257896 337214 257948 337220
rect 258172 334620 258224 334626
rect 258172 334562 258224 334568
rect 257986 29336 258042 29345
rect 257986 29271 258042 29280
rect 258000 29073 258028 29271
rect 257986 29064 258042 29073
rect 257986 28999 258042 29008
rect 258184 13190 258212 334562
rect 258172 13184 258224 13190
rect 258172 13126 258224 13132
rect 258276 6458 258304 340054
rect 258552 334626 258580 340054
rect 259380 337550 259408 340068
rect 259472 340054 259854 340082
rect 260116 340054 260406 340082
rect 259368 337544 259420 337550
rect 259368 337486 259420 337492
rect 258816 337476 258868 337482
rect 258816 337418 258868 337424
rect 258724 337272 258776 337278
rect 258724 337214 258776 337220
rect 258540 334620 258592 334626
rect 258540 334562 258592 334568
rect 258264 6452 258316 6458
rect 258264 6394 258316 6400
rect 257436 4004 257488 4010
rect 257436 3946 257488 3952
rect 257344 3120 257396 3126
rect 257344 3062 257396 3068
rect 257448 480 257476 3946
rect 258632 3528 258684 3534
rect 258632 3470 258684 3476
rect 258644 480 258672 3470
rect 258736 3058 258764 337214
rect 258724 3052 258776 3058
rect 258724 2994 258776 3000
rect 258828 2990 258856 337418
rect 259366 64016 259422 64025
rect 259366 63951 259422 63960
rect 259380 63617 259408 63951
rect 259366 63608 259422 63617
rect 259366 63543 259422 63552
rect 259472 6526 259500 340054
rect 260116 337822 260144 340054
rect 259644 337816 259696 337822
rect 259644 337758 259696 337764
rect 260104 337816 260156 337822
rect 260104 337758 260156 337764
rect 259656 331226 259684 337758
rect 260104 337680 260156 337686
rect 260104 337622 260156 337628
rect 259644 331220 259696 331226
rect 259644 331162 259696 331168
rect 259828 331220 259880 331226
rect 259828 331162 259880 331168
rect 259840 328438 259868 331162
rect 259828 328432 259880 328438
rect 259828 328374 259880 328380
rect 259920 318844 259972 318850
rect 259920 318786 259972 318792
rect 259932 307834 259960 318786
rect 259736 307828 259788 307834
rect 259736 307770 259788 307776
rect 259920 307828 259972 307834
rect 259920 307770 259972 307776
rect 259748 306377 259776 307770
rect 259734 306368 259790 306377
rect 259734 306303 259790 306312
rect 259918 306368 259974 306377
rect 259918 306303 259974 306312
rect 259932 295361 259960 306303
rect 259642 295352 259698 295361
rect 259642 295287 259698 295296
rect 259918 295352 259974 295361
rect 259918 295287 259974 295296
rect 259656 292618 259684 295287
rect 259564 292590 259684 292618
rect 259564 285666 259592 292590
rect 259552 285660 259604 285666
rect 259552 285602 259604 285608
rect 259920 285660 259972 285666
rect 259920 285602 259972 285608
rect 259932 258097 259960 285602
rect 259734 258088 259790 258097
rect 259734 258023 259790 258032
rect 259918 258088 259974 258097
rect 259918 258023 259974 258032
rect 259748 251190 259776 258023
rect 259736 251184 259788 251190
rect 259736 251126 259788 251132
rect 259644 242684 259696 242690
rect 259644 242626 259696 242632
rect 259656 240145 259684 242626
rect 259642 240136 259698 240145
rect 259642 240071 259698 240080
rect 259826 240136 259882 240145
rect 259826 240071 259882 240080
rect 259840 230518 259868 240071
rect 259552 230512 259604 230518
rect 259552 230454 259604 230460
rect 259828 230512 259880 230518
rect 259828 230454 259880 230460
rect 259564 227066 259592 230454
rect 259564 227038 259684 227066
rect 259656 222193 259684 227038
rect 259642 222184 259698 222193
rect 259642 222119 259698 222128
rect 259734 221912 259790 221921
rect 259734 221847 259790 221856
rect 259748 205578 259776 221847
rect 259656 205550 259776 205578
rect 259656 202881 259684 205550
rect 259642 202872 259698 202881
rect 259642 202807 259698 202816
rect 259918 202872 259974 202881
rect 259918 202807 259974 202816
rect 259932 193254 259960 202807
rect 259736 193248 259788 193254
rect 259736 193190 259788 193196
rect 259920 193248 259972 193254
rect 259920 193190 259972 193196
rect 259748 186266 259776 193190
rect 259656 186238 259776 186266
rect 259656 173942 259684 186238
rect 259644 173936 259696 173942
rect 259644 173878 259696 173884
rect 259644 172576 259696 172582
rect 259644 172518 259696 172524
rect 259656 161498 259684 172518
rect 259552 161492 259604 161498
rect 259552 161434 259604 161440
rect 259644 161492 259696 161498
rect 259644 161434 259696 161440
rect 259564 143562 259592 161434
rect 259564 143534 259684 143562
rect 259656 142118 259684 143534
rect 259644 142112 259696 142118
rect 259644 142054 259696 142060
rect 259736 132524 259788 132530
rect 259736 132466 259788 132472
rect 259748 113218 259776 132466
rect 259644 113212 259696 113218
rect 259644 113154 259696 113160
rect 259736 113212 259788 113218
rect 259736 113154 259788 113160
rect 259656 109018 259684 113154
rect 259656 108990 259868 109018
rect 259840 106282 259868 108990
rect 259552 106276 259604 106282
rect 259552 106218 259604 106224
rect 259828 106276 259880 106282
rect 259828 106218 259880 106224
rect 259564 96665 259592 106218
rect 259550 96656 259606 96665
rect 259550 96591 259606 96600
rect 259734 96656 259790 96665
rect 259734 96591 259790 96600
rect 259748 91746 259776 96591
rect 259748 91718 259868 91746
rect 259840 86986 259868 91718
rect 259840 86958 259960 86986
rect 259932 77738 259960 86958
rect 259748 77710 259960 77738
rect 259748 60738 259776 77710
rect 259656 60722 259776 60738
rect 259644 60716 259776 60722
rect 259696 60710 259776 60716
rect 259828 60716 259880 60722
rect 259644 60658 259696 60664
rect 259828 60658 259880 60664
rect 259840 47002 259868 60658
rect 259656 46974 259868 47002
rect 259656 46918 259684 46974
rect 259644 46912 259696 46918
rect 259644 46854 259696 46860
rect 259736 46912 259788 46918
rect 259736 46854 259788 46860
rect 259748 22114 259776 46854
rect 259656 22086 259776 22114
rect 259656 14482 259684 22086
rect 259644 14476 259696 14482
rect 259644 14418 259696 14424
rect 259828 8084 259880 8090
rect 259828 8026 259880 8032
rect 259460 6520 259512 6526
rect 259460 6462 259512 6468
rect 258816 2984 258868 2990
rect 258816 2926 258868 2932
rect 259840 480 259868 8026
rect 260116 2922 260144 337622
rect 260852 337346 260880 340068
rect 261036 340054 261326 340082
rect 261496 340054 261878 340082
rect 260840 337340 260892 337346
rect 260840 337282 260892 337288
rect 260932 335640 260984 335646
rect 260932 335582 260984 335588
rect 260654 87136 260710 87145
rect 260654 87071 260656 87080
rect 260708 87071 260710 87080
rect 260656 87042 260708 87048
rect 260944 14550 260972 335582
rect 260932 14544 260984 14550
rect 260932 14486 260984 14492
rect 261036 6594 261064 340054
rect 261392 337612 261444 337618
rect 261392 337554 261444 337560
rect 261404 334370 261432 337554
rect 261496 335646 261524 340054
rect 262324 337754 262352 340068
rect 262416 340054 262798 340082
rect 263060 340054 263350 340082
rect 262312 337748 262364 337754
rect 262312 337690 262364 337696
rect 261484 335640 261536 335646
rect 261484 335582 261536 335588
rect 261404 334342 261524 334370
rect 261024 6588 261076 6594
rect 261024 6530 261076 6536
rect 260104 2916 260156 2922
rect 260104 2858 260156 2864
rect 261496 2854 261524 334342
rect 262416 8158 262444 340054
rect 263060 336734 263088 340054
rect 263796 337210 263824 340068
rect 263888 340054 264270 340082
rect 264440 340054 264822 340082
rect 263784 337204 263836 337210
rect 263784 337146 263836 337152
rect 262864 336728 262916 336734
rect 262864 336670 262916 336676
rect 263048 336728 263100 336734
rect 263048 336670 263100 336676
rect 262876 325718 262904 336670
rect 263692 335640 263744 335646
rect 263692 335582 263744 335588
rect 262680 325712 262732 325718
rect 262680 325654 262732 325660
rect 262864 325712 262916 325718
rect 262864 325654 262916 325660
rect 262692 298178 262720 325654
rect 262496 298172 262548 298178
rect 262496 298114 262548 298120
rect 262680 298172 262732 298178
rect 262680 298114 262732 298120
rect 262508 289882 262536 298114
rect 262496 289876 262548 289882
rect 262496 289818 262548 289824
rect 262680 289876 262732 289882
rect 262680 289818 262732 289824
rect 262692 283642 262720 289818
rect 262600 283614 262720 283642
rect 262600 269142 262628 283614
rect 262588 269136 262640 269142
rect 262588 269078 262640 269084
rect 262680 269136 262732 269142
rect 262680 269078 262732 269084
rect 262692 251190 262720 269078
rect 262680 251184 262732 251190
rect 262680 251126 262732 251132
rect 262772 251184 262824 251190
rect 262772 251126 262824 251132
rect 262784 231878 262812 251126
rect 262680 231872 262732 231878
rect 262680 231814 262732 231820
rect 262772 231872 262824 231878
rect 262772 231814 262824 231820
rect 262692 212514 262720 231814
rect 262600 212486 262720 212514
rect 262600 196042 262628 212486
rect 262588 196036 262640 196042
rect 262588 195978 262640 195984
rect 262680 195968 262732 195974
rect 262680 195910 262732 195916
rect 262692 186266 262720 195910
rect 262600 186238 262720 186266
rect 262600 173942 262628 186238
rect 262588 173936 262640 173942
rect 262588 173878 262640 173884
rect 262680 173936 262732 173942
rect 262680 173878 262732 173884
rect 262692 164234 262720 173878
rect 262600 164206 262720 164234
rect 262600 157434 262628 164206
rect 262508 157406 262628 157434
rect 262508 153218 262536 157406
rect 262508 153190 262628 153218
rect 262600 144906 262628 153190
rect 262588 144900 262640 144906
rect 262588 144842 262640 144848
rect 262772 144900 262824 144906
rect 262772 144842 262824 144848
rect 262784 139890 262812 144842
rect 262692 139862 262812 139890
rect 262692 128466 262720 139862
rect 262600 128438 262720 128466
rect 262600 128330 262628 128438
rect 262600 128302 262720 128330
rect 262692 120714 262720 128302
rect 262600 120686 262720 120714
rect 262600 109018 262628 120686
rect 262600 108990 262812 109018
rect 262784 101402 262812 108990
rect 262600 101374 262812 101402
rect 262600 99226 262628 101374
rect 262600 99198 262720 99226
rect 262692 87038 262720 99198
rect 262588 87032 262640 87038
rect 262588 86974 262640 86980
rect 262680 87032 262732 87038
rect 262680 86974 262732 86980
rect 262600 77314 262628 86974
rect 262588 77308 262640 77314
rect 262588 77250 262640 77256
rect 262680 77308 262732 77314
rect 262680 77250 262732 77256
rect 262692 60738 262720 77250
rect 262600 60722 262720 60738
rect 262588 60716 262720 60722
rect 262640 60710 262720 60716
rect 262772 60716 262824 60722
rect 262588 60658 262640 60664
rect 262772 60658 262824 60664
rect 262784 52290 262812 60658
rect 262588 52284 262640 52290
rect 262588 52226 262640 52232
rect 262772 52284 262824 52290
rect 262772 52226 262824 52232
rect 262600 41154 262628 52226
rect 262600 41126 262720 41154
rect 262692 22114 262720 41126
rect 263414 29336 263470 29345
rect 263598 29336 263654 29345
rect 263470 29294 263598 29322
rect 263414 29271 263470 29280
rect 263598 29271 263654 29280
rect 262600 22086 262720 22114
rect 262600 14618 262628 22086
rect 263704 14686 263732 335582
rect 263692 14680 263744 14686
rect 263692 14622 263744 14628
rect 262588 14612 262640 14618
rect 262588 14554 262640 14560
rect 263888 8226 263916 340054
rect 264440 335646 264468 340054
rect 265268 337074 265296 340068
rect 265452 340054 265742 340082
rect 265912 340054 266294 340082
rect 265256 337068 265308 337074
rect 265256 337010 265308 337016
rect 264428 335640 264480 335646
rect 264428 335582 264480 335588
rect 265072 335640 265124 335646
rect 265452 335594 265480 340054
rect 265912 335646 265940 340054
rect 266740 337414 266768 340068
rect 266924 340054 267214 340082
rect 267384 340054 267674 340082
rect 266728 337408 266780 337414
rect 266728 337350 266780 337356
rect 265072 335582 265124 335588
rect 264978 314664 265034 314673
rect 264978 314599 265034 314608
rect 264992 305017 265020 314599
rect 264978 305008 265034 305017
rect 264978 304943 265034 304952
rect 264980 262948 265032 262954
rect 264980 262890 265032 262896
rect 264992 258097 265020 262890
rect 264978 258088 265034 258097
rect 264978 258023 265034 258032
rect 264980 201476 265032 201482
rect 264980 201418 265032 201424
rect 264992 189990 265020 201418
rect 264980 189984 265032 189990
rect 264980 189926 265032 189932
rect 265084 14754 265112 335582
rect 265268 335566 265480 335594
rect 265900 335640 265952 335646
rect 265900 335582 265952 335588
rect 266452 335640 266504 335646
rect 266924 335594 266952 340054
rect 267384 335646 267412 340054
rect 268212 336938 268240 340068
rect 268396 340054 268686 340082
rect 269146 340054 269252 340082
rect 268200 336932 268252 336938
rect 268200 336874 268252 336880
rect 266452 335582 266504 335588
rect 265268 335306 265296 335566
rect 265256 335300 265308 335306
rect 265256 335242 265308 335248
rect 265256 325712 265308 325718
rect 265256 325654 265308 325660
rect 265268 317506 265296 325654
rect 265268 317478 265388 317506
rect 265360 316062 265388 317478
rect 265164 316056 265216 316062
rect 265164 315998 265216 316004
rect 265348 316056 265400 316062
rect 265348 315998 265400 316004
rect 265176 314673 265204 315998
rect 265162 314664 265218 314673
rect 265162 314599 265218 314608
rect 265254 305008 265310 305017
rect 265254 304943 265310 304952
rect 265268 278798 265296 304943
rect 265164 278792 265216 278798
rect 265164 278734 265216 278740
rect 265256 278792 265308 278798
rect 265256 278734 265308 278740
rect 265176 262954 265204 278734
rect 265164 262948 265216 262954
rect 265164 262890 265216 262896
rect 265162 258088 265218 258097
rect 265162 258023 265218 258032
rect 265176 251258 265204 258023
rect 265164 251252 265216 251258
rect 265164 251194 265216 251200
rect 265256 251252 265308 251258
rect 265256 251194 265308 251200
rect 265268 246378 265296 251194
rect 265268 246350 265388 246378
rect 265360 231878 265388 246350
rect 265256 231872 265308 231878
rect 265256 231814 265308 231820
rect 265348 231872 265400 231878
rect 265348 231814 265400 231820
rect 265268 222290 265296 231814
rect 265256 222284 265308 222290
rect 265256 222226 265308 222232
rect 265164 222216 265216 222222
rect 265164 222158 265216 222164
rect 265176 212566 265204 222158
rect 265164 212560 265216 212566
rect 265164 212502 265216 212508
rect 265256 212560 265308 212566
rect 265256 212502 265308 212508
rect 265268 211138 265296 212502
rect 265256 211132 265308 211138
rect 265256 211074 265308 211080
rect 265256 202768 265308 202774
rect 265256 202710 265308 202716
rect 265268 201482 265296 202710
rect 265256 201476 265308 201482
rect 265256 201418 265308 201424
rect 265164 189984 265216 189990
rect 265164 189926 265216 189932
rect 265176 180810 265204 189926
rect 265164 180804 265216 180810
rect 265164 180746 265216 180752
rect 265256 180804 265308 180810
rect 265256 180746 265308 180752
rect 265268 179382 265296 180746
rect 265256 179376 265308 179382
rect 265256 179318 265308 179324
rect 265164 161492 265216 161498
rect 265164 161434 265216 161440
rect 265176 153202 265204 161434
rect 265164 153196 265216 153202
rect 265164 153138 265216 153144
rect 265348 153196 265400 153202
rect 265348 153138 265400 153144
rect 265360 137714 265388 153138
rect 265268 137686 265388 137714
rect 265268 125610 265296 137686
rect 265176 125594 265296 125610
rect 265164 125588 265296 125594
rect 265216 125582 265296 125588
rect 265348 125588 265400 125594
rect 265164 125530 265216 125536
rect 265348 125530 265400 125536
rect 265360 118402 265388 125530
rect 265268 118374 265388 118402
rect 265268 104922 265296 118374
rect 265256 104916 265308 104922
rect 265256 104858 265308 104864
rect 265348 104916 265400 104922
rect 265348 104858 265400 104864
rect 265360 85610 265388 104858
rect 265256 85604 265308 85610
rect 265256 85546 265308 85552
rect 265348 85604 265400 85610
rect 265348 85546 265400 85552
rect 265268 71074 265296 85546
rect 265176 71046 265296 71074
rect 265176 66230 265204 71046
rect 265164 66224 265216 66230
rect 265164 66166 265216 66172
rect 265256 46980 265308 46986
rect 265256 46922 265308 46928
rect 265268 45558 265296 46922
rect 265256 45552 265308 45558
rect 265256 45494 265308 45500
rect 265256 35964 265308 35970
rect 265256 35906 265308 35912
rect 265268 31822 265296 35906
rect 265256 31816 265308 31822
rect 265256 31758 265308 31764
rect 265256 31680 265308 31686
rect 265256 31622 265308 31628
rect 265268 27606 265296 31622
rect 265256 27600 265308 27606
rect 265256 27542 265308 27548
rect 265256 19304 265308 19310
rect 265256 19246 265308 19252
rect 265268 17950 265296 19246
rect 265256 17944 265308 17950
rect 265256 17886 265308 17892
rect 265440 17944 265492 17950
rect 265440 17886 265492 17892
rect 265072 14748 265124 14754
rect 265072 14690 265124 14696
rect 265452 9625 265480 17886
rect 266464 14822 266492 335582
rect 266740 335566 266952 335594
rect 267372 335640 267424 335646
rect 268396 335594 268424 340054
rect 269028 337408 269080 337414
rect 269028 337350 269080 337356
rect 267372 335582 267424 335588
rect 267844 335566 268424 335594
rect 266740 317506 266768 335566
rect 267844 317506 267872 335566
rect 266648 317478 266768 317506
rect 267752 317478 267872 317506
rect 266648 317422 266676 317478
rect 267752 317422 267780 317478
rect 266636 317416 266688 317422
rect 266636 317358 266688 317364
rect 266728 317416 266780 317422
rect 266728 317358 266780 317364
rect 267740 317416 267792 317422
rect 267740 317358 267792 317364
rect 267832 317416 267884 317422
rect 267832 317358 267884 317364
rect 266740 260914 266768 317358
rect 267844 316033 267872 317358
rect 267830 316024 267886 316033
rect 267830 315959 267886 315968
rect 268014 316024 268070 316033
rect 268014 315959 268070 315968
rect 268028 306406 268056 315959
rect 267832 306400 267884 306406
rect 267832 306342 267884 306348
rect 268016 306400 268068 306406
rect 268016 306342 268068 306348
rect 267844 302954 267872 306342
rect 267844 302926 267964 302954
rect 267936 289882 267964 302926
rect 267832 289876 267884 289882
rect 267832 289818 267884 289824
rect 267924 289876 267976 289882
rect 267924 289818 267976 289824
rect 267844 278798 267872 289818
rect 267740 278792 267792 278798
rect 267740 278734 267792 278740
rect 267832 278792 267884 278798
rect 267832 278734 267884 278740
rect 267752 277409 267780 278734
rect 267738 277400 267794 277409
rect 267738 277335 267794 277344
rect 268014 277400 268070 277409
rect 268014 277335 268070 277344
rect 268028 267782 268056 277335
rect 267832 267776 267884 267782
rect 267832 267718 267884 267724
rect 268016 267776 268068 267782
rect 268016 267718 268068 267724
rect 266728 260908 266780 260914
rect 266728 260850 266780 260856
rect 266728 260772 266780 260778
rect 266728 260714 266780 260720
rect 266740 251190 266768 260714
rect 267844 259486 267872 267718
rect 267740 259480 267792 259486
rect 267740 259422 267792 259428
rect 267832 259480 267884 259486
rect 267832 259422 267884 259428
rect 267752 251258 267780 259422
rect 267740 251252 267792 251258
rect 267740 251194 267792 251200
rect 267832 251252 267884 251258
rect 267832 251194 267884 251200
rect 266728 251184 266780 251190
rect 266728 251126 266780 251132
rect 266728 251048 266780 251054
rect 266728 250990 266780 250996
rect 266740 231946 266768 250990
rect 267844 246378 267872 251194
rect 267844 246350 267964 246378
rect 267936 240145 267964 246350
rect 267922 240136 267978 240145
rect 267922 240071 267978 240080
rect 268106 240136 268162 240145
rect 268106 240071 268162 240080
rect 266728 231940 266780 231946
rect 266728 231882 266780 231888
rect 268120 230518 268148 240071
rect 266728 230512 266780 230518
rect 266728 230454 266780 230460
rect 267924 230512 267976 230518
rect 267924 230454 267976 230460
rect 268108 230512 268160 230518
rect 268108 230454 268160 230460
rect 266740 217410 266768 230454
rect 267936 220862 267964 230454
rect 267740 220856 267792 220862
rect 267740 220798 267792 220804
rect 267924 220856 267976 220862
rect 267924 220798 267976 220804
rect 266740 217382 266860 217410
rect 266832 212566 266860 217382
rect 267752 212566 267780 220798
rect 266636 212560 266688 212566
rect 266636 212502 266688 212508
rect 266820 212560 266872 212566
rect 266820 212502 266872 212508
rect 267740 212560 267792 212566
rect 267740 212502 267792 212508
rect 267832 212560 267884 212566
rect 267832 212502 267884 212508
rect 266648 201482 266676 212502
rect 267752 202910 267780 202941
rect 267844 202910 267872 212502
rect 267740 202904 267792 202910
rect 267832 202904 267884 202910
rect 267792 202852 267832 202858
rect 267740 202846 267884 202852
rect 267752 202830 267872 202846
rect 266636 201476 266688 201482
rect 266636 201418 266688 201424
rect 266820 201476 266872 201482
rect 266820 201418 266872 201424
rect 266832 186266 266860 201418
rect 267844 198098 267872 202830
rect 267752 198070 267872 198098
rect 267752 186386 267780 198070
rect 267740 186380 267792 186386
rect 267740 186322 267792 186328
rect 266740 186238 266860 186266
rect 266740 174078 266768 186238
rect 267740 183592 267792 183598
rect 267738 183560 267740 183569
rect 267792 183560 267794 183569
rect 267738 183495 267794 183504
rect 267922 183560 267978 183569
rect 267922 183495 267978 183504
rect 266728 174072 266780 174078
rect 266728 174014 266780 174020
rect 267936 173942 267964 183495
rect 266636 173936 266688 173942
rect 266636 173878 266688 173884
rect 267832 173936 267884 173942
rect 267832 173878 267884 173884
rect 267924 173936 267976 173942
rect 267924 173878 267976 173884
rect 266648 171034 266676 173878
rect 266648 171006 266768 171034
rect 266740 153218 266768 171006
rect 267844 164234 267872 173878
rect 267752 164206 267872 164234
rect 267752 157418 267780 164206
rect 267740 157412 267792 157418
rect 267740 157354 267792 157360
rect 267740 157276 267792 157282
rect 267740 157218 267792 157224
rect 266648 153202 266768 153218
rect 266636 153196 266768 153202
rect 266688 153190 266768 153196
rect 266636 153138 266688 153144
rect 266648 153107 266676 153138
rect 267752 144906 267780 157218
rect 266636 144900 266688 144906
rect 266636 144842 266688 144848
rect 267740 144900 267792 144906
rect 267740 144842 267792 144848
rect 267924 144900 267976 144906
rect 267924 144842 267976 144848
rect 266648 143562 266676 144842
rect 266648 143534 266768 143562
rect 266740 138394 266768 143534
rect 267936 139890 267964 144842
rect 267844 139862 267964 139890
rect 266740 138366 266860 138394
rect 266832 135289 266860 138366
rect 266634 135280 266690 135289
rect 266634 135215 266690 135224
rect 266818 135280 266874 135289
rect 267844 135250 267872 139862
rect 266818 135215 266874 135224
rect 267740 135244 267792 135250
rect 266648 134722 266676 135215
rect 267740 135186 267792 135192
rect 267832 135244 267884 135250
rect 267832 135186 267884 135192
rect 266648 134694 266860 134722
rect 266832 128330 266860 134694
rect 266740 128302 266860 128330
rect 266740 125576 266768 128302
rect 267752 125594 267780 135186
rect 267740 125588 267792 125594
rect 266740 125548 266860 125576
rect 266832 115977 266860 125548
rect 267740 125530 267792 125536
rect 267924 125588 267976 125594
rect 267924 125530 267976 125536
rect 267936 120578 267964 125530
rect 267844 120550 267964 120578
rect 266634 115968 266690 115977
rect 266634 115903 266690 115912
rect 266818 115968 266874 115977
rect 266818 115903 266874 115912
rect 266648 109070 266676 115903
rect 267844 114510 267872 120550
rect 267832 114504 267884 114510
rect 267832 114446 267884 114452
rect 266636 109064 266688 109070
rect 266636 109006 266688 109012
rect 266728 108996 266780 109002
rect 266728 108938 266780 108944
rect 266740 96801 266768 108938
rect 266726 96792 266782 96801
rect 266726 96727 266782 96736
rect 266634 96656 266690 96665
rect 266634 96591 266690 96600
rect 266648 95198 266676 96591
rect 266636 95192 266688 95198
rect 266636 95134 266688 95140
rect 267740 93900 267792 93906
rect 267740 93842 267792 93848
rect 267752 85610 267780 93842
rect 266728 85604 266780 85610
rect 266728 85546 266780 85552
rect 267740 85604 267792 85610
rect 267740 85546 267792 85552
rect 267832 85604 267884 85610
rect 267832 85546 267884 85552
rect 266740 84182 266768 85546
rect 267844 84182 267872 85546
rect 266728 84176 266780 84182
rect 266728 84118 266780 84124
rect 267832 84176 267884 84182
rect 267832 84118 267884 84124
rect 266820 74588 266872 74594
rect 266820 74530 266872 74536
rect 267740 74588 267792 74594
rect 267740 74530 267792 74536
rect 266832 66298 266860 74530
rect 266636 66292 266688 66298
rect 266636 66234 266688 66240
rect 266820 66292 266872 66298
rect 266820 66234 266872 66240
rect 266648 61470 266676 66234
rect 267752 64870 267780 74530
rect 267740 64864 267792 64870
rect 267740 64806 267792 64812
rect 266636 61464 266688 61470
rect 266636 61406 266688 61412
rect 268108 55276 268160 55282
rect 268108 55218 268160 55224
rect 266636 48340 266688 48346
rect 266636 48282 266688 48288
rect 266648 42106 266676 48282
rect 268120 45966 268148 55218
rect 268108 45960 268160 45966
rect 268108 45902 268160 45908
rect 267832 45620 267884 45626
rect 267832 45562 267884 45568
rect 266648 42078 266860 42106
rect 266832 31618 266860 42078
rect 267844 37262 267872 45562
rect 267832 37256 267884 37262
rect 267832 37198 267884 37204
rect 268016 37256 268068 37262
rect 268016 37198 268068 37204
rect 266636 31612 266688 31618
rect 266636 31554 266688 31560
rect 266820 31612 266872 31618
rect 266820 31554 266872 31560
rect 266648 17898 266676 31554
rect 267740 29232 267792 29238
rect 267738 29200 267740 29209
rect 267792 29200 267794 29209
rect 267738 29135 267794 29144
rect 268028 27742 268056 37198
rect 268016 27736 268068 27742
rect 268016 27678 268068 27684
rect 267924 27600 267976 27606
rect 267924 27542 267976 27548
rect 267936 26246 267964 27542
rect 267924 26240 267976 26246
rect 267924 26182 267976 26188
rect 266648 17870 266768 17898
rect 266452 14816 266504 14822
rect 266452 14758 266504 14764
rect 266740 10606 266768 17870
rect 266728 10600 266780 10606
rect 266728 10542 266780 10548
rect 265254 9616 265310 9625
rect 265254 9551 265310 9560
rect 265438 9616 265494 9625
rect 265438 9551 265494 9560
rect 265268 8378 265296 9551
rect 265176 8350 265296 8378
rect 265176 8294 265204 8350
rect 265164 8288 265216 8294
rect 265164 8230 265216 8236
rect 263876 8220 263928 8226
rect 263876 8162 263928 8168
rect 267004 8220 267056 8226
rect 267004 8162 267056 8168
rect 262404 8152 262456 8158
rect 262404 8094 262456 8100
rect 263416 8152 263468 8158
rect 263416 8094 263468 8100
rect 262220 3664 262272 3670
rect 262220 3606 262272 3612
rect 261484 2848 261536 2854
rect 261484 2790 261536 2796
rect 261024 1148 261076 1154
rect 261024 1090 261076 1096
rect 261036 480 261064 1090
rect 262232 480 262260 3606
rect 263428 480 263456 8094
rect 264612 3868 264664 3874
rect 264612 3810 264664 3816
rect 264624 480 264652 3810
rect 265808 3596 265860 3602
rect 265808 3538 265860 3544
rect 265820 480 265848 3538
rect 267016 480 267044 8162
rect 269040 4146 269068 337350
rect 269224 14890 269252 340054
rect 269684 337482 269712 340068
rect 269868 340054 270158 340082
rect 269672 337476 269724 337482
rect 269672 337418 269724 337424
rect 269868 335594 269896 340054
rect 269316 335566 269896 335594
rect 269212 14884 269264 14890
rect 269212 14826 269264 14832
rect 269316 10742 269344 335566
rect 270498 183560 270554 183569
rect 270498 183495 270554 183504
rect 270512 174010 270540 183495
rect 270500 174004 270552 174010
rect 270500 173946 270552 173952
rect 270500 169108 270552 169114
rect 270500 169050 270552 169056
rect 270512 164257 270540 169050
rect 270498 164248 270554 164257
rect 270498 164183 270554 164192
rect 270500 98116 270552 98122
rect 270500 98058 270552 98064
rect 270512 75954 270540 98058
rect 270500 75948 270552 75954
rect 270500 75890 270552 75896
rect 270500 22160 270552 22166
rect 270500 22102 270552 22108
rect 270512 10810 270540 22102
rect 270604 18018 270632 340068
rect 271156 337142 271184 340068
rect 271248 340054 271630 340082
rect 271984 340054 272090 340082
rect 271144 337136 271196 337142
rect 271144 337078 271196 337084
rect 271248 334354 271276 340054
rect 271788 337476 271840 337482
rect 271788 337418 271840 337424
rect 271328 337272 271380 337278
rect 271328 337214 271380 337220
rect 271236 334348 271288 334354
rect 271236 334290 271288 334296
rect 271340 334234 271368 337214
rect 271156 334206 271368 334234
rect 270776 328500 270828 328506
rect 270776 328442 270828 328448
rect 270788 307850 270816 328442
rect 270696 307822 270816 307850
rect 270696 302326 270724 307822
rect 270684 302320 270736 302326
rect 270684 302262 270736 302268
rect 270776 302116 270828 302122
rect 270776 302058 270828 302064
rect 270788 289814 270816 302058
rect 270684 289808 270736 289814
rect 270684 289750 270736 289756
rect 270776 289808 270828 289814
rect 270776 289750 270828 289756
rect 270696 280158 270724 289750
rect 270684 280152 270736 280158
rect 270684 280094 270736 280100
rect 270684 275324 270736 275330
rect 270684 275266 270736 275272
rect 270696 263634 270724 275266
rect 270684 263628 270736 263634
rect 270684 263570 270736 263576
rect 270684 263492 270736 263498
rect 270684 263434 270736 263440
rect 270696 260846 270724 263434
rect 270684 260840 270736 260846
rect 270684 260782 270736 260788
rect 270684 256012 270736 256018
rect 270684 255954 270736 255960
rect 270696 244322 270724 255954
rect 270684 244316 270736 244322
rect 270684 244258 270736 244264
rect 270684 241596 270736 241602
rect 270684 241538 270736 241544
rect 270696 241466 270724 241538
rect 270684 241460 270736 241466
rect 270684 241402 270736 241408
rect 270684 232076 270736 232082
rect 270684 232018 270736 232024
rect 270696 225010 270724 232018
rect 270684 225004 270736 225010
rect 270684 224946 270736 224952
rect 270684 222284 270736 222290
rect 270684 222226 270736 222232
rect 270696 222154 270724 222226
rect 270684 222148 270736 222154
rect 270684 222090 270736 222096
rect 270684 212764 270736 212770
rect 270684 212706 270736 212712
rect 270696 202881 270724 212706
rect 270682 202872 270738 202881
rect 270682 202807 270738 202816
rect 270682 202736 270738 202745
rect 270682 202671 270738 202680
rect 270696 186386 270724 202671
rect 270684 186380 270736 186386
rect 270684 186322 270736 186328
rect 270684 183592 270736 183598
rect 270682 183560 270684 183569
rect 270736 183560 270738 183569
rect 270682 183495 270738 183504
rect 270684 174004 270736 174010
rect 270684 173946 270736 173952
rect 270696 169114 270724 173946
rect 270684 169108 270736 169114
rect 270684 169050 270736 169056
rect 270682 164248 270738 164257
rect 270682 164183 270738 164192
rect 270696 157214 270724 164183
rect 270684 157208 270736 157214
rect 270684 157150 270736 157156
rect 270776 157140 270828 157146
rect 270776 157082 270828 157088
rect 270788 147914 270816 157082
rect 270696 147886 270816 147914
rect 270696 144906 270724 147886
rect 270684 144900 270736 144906
rect 270684 144842 270736 144848
rect 270960 144900 271012 144906
rect 270960 144842 271012 144848
rect 270972 143546 271000 144842
rect 270960 143540 271012 143546
rect 270960 143482 271012 143488
rect 270960 135108 271012 135114
rect 270960 135050 271012 135056
rect 270972 125633 271000 135050
rect 270682 125624 270738 125633
rect 270682 125559 270684 125568
rect 270736 125559 270738 125568
rect 270958 125624 271014 125633
rect 270958 125559 270960 125568
rect 270684 125530 270736 125536
rect 271012 125559 271014 125568
rect 270960 125530 271012 125536
rect 270972 115938 271000 125530
rect 270684 115932 270736 115938
rect 270684 115874 270736 115880
rect 270960 115932 271012 115938
rect 270960 115874 271012 115880
rect 270696 106282 270724 115874
rect 270684 106276 270736 106282
rect 270684 106218 270736 106224
rect 270960 106276 271012 106282
rect 270960 106218 271012 106224
rect 270972 98122 271000 106218
rect 270960 98116 271012 98122
rect 270960 98058 271012 98064
rect 270684 75948 270736 75954
rect 270684 75890 270736 75896
rect 270696 66366 270724 75890
rect 270684 66360 270736 66366
rect 270684 66302 270736 66308
rect 270776 66292 270828 66298
rect 270776 66234 270828 66240
rect 270788 57882 270816 66234
rect 270696 57854 270816 57882
rect 270696 38690 270724 57854
rect 270684 38684 270736 38690
rect 270684 38626 270736 38632
rect 270776 38684 270828 38690
rect 270776 38626 270828 38632
rect 270788 22166 270816 38626
rect 270776 22160 270828 22166
rect 270776 22102 270828 22108
rect 270592 18012 270644 18018
rect 270592 17954 270644 17960
rect 270592 17876 270644 17882
rect 270592 17818 270644 17824
rect 270604 14958 270632 17818
rect 270592 14952 270644 14958
rect 270592 14894 270644 14900
rect 270500 10804 270552 10810
rect 270500 10746 270552 10752
rect 269304 10736 269356 10742
rect 269304 10678 269356 10684
rect 270500 8288 270552 8294
rect 270500 8230 270552 8236
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 269028 4140 269080 4146
rect 269028 4082 269080 4088
rect 268120 480 268148 4082
rect 269304 3256 269356 3262
rect 269304 3198 269356 3204
rect 269316 480 269344 3198
rect 270512 480 270540 8230
rect 271156 4418 271184 334206
rect 271144 4412 271196 4418
rect 271144 4354 271196 4360
rect 271800 626 271828 337418
rect 271984 18018 272012 340054
rect 272628 337346 272656 340068
rect 272720 340054 273102 340082
rect 273364 340054 273562 340082
rect 272616 337340 272668 337346
rect 272616 337282 272668 337288
rect 272720 334354 272748 340054
rect 272800 337340 272852 337346
rect 272800 337282 272852 337288
rect 272708 334348 272760 334354
rect 272708 334290 272760 334296
rect 272812 334234 272840 337282
rect 272536 334206 272840 334234
rect 272248 328500 272300 328506
rect 272248 328442 272300 328448
rect 272260 312610 272288 328442
rect 272168 312582 272288 312610
rect 272168 302326 272196 312582
rect 272156 302320 272208 302326
rect 272156 302262 272208 302268
rect 272248 302116 272300 302122
rect 272248 302058 272300 302064
rect 272260 289814 272288 302058
rect 272248 289808 272300 289814
rect 272248 289750 272300 289756
rect 272340 283620 272392 283626
rect 272340 283562 272392 283568
rect 272352 278769 272380 283562
rect 272154 278760 272210 278769
rect 272154 278695 272210 278704
rect 272338 278760 272394 278769
rect 272338 278695 272394 278704
rect 272168 270042 272196 278695
rect 272168 270014 272380 270042
rect 272352 260982 272380 270014
rect 272340 260976 272392 260982
rect 272340 260918 272392 260924
rect 272156 260772 272208 260778
rect 272156 260714 272208 260720
rect 272168 244390 272196 260714
rect 272156 244384 272208 244390
rect 272156 244326 272208 244332
rect 272156 244248 272208 244254
rect 272156 244190 272208 244196
rect 272168 241505 272196 244190
rect 272154 241496 272210 241505
rect 272154 241431 272210 241440
rect 272338 241360 272394 241369
rect 272338 241295 272394 241304
rect 272352 231826 272380 241295
rect 272076 231798 272380 231826
rect 272076 224890 272104 231798
rect 272076 224862 272196 224890
rect 272168 222193 272196 224862
rect 272154 222184 272210 222193
rect 272154 222119 272210 222128
rect 272246 222048 272302 222057
rect 272246 221983 272302 221992
rect 272260 220810 272288 221983
rect 272168 220782 272288 220810
rect 272168 212566 272196 220782
rect 272156 212560 272208 212566
rect 272156 212502 272208 212508
rect 272156 211200 272208 211206
rect 272156 211142 272208 211148
rect 272168 202881 272196 211142
rect 272154 202872 272210 202881
rect 272154 202807 272210 202816
rect 272246 202736 272302 202745
rect 272246 202671 272302 202680
rect 272260 186538 272288 202671
rect 272168 186510 272288 186538
rect 272168 183598 272196 186510
rect 272156 183592 272208 183598
rect 272156 183534 272208 183540
rect 272248 183524 272300 183530
rect 272248 183466 272300 183472
rect 272260 173890 272288 183466
rect 272168 173862 272288 173890
rect 272168 167074 272196 173862
rect 272156 167068 272208 167074
rect 272156 167010 272208 167016
rect 272248 167000 272300 167006
rect 272248 166942 272300 166948
rect 272260 164257 272288 166942
rect 272062 164248 272118 164257
rect 272062 164183 272118 164192
rect 272246 164248 272302 164257
rect 272246 164183 272302 164192
rect 272076 162858 272104 164183
rect 272064 162852 272116 162858
rect 272064 162794 272116 162800
rect 272248 154556 272300 154562
rect 272248 154498 272300 154504
rect 272260 153218 272288 154498
rect 272168 153190 272288 153218
rect 272168 144906 272196 153190
rect 272156 144900 272208 144906
rect 272156 144842 272208 144848
rect 272432 144900 272484 144906
rect 272432 144842 272484 144848
rect 272444 143546 272472 144842
rect 272340 143540 272392 143546
rect 272340 143482 272392 143488
rect 272432 143540 272484 143546
rect 272432 143482 272484 143488
rect 272352 133929 272380 143482
rect 272154 133920 272210 133929
rect 272154 133855 272210 133864
rect 272338 133920 272394 133929
rect 272338 133855 272394 133864
rect 272168 125594 272196 133855
rect 272156 125588 272208 125594
rect 272156 125530 272208 125536
rect 272432 125588 272484 125594
rect 272432 125530 272484 125536
rect 272444 124166 272472 125530
rect 272432 124160 272484 124166
rect 272432 124102 272484 124108
rect 272156 114572 272208 114578
rect 272156 114514 272208 114520
rect 272168 106282 272196 114514
rect 272156 106276 272208 106282
rect 272156 106218 272208 106224
rect 272432 106276 272484 106282
rect 272432 106218 272484 106224
rect 272444 103494 272472 106218
rect 272432 103488 272484 103494
rect 272432 103430 272484 103436
rect 272340 93900 272392 93906
rect 272340 93842 272392 93848
rect 272352 85610 272380 93842
rect 272156 85604 272208 85610
rect 272156 85546 272208 85552
rect 272340 85604 272392 85610
rect 272340 85546 272392 85552
rect 272168 82634 272196 85546
rect 272168 82606 272288 82634
rect 272260 72486 272288 82606
rect 272248 72480 272300 72486
rect 272248 72422 272300 72428
rect 272156 67652 272208 67658
rect 272156 67594 272208 67600
rect 272168 58070 272196 67594
rect 272156 58064 272208 58070
rect 272156 58006 272208 58012
rect 272156 57928 272208 57934
rect 272156 57870 272208 57876
rect 272168 38690 272196 57870
rect 272156 38684 272208 38690
rect 272156 38626 272208 38632
rect 272248 38684 272300 38690
rect 272248 38626 272300 38632
rect 272260 22250 272288 38626
rect 272260 22222 272380 22250
rect 271972 18012 272024 18018
rect 271972 17954 272024 17960
rect 271972 17876 272024 17882
rect 271972 17818 272024 17824
rect 271880 17808 271932 17814
rect 271880 17750 271932 17756
rect 271892 10878 271920 17750
rect 271984 15026 272012 17818
rect 272352 17814 272380 22222
rect 272340 17808 272392 17814
rect 272340 17750 272392 17756
rect 271972 15020 272024 15026
rect 271972 14962 272024 14968
rect 271880 10872 271932 10878
rect 271880 10814 271932 10820
rect 272536 4350 272564 334206
rect 273260 317416 273312 317422
rect 273260 317358 273312 317364
rect 273272 316033 273300 317358
rect 273074 316024 273130 316033
rect 273074 315959 273130 315968
rect 273258 316024 273314 316033
rect 273258 315959 273314 315968
rect 273088 306406 273116 315959
rect 273076 306400 273128 306406
rect 273076 306342 273128 306348
rect 273260 306400 273312 306406
rect 273260 306342 273312 306348
rect 273272 296750 273300 306342
rect 273260 296744 273312 296750
rect 273260 296686 273312 296692
rect 273364 15094 273392 340054
rect 274100 337006 274128 340068
rect 274284 340054 274574 340082
rect 274744 340054 275034 340082
rect 274088 337000 274140 337006
rect 274088 336942 274140 336948
rect 274284 331242 274312 340054
rect 273640 331214 274312 331242
rect 273640 327078 273668 331214
rect 273628 327072 273680 327078
rect 273628 327014 273680 327020
rect 273536 321564 273588 321570
rect 273536 321506 273588 321512
rect 273548 317422 273576 321506
rect 273536 317416 273588 317422
rect 273536 317358 273588 317364
rect 273548 296750 273576 296781
rect 273536 296744 273588 296750
rect 273588 296692 273668 296698
rect 273536 296686 273668 296692
rect 273548 296682 273668 296686
rect 273548 296676 273680 296682
rect 273548 296670 273628 296676
rect 273628 296618 273680 296624
rect 273628 287088 273680 287094
rect 273628 287030 273680 287036
rect 273640 285002 273668 287030
rect 273548 284974 273668 285002
rect 273548 280158 273576 284974
rect 273536 280152 273588 280158
rect 273536 280094 273588 280100
rect 273628 270564 273680 270570
rect 273628 270506 273680 270512
rect 273640 263514 273668 270506
rect 273548 263486 273668 263514
rect 273548 260846 273576 263486
rect 273536 260840 273588 260846
rect 273536 260782 273588 260788
rect 273628 251252 273680 251258
rect 273628 251194 273680 251200
rect 273640 244202 273668 251194
rect 273548 244174 273668 244202
rect 273548 236722 273576 244174
rect 273548 236694 273668 236722
rect 273640 224890 273668 236694
rect 273548 224862 273668 224890
rect 273548 217410 273576 224862
rect 273548 217382 273668 217410
rect 273640 205578 273668 217382
rect 273548 205550 273668 205578
rect 273548 202858 273576 205550
rect 273548 202830 273668 202858
rect 273640 186266 273668 202830
rect 273548 186238 273668 186266
rect 273548 183546 273576 186238
rect 273548 183518 273668 183546
rect 273640 166954 273668 183518
rect 273548 166926 273668 166954
rect 273548 157486 273576 166926
rect 273536 157480 273588 157486
rect 273536 157422 273588 157428
rect 273536 157344 273588 157350
rect 273536 157286 273588 157292
rect 273548 144906 273576 157286
rect 273536 144900 273588 144906
rect 273536 144842 273588 144848
rect 273536 137964 273588 137970
rect 273536 137906 273588 137912
rect 273548 135266 273576 137906
rect 273548 135238 273668 135266
rect 273640 128330 273668 135238
rect 273548 128302 273668 128330
rect 273548 125594 273576 128302
rect 273536 125588 273588 125594
rect 273536 125530 273588 125536
rect 273536 116000 273588 116006
rect 273536 115942 273588 115948
rect 273548 106282 273576 115942
rect 273536 106276 273588 106282
rect 273536 106218 273588 106224
rect 273536 99340 273588 99346
rect 273536 99282 273588 99288
rect 273548 96642 273576 99282
rect 273548 96614 273668 96642
rect 273640 79914 273668 96614
rect 273548 79886 273668 79914
rect 273548 72434 273576 79886
rect 273548 72406 273760 72434
rect 273732 70258 273760 72406
rect 273640 70230 273760 70258
rect 273640 67590 273668 70230
rect 273628 67584 273680 67590
rect 273628 67526 273680 67532
rect 273628 57996 273680 58002
rect 273628 57938 273680 57944
rect 273640 51218 273668 57938
rect 273640 51190 273760 51218
rect 273732 50946 273760 51190
rect 273548 50918 273760 50946
rect 273548 48278 273576 50918
rect 273536 48272 273588 48278
rect 273536 48214 273588 48220
rect 273536 38684 273588 38690
rect 273536 38626 273588 38632
rect 273548 22114 273576 38626
rect 273456 22086 273576 22114
rect 273456 17950 273484 22086
rect 273444 17944 273496 17950
rect 273444 17886 273496 17892
rect 274744 15162 274772 340054
rect 275572 337550 275600 340068
rect 275560 337544 275612 337550
rect 275560 337486 275612 337492
rect 275928 337544 275980 337550
rect 275928 337486 275980 337492
rect 275558 63880 275614 63889
rect 275558 63815 275614 63824
rect 275572 63617 275600 63815
rect 275558 63608 275614 63617
rect 275558 63543 275614 63552
rect 274732 15156 274784 15162
rect 274732 15098 274784 15104
rect 273352 15088 273404 15094
rect 273352 15030 273404 15036
rect 274088 6180 274140 6186
rect 274088 6122 274140 6128
rect 272524 4344 272576 4350
rect 272524 4286 272576 4292
rect 272892 3188 272944 3194
rect 272892 3130 272944 3136
rect 271708 598 271828 626
rect 271708 480 271736 598
rect 272904 480 272932 3130
rect 274100 480 274128 6122
rect 275940 2922 275968 337486
rect 276032 11014 276060 340068
rect 276124 340054 276506 340082
rect 276124 14414 276152 340054
rect 277044 337686 277072 340068
rect 277518 340054 277624 340082
rect 277032 337680 277084 337686
rect 277032 337622 277084 337628
rect 277306 29336 277362 29345
rect 277306 29271 277362 29280
rect 277320 29238 277348 29271
rect 277308 29232 277360 29238
rect 277308 29174 277360 29180
rect 276112 14408 276164 14414
rect 276112 14350 276164 14356
rect 276020 11008 276072 11014
rect 276020 10950 276072 10956
rect 277596 10266 277624 340054
rect 277688 340054 277978 340082
rect 277688 14346 277716 340054
rect 278516 336870 278544 340068
rect 278792 340054 278990 340082
rect 279068 340054 279450 340082
rect 278504 336864 278556 336870
rect 278504 336806 278556 336812
rect 278792 334830 278820 340054
rect 278780 334824 278832 334830
rect 278780 334766 278832 334772
rect 278964 334824 279016 334830
rect 278964 334766 279016 334772
rect 278872 328500 278924 328506
rect 278872 328442 278924 328448
rect 278778 110800 278834 110809
rect 278778 110735 278834 110744
rect 278792 110673 278820 110735
rect 278778 110664 278834 110673
rect 278778 110599 278834 110608
rect 278884 109154 278912 328442
rect 278792 109126 278912 109154
rect 278792 109002 278820 109126
rect 278780 108996 278832 109002
rect 278780 108938 278832 108944
rect 278872 99408 278924 99414
rect 278872 99350 278924 99356
rect 278884 80186 278912 99350
rect 278792 80158 278912 80186
rect 278792 80050 278820 80158
rect 278792 80022 278912 80050
rect 278884 31770 278912 80022
rect 278792 31742 278912 31770
rect 277676 14340 277728 14346
rect 277676 14282 277728 14288
rect 278792 14278 278820 31742
rect 278780 14272 278832 14278
rect 278780 14214 278832 14220
rect 277584 10260 277636 10266
rect 277584 10202 277636 10208
rect 278976 10198 279004 334766
rect 279068 328506 279096 340054
rect 279988 337618 280016 340068
rect 280356 340054 280462 340082
rect 280632 340054 280922 340082
rect 281184 340054 281474 340082
rect 281644 340054 281934 340082
rect 282104 340054 282394 340082
rect 282946 340054 283144 340082
rect 279976 337612 280028 337618
rect 279976 337554 280028 337560
rect 280252 335640 280304 335646
rect 280252 335582 280304 335588
rect 279056 328500 279108 328506
rect 279056 328442 279108 328448
rect 279056 108996 279108 109002
rect 279056 108938 279108 108944
rect 279068 99414 279096 108938
rect 279056 99408 279108 99414
rect 279056 99350 279108 99356
rect 279974 40352 280030 40361
rect 280158 40352 280214 40361
rect 280030 40310 280158 40338
rect 279974 40287 280030 40296
rect 280158 40287 280214 40296
rect 280264 14210 280292 335582
rect 280252 14204 280304 14210
rect 280252 14146 280304 14152
rect 278964 10192 279016 10198
rect 278964 10134 279016 10140
rect 280356 10130 280384 340054
rect 280632 335646 280660 340054
rect 281184 336802 281212 340054
rect 281448 337612 281500 337618
rect 281448 337554 281500 337560
rect 281172 336796 281224 336802
rect 281172 336738 281224 336744
rect 280620 335640 280672 335646
rect 280620 335582 280672 335588
rect 280344 10124 280396 10130
rect 280344 10066 280396 10072
rect 280068 6248 280120 6254
rect 280068 6190 280120 6196
rect 278872 3800 278924 3806
rect 278872 3742 278924 3748
rect 276480 3256 276532 3262
rect 276480 3198 276532 3204
rect 275284 2916 275336 2922
rect 275284 2858 275336 2864
rect 275928 2916 275980 2922
rect 275928 2858 275980 2864
rect 275296 480 275324 2858
rect 276492 480 276520 3198
rect 277676 3188 277728 3194
rect 277676 3130 277728 3136
rect 277688 480 277716 3130
rect 278884 480 278912 3742
rect 280080 480 280108 6190
rect 281460 610 281488 337554
rect 281540 335640 281592 335646
rect 281540 335582 281592 335588
rect 281552 11898 281580 335582
rect 281540 11892 281592 11898
rect 281540 11834 281592 11840
rect 281644 11830 281672 340054
rect 282104 335646 282132 340054
rect 282092 335640 282144 335646
rect 282092 335582 282144 335588
rect 283012 335640 283064 335646
rect 283012 335582 283064 335588
rect 281632 11824 281684 11830
rect 281632 11766 281684 11772
rect 283024 6662 283052 335582
rect 283116 7585 283144 340054
rect 283208 340054 283406 340082
rect 283576 340054 283866 340082
rect 283102 7576 283158 7585
rect 283102 7511 283158 7520
rect 283012 6656 283064 6662
rect 283012 6598 283064 6604
rect 283208 5370 283236 340054
rect 283576 335646 283604 340054
rect 284404 336734 284432 340068
rect 284588 340054 284878 340082
rect 285140 340054 285338 340082
rect 285798 340054 285904 340082
rect 284392 336728 284444 336734
rect 284392 336670 284444 336676
rect 283564 335640 283616 335646
rect 283564 335582 283616 335588
rect 284484 335232 284536 335238
rect 284484 335174 284536 335180
rect 284300 329588 284352 329594
rect 284300 329530 284352 329536
rect 283470 87136 283526 87145
rect 283654 87136 283710 87145
rect 283526 87094 283654 87122
rect 283470 87071 283526 87080
rect 283654 87071 283710 87080
rect 284312 5438 284340 329530
rect 284496 8945 284524 335174
rect 284588 329594 284616 340054
rect 285140 332586 285168 340054
rect 285588 337680 285640 337686
rect 285588 337622 285640 337628
rect 284668 332580 284720 332586
rect 284668 332522 284720 332528
rect 285128 332580 285180 332586
rect 285128 332522 285180 332528
rect 284576 329588 284628 329594
rect 284576 329530 284628 329536
rect 284680 327078 284708 332522
rect 284668 327072 284720 327078
rect 284668 327014 284720 327020
rect 284760 327072 284812 327078
rect 284760 327014 284812 327020
rect 284772 316010 284800 327014
rect 284680 315982 284800 316010
rect 284680 311914 284708 315982
rect 284668 311908 284720 311914
rect 284668 311850 284720 311856
rect 284576 306400 284628 306406
rect 284576 306342 284628 306348
rect 284588 289814 284616 306342
rect 284576 289808 284628 289814
rect 284576 289750 284628 289756
rect 284760 289740 284812 289746
rect 284760 289682 284812 289688
rect 284772 280158 284800 289682
rect 284576 280152 284628 280158
rect 284576 280094 284628 280100
rect 284760 280152 284812 280158
rect 284760 280094 284812 280100
rect 284588 278769 284616 280094
rect 284574 278760 284630 278769
rect 284574 278695 284630 278704
rect 284758 278760 284814 278769
rect 284758 278695 284814 278704
rect 284772 269142 284800 278695
rect 284576 269136 284628 269142
rect 284576 269078 284628 269084
rect 284760 269136 284812 269142
rect 284760 269078 284812 269084
rect 284588 260914 284616 269078
rect 284576 260908 284628 260914
rect 284576 260850 284628 260856
rect 284760 260908 284812 260914
rect 284760 260850 284812 260856
rect 284772 249898 284800 260850
rect 284668 249892 284720 249898
rect 284668 249834 284720 249840
rect 284760 249892 284812 249898
rect 284760 249834 284812 249840
rect 284680 249762 284708 249834
rect 284668 249756 284720 249762
rect 284668 249698 284720 249704
rect 284852 240168 284904 240174
rect 284852 240110 284904 240116
rect 284864 225078 284892 240110
rect 284852 225072 284904 225078
rect 284852 225014 284904 225020
rect 284852 224936 284904 224942
rect 284852 224878 284904 224884
rect 284864 220833 284892 224878
rect 284666 220824 284722 220833
rect 284666 220759 284722 220768
rect 284850 220824 284906 220833
rect 284850 220759 284906 220768
rect 284680 212498 284708 220759
rect 284668 212492 284720 212498
rect 284668 212434 284720 212440
rect 284852 212492 284904 212498
rect 284852 212434 284904 212440
rect 284864 211154 284892 212434
rect 284864 211138 284984 211154
rect 284668 211132 284720 211138
rect 284864 211132 284996 211138
rect 284864 211126 284944 211132
rect 284668 211074 284720 211080
rect 284944 211074 284996 211080
rect 284680 209778 284708 211074
rect 284956 211043 284984 211074
rect 284668 209772 284720 209778
rect 284668 209714 284720 209720
rect 284760 209772 284812 209778
rect 284760 209714 284812 209720
rect 284772 200138 284800 209714
rect 284772 200122 284892 200138
rect 284668 200116 284720 200122
rect 284772 200116 284904 200122
rect 284772 200110 284852 200116
rect 284668 200058 284720 200064
rect 284852 200058 284904 200064
rect 284680 198694 284708 200058
rect 284668 198688 284720 198694
rect 284668 198630 284720 198636
rect 284668 183524 284720 183530
rect 284668 183466 284720 183472
rect 284680 180810 284708 183466
rect 284668 180804 284720 180810
rect 284668 180746 284720 180752
rect 284668 162920 284720 162926
rect 284668 162862 284720 162868
rect 284680 147762 284708 162862
rect 284668 147756 284720 147762
rect 284668 147698 284720 147704
rect 284668 147620 284720 147626
rect 284668 147562 284720 147568
rect 284680 132818 284708 147562
rect 284680 132790 284800 132818
rect 284772 132546 284800 132790
rect 284680 132518 284800 132546
rect 284680 132462 284708 132518
rect 284668 132456 284720 132462
rect 284668 132398 284720 132404
rect 284852 122868 284904 122874
rect 284852 122810 284904 122816
rect 284864 106350 284892 122810
rect 284852 106344 284904 106350
rect 284852 106286 284904 106292
rect 284760 106276 284812 106282
rect 284760 106218 284812 106224
rect 284772 95198 284800 106218
rect 284760 95192 284812 95198
rect 284760 95134 284812 95140
rect 284760 93900 284812 93906
rect 284760 93842 284812 93848
rect 284772 84182 284800 93842
rect 284760 84176 284812 84182
rect 284760 84118 284812 84124
rect 284668 66292 284720 66298
rect 284668 66234 284720 66240
rect 284680 57050 284708 66234
rect 284668 57044 284720 57050
rect 284668 56986 284720 56992
rect 284760 48340 284812 48346
rect 284760 48282 284812 48288
rect 284772 41478 284800 48282
rect 284760 41472 284812 41478
rect 284760 41414 284812 41420
rect 284668 41404 284720 41410
rect 284668 41346 284720 41352
rect 284680 29034 284708 41346
rect 284668 29028 284720 29034
rect 284668 28970 284720 28976
rect 284760 29028 284812 29034
rect 284760 28970 284812 28976
rect 284772 27606 284800 28970
rect 284760 27600 284812 27606
rect 284760 27542 284812 27548
rect 284576 18012 284628 18018
rect 284576 17954 284628 17960
rect 284482 8936 284538 8945
rect 284482 8871 284538 8880
rect 284588 7546 284616 17954
rect 284576 7540 284628 7546
rect 284576 7482 284628 7488
rect 284300 5432 284352 5438
rect 284300 5374 284352 5380
rect 283196 5364 283248 5370
rect 283196 5306 283248 5312
rect 283656 5296 283708 5302
rect 283656 5238 283708 5244
rect 282460 3936 282512 3942
rect 282460 3878 282512 3884
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281448 604 281500 610
rect 281448 546 281500 552
rect 281276 480 281304 546
rect 282472 480 282500 3878
rect 283668 480 283696 5238
rect 285600 4146 285628 337622
rect 285680 335640 285732 335646
rect 285680 335582 285732 335588
rect 285692 5506 285720 335582
rect 285772 306468 285824 306474
rect 285772 306410 285824 306416
rect 285784 296750 285812 306410
rect 285772 296744 285824 296750
rect 285772 296686 285824 296692
rect 285772 291916 285824 291922
rect 285772 291858 285824 291864
rect 285784 278798 285812 291858
rect 285772 278792 285824 278798
rect 285772 278734 285824 278740
rect 285770 202872 285826 202881
rect 285770 202807 285826 202816
rect 285784 198082 285812 202807
rect 285772 198076 285824 198082
rect 285772 198018 285824 198024
rect 285876 9314 285904 340054
rect 285968 340054 286350 340082
rect 286612 340054 286810 340082
rect 287164 340054 287270 340082
rect 287348 340054 287822 340082
rect 287992 340054 288282 340082
rect 288544 340054 288742 340082
rect 289004 340054 289294 340082
rect 289464 340054 289754 340082
rect 289832 340054 290214 340082
rect 285968 335646 285996 340054
rect 286612 335646 286640 340054
rect 285956 335640 286008 335646
rect 285956 335582 286008 335588
rect 286048 335640 286100 335646
rect 286048 335582 286100 335588
rect 286600 335640 286652 335646
rect 286600 335582 286652 335588
rect 287060 335640 287112 335646
rect 287060 335582 287112 335588
rect 286060 327078 286088 335582
rect 286048 327072 286100 327078
rect 286048 327014 286100 327020
rect 285956 317552 286008 317558
rect 285956 317494 286008 317500
rect 285968 311914 285996 317494
rect 285956 311908 286008 311914
rect 285956 311850 286008 311856
rect 286048 296744 286100 296750
rect 286048 296686 286100 296692
rect 286060 291922 286088 296686
rect 286048 291916 286100 291922
rect 286048 291858 286100 291864
rect 286048 278792 286100 278798
rect 286048 278734 286100 278740
rect 286060 261089 286088 278734
rect 286046 261080 286102 261089
rect 286046 261015 286102 261024
rect 285954 260944 286010 260953
rect 285954 260879 286010 260888
rect 285968 249830 285996 260879
rect 285956 249824 286008 249830
rect 286048 249824 286100 249830
rect 285956 249766 286008 249772
rect 286046 249792 286048 249801
rect 286100 249792 286102 249801
rect 286046 249727 286102 249736
rect 285954 249656 286010 249665
rect 285954 249591 286010 249600
rect 285968 245002 285996 249591
rect 285956 244996 286008 245002
rect 285956 244938 286008 244944
rect 285956 234524 286008 234530
rect 285956 234466 286008 234472
rect 285968 222193 285996 234466
rect 285954 222184 286010 222193
rect 285954 222119 286010 222128
rect 286138 222184 286194 222193
rect 286138 222119 286194 222128
rect 286152 220833 286180 222119
rect 285954 220824 286010 220833
rect 285954 220759 286010 220768
rect 286138 220824 286194 220833
rect 286138 220759 286194 220768
rect 285968 211834 285996 220759
rect 285968 211806 286180 211834
rect 286152 202910 286180 211806
rect 285956 202904 286008 202910
rect 285954 202872 285956 202881
rect 286140 202904 286192 202910
rect 286008 202872 286010 202881
rect 286140 202846 286192 202852
rect 285954 202807 286010 202816
rect 285956 198076 286008 198082
rect 285956 198018 286008 198024
rect 285968 183734 285996 198018
rect 285956 183728 286008 183734
rect 285956 183670 286008 183676
rect 285956 183592 286008 183598
rect 285956 183534 286008 183540
rect 285968 180810 285996 183534
rect 285956 180804 286008 180810
rect 285956 180746 286008 180752
rect 285956 175976 286008 175982
rect 285956 175918 286008 175924
rect 285968 153202 285996 175918
rect 285956 153196 286008 153202
rect 285956 153138 286008 153144
rect 286048 153196 286100 153202
rect 286048 153138 286100 153144
rect 286060 149410 286088 153138
rect 286060 149382 286180 149410
rect 286152 142118 286180 149382
rect 286140 142112 286192 142118
rect 286140 142054 286192 142060
rect 286048 132524 286100 132530
rect 286048 132466 286100 132472
rect 286060 129010 286088 132466
rect 285968 128982 286088 129010
rect 285968 124137 285996 128982
rect 285954 124128 286010 124137
rect 285954 124063 286010 124072
rect 286230 123992 286286 124001
rect 286230 123927 286286 123936
rect 286244 114510 286272 123927
rect 285956 114504 286008 114510
rect 285956 114446 286008 114452
rect 286232 114504 286284 114510
rect 286232 114446 286284 114452
rect 285968 95266 285996 114446
rect 285956 95260 286008 95266
rect 285956 95202 286008 95208
rect 286048 95260 286100 95266
rect 286048 95202 286100 95208
rect 286060 85592 286088 95202
rect 285968 85564 286088 85592
rect 285968 85490 285996 85564
rect 285968 85462 286088 85490
rect 286060 84182 286088 85462
rect 286048 84176 286100 84182
rect 286048 84118 286100 84124
rect 285956 66292 286008 66298
rect 285956 66234 286008 66240
rect 285968 61826 285996 66234
rect 285968 61798 286180 61826
rect 286152 61554 286180 61798
rect 286060 61526 286180 61554
rect 286060 56574 286088 61526
rect 286048 56568 286100 56574
rect 286048 56510 286100 56516
rect 285956 46980 286008 46986
rect 285956 46922 286008 46928
rect 285968 46866 285996 46922
rect 285968 46838 286088 46866
rect 286060 29102 286088 46838
rect 286048 29096 286100 29102
rect 286048 29038 286100 29044
rect 285956 29028 286008 29034
rect 285956 28970 286008 28976
rect 285968 27606 285996 28970
rect 285956 27600 286008 27606
rect 285956 27542 286008 27548
rect 285956 18012 286008 18018
rect 285956 17954 286008 17960
rect 285864 9308 285916 9314
rect 285864 9250 285916 9256
rect 285968 7478 285996 17954
rect 285956 7472 286008 7478
rect 285956 7414 286008 7420
rect 287072 7410 287100 335582
rect 287164 9382 287192 340054
rect 287348 11966 287376 340054
rect 287992 335646 288020 340054
rect 288256 337816 288308 337822
rect 288256 337758 288308 337764
rect 287980 335640 288032 335646
rect 287980 335582 288032 335588
rect 287336 11960 287388 11966
rect 287336 11902 287388 11908
rect 287152 9376 287204 9382
rect 287152 9318 287204 9324
rect 287060 7404 287112 7410
rect 287060 7346 287112 7352
rect 285680 5500 285732 5506
rect 285680 5442 285732 5448
rect 287152 5364 287204 5370
rect 287152 5306 287204 5312
rect 284760 4140 284812 4146
rect 284760 4082 284812 4088
rect 285588 4140 285640 4146
rect 285588 4082 285640 4088
rect 284772 480 284800 4082
rect 285956 3800 286008 3806
rect 285956 3742 286008 3748
rect 285968 480 285996 3742
rect 287164 480 287192 5306
rect 288268 626 288296 337758
rect 288440 335640 288492 335646
rect 288440 335582 288492 335588
rect 288346 16824 288402 16833
rect 288346 16759 288402 16768
rect 288360 16289 288388 16759
rect 288346 16280 288402 16289
rect 288346 16215 288402 16224
rect 288452 7342 288480 335582
rect 288544 10062 288572 340054
rect 289004 336734 289032 340054
rect 288992 336728 289044 336734
rect 288992 336670 289044 336676
rect 289464 335646 289492 340054
rect 289452 335640 289504 335646
rect 289452 335582 289504 335588
rect 288992 318640 289044 318646
rect 288992 318582 289044 318588
rect 289004 308446 289032 318582
rect 288992 308440 289044 308446
rect 288992 308382 289044 308388
rect 288716 290012 288768 290018
rect 288716 289954 288768 289960
rect 288728 289814 288756 289954
rect 288716 289808 288768 289814
rect 288716 289750 288768 289756
rect 288808 289808 288860 289814
rect 288808 289750 288860 289756
rect 288820 280158 288848 289750
rect 288808 280152 288860 280158
rect 288808 280094 288860 280100
rect 288900 280152 288952 280158
rect 288900 280094 288952 280100
rect 288912 269142 288940 280094
rect 288808 269136 288860 269142
rect 288808 269078 288860 269084
rect 288900 269136 288952 269142
rect 288900 269078 288952 269084
rect 288820 258058 288848 269078
rect 288808 258052 288860 258058
rect 288808 257994 288860 258000
rect 288992 258052 289044 258058
rect 288992 257994 289044 258000
rect 289004 248441 289032 257994
rect 288806 248432 288862 248441
rect 288806 248367 288862 248376
rect 288990 248432 289046 248441
rect 288990 248367 289046 248376
rect 288820 230466 288848 248367
rect 288820 230438 288940 230466
rect 288912 222170 288940 230438
rect 288820 222142 288940 222170
rect 288820 211002 288848 222142
rect 288808 210996 288860 211002
rect 288808 210938 288860 210944
rect 289176 210996 289228 211002
rect 289176 210938 289228 210944
rect 289188 201362 289216 210938
rect 288912 201334 289216 201362
rect 288912 190534 288940 201334
rect 288808 190528 288860 190534
rect 288808 190470 288860 190476
rect 288900 190528 288952 190534
rect 288900 190470 288952 190476
rect 288820 190398 288848 190470
rect 288808 190392 288860 190398
rect 288808 190334 288860 190340
rect 288992 190392 289044 190398
rect 288992 190334 289044 190340
rect 289004 180849 289032 190334
rect 288806 180840 288862 180849
rect 288728 180810 288806 180826
rect 288716 180804 288806 180810
rect 288768 180798 288806 180804
rect 288806 180775 288862 180784
rect 288990 180840 289046 180849
rect 288990 180775 289046 180784
rect 288716 180746 288768 180752
rect 289084 177880 289136 177886
rect 289084 177822 289136 177828
rect 289096 169726 289124 177822
rect 289084 169720 289136 169726
rect 289084 169662 289136 169668
rect 289084 160132 289136 160138
rect 289084 160074 289136 160080
rect 289096 155258 289124 160074
rect 288912 155230 289124 155258
rect 288912 150498 288940 155230
rect 288912 150470 289032 150498
rect 289004 150414 289032 150470
rect 288992 150408 289044 150414
rect 288992 150350 289044 150356
rect 288808 140820 288860 140826
rect 288808 140762 288860 140768
rect 288820 131238 288848 140762
rect 288808 131232 288860 131238
rect 288808 131174 288860 131180
rect 288716 131164 288768 131170
rect 288716 131106 288768 131112
rect 288728 126290 288756 131106
rect 288728 126262 289032 126290
rect 289004 104922 289032 126262
rect 288808 104916 288860 104922
rect 288808 104858 288860 104864
rect 288992 104916 289044 104922
rect 288992 104858 289044 104864
rect 288820 102134 288848 104858
rect 288808 102128 288860 102134
rect 288808 102070 288860 102076
rect 288716 92540 288768 92546
rect 288716 92482 288768 92488
rect 288728 84182 288756 92482
rect 288716 84176 288768 84182
rect 288716 84118 288768 84124
rect 288900 75812 288952 75818
rect 288900 75754 288952 75760
rect 288912 48226 288940 75754
rect 288820 48198 288940 48226
rect 288820 45490 288848 48198
rect 288808 45484 288860 45490
rect 288808 45426 288860 45432
rect 289084 45484 289136 45490
rect 289084 45426 289136 45432
rect 289096 44169 289124 45426
rect 288898 44160 288954 44169
rect 288898 44095 288954 44104
rect 289082 44160 289138 44169
rect 289082 44095 289138 44104
rect 288912 35306 288940 44095
rect 288912 35278 289124 35306
rect 289096 29850 289124 35278
rect 289084 29844 289136 29850
rect 289084 29786 289136 29792
rect 288808 19304 288860 19310
rect 288808 19246 288860 19252
rect 288820 12034 288848 19246
rect 289266 16824 289322 16833
rect 289266 16759 289268 16768
rect 289320 16759 289322 16768
rect 289268 16730 289320 16736
rect 288808 12028 288860 12034
rect 288808 11970 288860 11976
rect 288532 10056 288584 10062
rect 288532 9998 288584 10004
rect 289832 9994 289860 340054
rect 290292 331242 290320 340190
rect 290464 337884 290516 337890
rect 290464 337826 290516 337832
rect 290108 331214 290320 331242
rect 290108 313274 290136 331214
rect 290096 313268 290148 313274
rect 290096 313210 290148 313216
rect 290188 306332 290240 306338
rect 290188 306274 290240 306280
rect 290200 303634 290228 306274
rect 290200 303606 290320 303634
rect 290292 284345 290320 303606
rect 290002 284336 290058 284345
rect 290002 284271 290058 284280
rect 290278 284336 290334 284345
rect 290278 284271 290334 284280
rect 290016 277438 290044 284271
rect 290004 277432 290056 277438
rect 290004 277374 290056 277380
rect 290096 277432 290148 277438
rect 290096 277374 290148 277380
rect 290108 258058 290136 277374
rect 290096 258052 290148 258058
rect 290096 257994 290148 258000
rect 290004 248464 290056 248470
rect 290004 248406 290056 248412
rect 290016 245886 290044 248406
rect 290004 245880 290056 245886
rect 290004 245822 290056 245828
rect 290372 245880 290424 245886
rect 290372 245822 290424 245828
rect 290384 220862 290412 245822
rect 290188 220856 290240 220862
rect 290188 220798 290240 220804
rect 290372 220856 290424 220862
rect 290372 220798 290424 220804
rect 290200 212634 290228 220798
rect 290188 212628 290240 212634
rect 290188 212570 290240 212576
rect 290188 212492 290240 212498
rect 290188 212434 290240 212440
rect 290200 196654 290228 212434
rect 290004 196648 290056 196654
rect 290004 196590 290056 196596
rect 290188 196648 290240 196654
rect 290188 196590 290240 196596
rect 290016 172689 290044 196590
rect 290002 172680 290058 172689
rect 290002 172615 290058 172624
rect 290002 172544 290058 172553
rect 290002 172479 290058 172488
rect 290016 154544 290044 172479
rect 290016 154516 290136 154544
rect 290108 131186 290136 154516
rect 290016 131158 290136 131186
rect 290016 122874 290044 131158
rect 290004 122868 290056 122874
rect 290004 122810 290056 122816
rect 290096 122732 290148 122738
rect 290096 122674 290148 122680
rect 290108 102105 290136 122674
rect 290094 102096 290150 102105
rect 290094 102031 290150 102040
rect 289910 101960 289966 101969
rect 289910 101895 289966 101904
rect 289924 84182 289952 101895
rect 289912 84176 289964 84182
rect 289912 84118 289964 84124
rect 290004 74588 290056 74594
rect 290004 74530 290056 74536
rect 290016 57934 290044 74530
rect 290004 57928 290056 57934
rect 290004 57870 290056 57876
rect 290096 57928 290148 57934
rect 290096 57870 290148 57876
rect 290108 45558 290136 57870
rect 290096 45552 290148 45558
rect 290096 45494 290148 45500
rect 290188 45484 290240 45490
rect 290188 45426 290240 45432
rect 290200 22794 290228 45426
rect 290200 22766 290320 22794
rect 289912 16788 289964 16794
rect 289912 16730 289964 16736
rect 289924 16561 289952 16730
rect 289910 16552 289966 16561
rect 289910 16487 289966 16496
rect 290292 12102 290320 22766
rect 290280 12096 290332 12102
rect 290280 12038 290332 12044
rect 289820 9988 289872 9994
rect 289820 9930 289872 9936
rect 288440 7336 288492 7342
rect 288440 7278 288492 7284
rect 289820 6520 289872 6526
rect 289820 6462 289872 6468
rect 288440 6452 288492 6458
rect 288440 6394 288492 6400
rect 288452 3330 288480 6394
rect 288532 6384 288584 6390
rect 288532 6326 288584 6332
rect 288440 3324 288492 3330
rect 288440 3266 288492 3272
rect 288544 3262 288572 6326
rect 289544 3868 289596 3874
rect 289544 3810 289596 3816
rect 288532 3256 288584 3262
rect 288532 3198 288584 3204
rect 288268 598 288388 626
rect 288360 480 288388 598
rect 289556 480 289584 3810
rect 289832 3398 289860 6462
rect 289820 3392 289872 3398
rect 289820 3334 289872 3340
rect 290476 3194 290504 337826
rect 291212 7274 291240 340068
rect 291304 340054 291686 340082
rect 291304 9926 291332 340054
rect 291764 335594 291792 340190
rect 291580 335566 291792 335594
rect 292592 340054 292698 340082
rect 292868 340054 293158 340082
rect 293328 340054 293710 340082
rect 293972 340054 294170 340082
rect 294248 340054 294630 340082
rect 291580 309194 291608 335566
rect 291476 309188 291528 309194
rect 291476 309130 291528 309136
rect 291568 309188 291620 309194
rect 291568 309130 291620 309136
rect 291488 302954 291516 309130
rect 291488 302926 291608 302954
rect 291580 298058 291608 302926
rect 291580 298030 291700 298058
rect 291672 270586 291700 298030
rect 291580 270558 291700 270586
rect 291580 251258 291608 270558
rect 291476 251252 291528 251258
rect 291476 251194 291528 251200
rect 291568 251252 291620 251258
rect 291568 251194 291620 251200
rect 291488 248402 291516 251194
rect 291476 248396 291528 248402
rect 291476 248338 291528 248344
rect 291752 240100 291804 240106
rect 291752 240042 291804 240048
rect 291764 238762 291792 240042
rect 291764 238734 291884 238762
rect 291856 220862 291884 238734
rect 291660 220856 291712 220862
rect 291660 220798 291712 220804
rect 291844 220856 291896 220862
rect 291844 220798 291896 220804
rect 291672 212634 291700 220798
rect 291660 212628 291712 212634
rect 291660 212570 291712 212576
rect 291660 212492 291712 212498
rect 291660 212434 291712 212440
rect 291672 200122 291700 212434
rect 291660 200116 291712 200122
rect 291660 200058 291712 200064
rect 291476 190528 291528 190534
rect 291476 190470 291528 190476
rect 291488 172689 291516 190470
rect 291474 172680 291530 172689
rect 291474 172615 291530 172624
rect 291474 172544 291530 172553
rect 291474 172479 291530 172488
rect 291488 154544 291516 172479
rect 291488 154516 291608 154544
rect 291580 139398 291608 154516
rect 291568 139392 291620 139398
rect 291568 139334 291620 139340
rect 291752 139392 291804 139398
rect 291752 139334 291804 139340
rect 291764 137970 291792 139334
rect 291752 137964 291804 137970
rect 291752 137906 291804 137912
rect 291568 120148 291620 120154
rect 291568 120090 291620 120096
rect 291580 115258 291608 120090
rect 291568 115252 291620 115258
rect 291568 115194 291620 115200
rect 291476 103556 291528 103562
rect 291476 103498 291528 103504
rect 291488 93838 291516 103498
rect 291476 93832 291528 93838
rect 291476 93774 291528 93780
rect 291384 89004 291436 89010
rect 291384 88946 291436 88952
rect 291396 75834 291424 88946
rect 291396 75806 291516 75834
rect 291488 57934 291516 75806
rect 291476 57928 291528 57934
rect 291476 57870 291528 57876
rect 291568 57928 291620 57934
rect 291568 57870 291620 57876
rect 291580 45558 291608 57870
rect 291568 45552 291620 45558
rect 291568 45494 291620 45500
rect 291660 45484 291712 45490
rect 291660 45426 291712 45432
rect 291672 19802 291700 45426
rect 291488 19774 291700 19802
rect 291488 19258 291516 19774
rect 291488 19230 291608 19258
rect 291580 12170 291608 19230
rect 291568 12164 291620 12170
rect 291568 12106 291620 12112
rect 291292 9920 291344 9926
rect 291292 9862 291344 9868
rect 291200 7268 291252 7274
rect 291200 7210 291252 7216
rect 292592 7206 292620 340054
rect 292764 335640 292816 335646
rect 292764 335582 292816 335588
rect 292776 13258 292804 335582
rect 292764 13252 292816 13258
rect 292764 13194 292816 13200
rect 292868 9858 292896 340054
rect 293328 335646 293356 340054
rect 293316 335640 293368 335646
rect 293316 335582 293368 335588
rect 292856 9852 292908 9858
rect 292856 9794 292908 9800
rect 292580 7200 292632 7206
rect 292580 7142 292632 7148
rect 293972 7138 294000 340054
rect 294248 335696 294276 340054
rect 294064 335668 294276 335696
rect 294064 9790 294092 335668
rect 294708 331242 294736 340190
rect 294248 331214 294736 331242
rect 295352 340054 295642 340082
rect 295720 340054 296102 340082
rect 296272 340054 296654 340082
rect 296732 340054 297114 340082
rect 297284 340054 297574 340082
rect 298126 340054 298232 340082
rect 294248 318730 294276 331214
rect 294248 318702 294368 318730
rect 294340 304978 294368 318702
rect 294328 304972 294380 304978
rect 294328 304914 294380 304920
rect 294236 304904 294288 304910
rect 294236 304846 294288 304852
rect 294248 295338 294276 304846
rect 295246 296712 295302 296721
rect 295246 296647 295302 296656
rect 294248 295310 294368 295338
rect 294340 276026 294368 295310
rect 295260 278798 295288 296647
rect 295248 278792 295300 278798
rect 295248 278734 295300 278740
rect 294248 275998 294368 276026
rect 294248 270638 294276 275998
rect 294236 270632 294288 270638
rect 294236 270574 294288 270580
rect 294144 270496 294196 270502
rect 294144 270438 294196 270444
rect 294156 267753 294184 270438
rect 294142 267744 294198 267753
rect 294142 267679 294198 267688
rect 294418 267744 294474 267753
rect 294418 267679 294474 267688
rect 294432 258097 294460 267679
rect 294234 258088 294290 258097
rect 294234 258023 294236 258032
rect 294288 258023 294290 258032
rect 294418 258088 294474 258097
rect 294418 258023 294474 258032
rect 294236 257994 294288 258000
rect 294236 248464 294288 248470
rect 294236 248406 294288 248412
rect 294248 241482 294276 248406
rect 294248 241454 294368 241482
rect 294340 237810 294368 241454
rect 294340 237782 294460 237810
rect 294432 220862 294460 237782
rect 294328 220856 294380 220862
rect 294328 220798 294380 220804
rect 294420 220856 294472 220862
rect 294420 220798 294472 220804
rect 294340 211138 294368 220798
rect 294236 211132 294288 211138
rect 294236 211074 294288 211080
rect 294328 211132 294380 211138
rect 294328 211074 294380 211080
rect 294248 198082 294276 211074
rect 294236 198076 294288 198082
rect 294236 198018 294288 198024
rect 294420 198076 294472 198082
rect 294420 198018 294472 198024
rect 294432 183598 294460 198018
rect 294236 183592 294288 183598
rect 294236 183534 294288 183540
rect 294420 183592 294472 183598
rect 294420 183534 294472 183540
rect 294248 178770 294276 183534
rect 294236 178764 294288 178770
rect 294236 178706 294288 178712
rect 294420 178764 294472 178770
rect 294420 178706 294472 178712
rect 294432 162926 294460 178706
rect 294328 162920 294380 162926
rect 294328 162862 294380 162868
rect 294420 162920 294472 162926
rect 294420 162862 294472 162868
rect 294340 153218 294368 162862
rect 295246 157992 295302 158001
rect 295246 157927 295302 157936
rect 295260 157593 295288 157927
rect 295246 157584 295302 157593
rect 295246 157519 295302 157528
rect 294248 153190 294368 153218
rect 294248 144922 294276 153190
rect 294248 144894 294460 144922
rect 294432 135946 294460 144894
rect 294248 135918 294460 135946
rect 294248 135130 294276 135918
rect 294248 135102 294368 135130
rect 294340 127650 294368 135102
rect 294340 127622 294460 127650
rect 294432 114594 294460 127622
rect 294248 114566 294460 114594
rect 294248 100094 294276 114566
rect 294236 100088 294288 100094
rect 294236 100030 294288 100036
rect 294420 100088 294472 100094
rect 294420 100030 294472 100036
rect 294432 87038 294460 100030
rect 294420 87032 294472 87038
rect 294420 86974 294472 86980
rect 294420 86896 294472 86902
rect 294420 86838 294472 86844
rect 294432 76498 294460 86838
rect 294236 76492 294288 76498
rect 294236 76434 294288 76440
rect 294420 76492 294472 76498
rect 294420 76434 294472 76440
rect 294248 64870 294276 76434
rect 294236 64864 294288 64870
rect 294236 64806 294288 64812
rect 294236 55276 294288 55282
rect 294236 55218 294288 55224
rect 294248 35970 294276 55218
rect 294144 35964 294196 35970
rect 294144 35906 294196 35912
rect 294236 35964 294288 35970
rect 294236 35906 294288 35912
rect 294156 27713 294184 35906
rect 294142 27704 294198 27713
rect 294142 27639 294198 27648
rect 294142 27568 294198 27577
rect 294142 27503 294198 27512
rect 294156 18018 294184 27503
rect 294144 18012 294196 18018
rect 294144 17954 294196 17960
rect 294236 18012 294288 18018
rect 294236 17954 294288 17960
rect 294248 13326 294276 17954
rect 294236 13320 294288 13326
rect 294236 13262 294288 13268
rect 294052 9784 294104 9790
rect 294052 9726 294104 9732
rect 293960 7132 294012 7138
rect 293960 7074 294012 7080
rect 295352 7070 295380 340054
rect 295720 335696 295748 340054
rect 295444 335668 295748 335696
rect 295444 9722 295472 335668
rect 296272 335594 296300 340054
rect 295536 335566 296300 335594
rect 295536 328438 295564 335566
rect 295524 328432 295576 328438
rect 295524 328374 295576 328380
rect 295708 328432 295760 328438
rect 295708 328374 295760 328380
rect 295720 323490 295748 328374
rect 295628 323462 295748 323490
rect 295628 298246 295656 323462
rect 295616 298240 295668 298246
rect 295616 298182 295668 298188
rect 295524 298036 295576 298042
rect 295524 297978 295576 297984
rect 295536 296721 295564 297978
rect 295522 296712 295578 296721
rect 295522 296647 295578 296656
rect 295524 278792 295576 278798
rect 295524 278734 295576 278740
rect 295536 277914 295564 278734
rect 295524 277908 295576 277914
rect 295524 277850 295576 277856
rect 295800 277908 295852 277914
rect 295800 277850 295852 277856
rect 295812 264330 295840 277850
rect 295720 264302 295840 264330
rect 295720 251190 295748 264302
rect 295524 251184 295576 251190
rect 295524 251126 295576 251132
rect 295708 251184 295760 251190
rect 295708 251126 295760 251132
rect 295536 241482 295564 251126
rect 295536 241454 295656 241482
rect 295536 222222 295564 222253
rect 295628 222222 295656 241454
rect 295524 222216 295576 222222
rect 295616 222216 295668 222222
rect 295576 222164 295616 222170
rect 295524 222158 295668 222164
rect 295536 222142 295656 222158
rect 295536 202910 295564 202941
rect 295628 202910 295656 222142
rect 295524 202904 295576 202910
rect 295616 202904 295668 202910
rect 295576 202852 295616 202858
rect 295524 202846 295668 202852
rect 295536 202830 295656 202846
rect 295628 186454 295656 202830
rect 295616 186448 295668 186454
rect 295616 186390 295668 186396
rect 295524 186312 295576 186318
rect 295524 186254 295576 186260
rect 295536 178770 295564 186254
rect 295524 178764 295576 178770
rect 295524 178706 295576 178712
rect 295708 178764 295760 178770
rect 295708 178706 295760 178712
rect 295720 157418 295748 178706
rect 295524 157412 295576 157418
rect 295524 157354 295576 157360
rect 295708 157412 295760 157418
rect 295708 157354 295760 157360
rect 295536 144922 295564 157354
rect 295536 144894 295748 144922
rect 295720 140758 295748 144894
rect 295708 140752 295760 140758
rect 295708 140694 295760 140700
rect 295616 131164 295668 131170
rect 295616 131106 295668 131112
rect 295628 127650 295656 131106
rect 295628 127622 295748 127650
rect 295720 114594 295748 127622
rect 295536 114566 295748 114594
rect 295536 104854 295564 114566
rect 295524 104848 295576 104854
rect 295524 104790 295576 104796
rect 295616 104848 295668 104854
rect 295616 104790 295668 104796
rect 295628 91746 295656 104790
rect 295628 91718 295748 91746
rect 295720 80730 295748 91718
rect 295536 80702 295748 80730
rect 295536 28966 295564 80702
rect 296534 76256 296590 76265
rect 296534 76191 296590 76200
rect 296548 75857 296576 76191
rect 296534 75848 296590 75857
rect 296534 75783 296590 75792
rect 295524 28960 295576 28966
rect 295524 28902 295576 28908
rect 295616 28960 295668 28966
rect 295616 28902 295668 28908
rect 295628 12510 295656 28902
rect 295616 12504 295668 12510
rect 295616 12446 295668 12452
rect 295432 9716 295484 9722
rect 295432 9658 295484 9664
rect 295340 7064 295392 7070
rect 295340 7006 295392 7012
rect 296732 6730 296760 340054
rect 297284 335696 297312 340054
rect 297916 337204 297968 337210
rect 297916 337146 297968 337152
rect 296824 335668 297312 335696
rect 296824 328438 296852 335668
rect 296812 328432 296864 328438
rect 296812 328374 296864 328380
rect 296996 328432 297048 328438
rect 296996 328374 297048 328380
rect 297008 323490 297036 328374
rect 296916 323462 297036 323490
rect 296916 296750 296944 323462
rect 296812 296744 296864 296750
rect 296812 296686 296864 296692
rect 296904 296744 296956 296750
rect 296904 296686 296956 296692
rect 296824 277438 296852 296686
rect 296812 277432 296864 277438
rect 296812 277374 296864 277380
rect 297088 277432 297140 277438
rect 297088 277374 297140 277380
rect 297100 259486 297128 277374
rect 296996 259480 297048 259486
rect 296996 259422 297048 259428
rect 297088 259480 297140 259486
rect 297088 259422 297140 259428
rect 297008 258058 297036 259422
rect 296996 258052 297048 258058
rect 296996 257994 297048 258000
rect 297180 258052 297232 258058
rect 297180 257994 297232 258000
rect 297192 248441 297220 257994
rect 296902 248432 296958 248441
rect 296902 248367 296958 248376
rect 297178 248432 297234 248441
rect 297178 248367 297234 248376
rect 296824 222222 296852 222253
rect 296916 222222 296944 248367
rect 296812 222216 296864 222222
rect 296904 222216 296956 222222
rect 296864 222164 296904 222170
rect 296812 222158 296956 222164
rect 296824 222142 296944 222158
rect 296824 202910 296852 202941
rect 296916 202910 296944 222142
rect 296812 202904 296864 202910
rect 296904 202904 296956 202910
rect 296864 202852 296904 202858
rect 296812 202846 296956 202852
rect 296824 202830 296944 202846
rect 296916 186454 296944 202830
rect 296904 186448 296956 186454
rect 296904 186390 296956 186396
rect 296812 186312 296864 186318
rect 296812 186254 296864 186260
rect 296824 172530 296852 186254
rect 296824 172514 296944 172530
rect 296824 172508 296956 172514
rect 296824 172502 296904 172508
rect 296904 172450 296956 172456
rect 296996 172508 297048 172514
rect 296996 172450 297048 172456
rect 296916 172419 296944 172450
rect 297008 157418 297036 172450
rect 296812 157412 296864 157418
rect 296812 157354 296864 157360
rect 296996 157412 297048 157418
rect 296996 157354 297048 157360
rect 296824 144922 296852 157354
rect 296824 144894 297036 144922
rect 297008 142118 297036 144894
rect 296996 142112 297048 142118
rect 296996 142054 297048 142060
rect 296904 132524 296956 132530
rect 296904 132466 296956 132472
rect 296916 122874 296944 132466
rect 296904 122868 296956 122874
rect 296904 122810 296956 122816
rect 297088 122868 297140 122874
rect 297088 122810 297140 122816
rect 297100 113218 297128 122810
rect 296996 113212 297048 113218
rect 296996 113154 297048 113160
rect 297088 113212 297140 113218
rect 297088 113154 297140 113160
rect 297008 108338 297036 113154
rect 296824 108310 297036 108338
rect 296824 93809 296852 108310
rect 296810 93800 296866 93809
rect 296810 93735 296866 93744
rect 297178 93664 297234 93673
rect 297178 93599 297234 93608
rect 297192 85490 297220 93599
rect 297546 87136 297602 87145
rect 297546 87071 297548 87080
rect 297600 87071 297602 87080
rect 297548 87042 297600 87048
rect 297008 85462 297220 85490
rect 297008 84182 297036 85462
rect 296996 84176 297048 84182
rect 296996 84118 297048 84124
rect 296904 74588 296956 74594
rect 296904 74530 296956 74536
rect 296916 74458 296944 74530
rect 296904 74452 296956 74458
rect 296904 74394 296956 74400
rect 296812 64932 296864 64938
rect 296812 64874 296864 64880
rect 296824 45558 296852 64874
rect 296812 45552 296864 45558
rect 296812 45494 296864 45500
rect 296812 38616 296864 38622
rect 296812 38558 296864 38564
rect 296824 29186 296852 38558
rect 296824 29158 296944 29186
rect 296916 13394 296944 29158
rect 296904 13388 296956 13394
rect 296904 13330 296956 13336
rect 296720 6724 296772 6730
rect 296720 6666 296772 6672
rect 297364 6724 297416 6730
rect 297364 6666 297416 6672
rect 295892 6588 295944 6594
rect 295892 6530 295944 6536
rect 294328 6316 294380 6322
rect 294328 6258 294380 6264
rect 290740 5432 290792 5438
rect 290740 5374 290792 5380
rect 290464 3188 290516 3194
rect 290464 3130 290516 3136
rect 290752 480 290780 5374
rect 291936 3256 291988 3262
rect 291936 3198 291988 3204
rect 291948 480 291976 3198
rect 293132 3052 293184 3058
rect 293132 2994 293184 3000
rect 293144 480 293172 2994
rect 294340 480 294368 6258
rect 295904 4146 295932 6530
rect 295892 4140 295944 4146
rect 295892 4082 295944 4088
rect 296720 4140 296772 4146
rect 296720 4082 296772 4088
rect 295524 3120 295576 3126
rect 295524 3062 295576 3068
rect 295536 480 295564 3062
rect 296732 480 296760 4082
rect 297376 4010 297404 6666
rect 297824 5500 297876 5506
rect 297824 5442 297876 5448
rect 297836 4026 297864 5442
rect 297928 4146 297956 337146
rect 298006 157584 298062 157593
rect 298006 157519 298008 157528
rect 298060 157519 298062 157528
rect 298008 157490 298060 157496
rect 298006 29472 298062 29481
rect 298006 29407 298062 29416
rect 298020 29209 298048 29407
rect 298006 29200 298062 29209
rect 298006 29135 298062 29144
rect 298100 16584 298152 16590
rect 298098 16552 298100 16561
rect 298152 16552 298154 16561
rect 298098 16487 298154 16496
rect 298204 12306 298232 340054
rect 298388 340054 298586 340082
rect 298664 340054 299046 340082
rect 298284 335640 298336 335646
rect 298284 335582 298336 335588
rect 298296 13462 298324 335582
rect 298284 13456 298336 13462
rect 298284 13398 298336 13404
rect 298192 12300 298244 12306
rect 298192 12242 298244 12248
rect 298388 6798 298416 340054
rect 298664 335646 298692 340054
rect 298652 335640 298704 335646
rect 298652 335582 298704 335588
rect 299584 331362 299612 340068
rect 299768 340054 300058 340082
rect 300228 340054 300518 340082
rect 300964 340054 301070 340082
rect 301240 340054 301530 340082
rect 301700 340054 301990 340082
rect 302344 340054 302542 340082
rect 302712 340054 303002 340082
rect 303080 340054 303462 340082
rect 303724 340054 303922 340082
rect 304184 340054 304474 340082
rect 304644 340054 304934 340082
rect 305104 340054 305394 340082
rect 305656 340054 305946 340082
rect 299572 331356 299624 331362
rect 299572 331298 299624 331304
rect 299768 331242 299796 340054
rect 299676 331214 299796 331242
rect 299572 331084 299624 331090
rect 299572 331026 299624 331032
rect 299480 331016 299532 331022
rect 299480 330958 299532 330964
rect 299492 241466 299520 330958
rect 299480 241460 299532 241466
rect 299480 241402 299532 241408
rect 299480 231872 299532 231878
rect 299480 231814 299532 231820
rect 299492 222154 299520 231814
rect 299480 222148 299532 222154
rect 299480 222090 299532 222096
rect 299480 212560 299532 212566
rect 299480 212502 299532 212508
rect 299492 202842 299520 212502
rect 299480 202836 299532 202842
rect 299480 202778 299532 202784
rect 299480 193248 299532 193254
rect 299480 193190 299532 193196
rect 298466 17096 298522 17105
rect 298466 17031 298522 17040
rect 298480 16590 298508 17031
rect 298468 16584 298520 16590
rect 298468 16526 298520 16532
rect 299492 6866 299520 193190
rect 299584 12374 299612 331026
rect 299676 331022 299704 331214
rect 299664 331016 299716 331022
rect 299664 330958 299716 330964
rect 300228 318850 300256 340054
rect 300860 335640 300912 335646
rect 300860 335582 300912 335588
rect 299848 318844 299900 318850
rect 299848 318786 299900 318792
rect 300216 318844 300268 318850
rect 300216 318786 300268 318792
rect 299860 317422 299888 318786
rect 299848 317416 299900 317422
rect 299848 317358 299900 317364
rect 299848 299532 299900 299538
rect 299848 299474 299900 299480
rect 299860 296682 299888 299474
rect 299848 296676 299900 296682
rect 299848 296618 299900 296624
rect 299940 296676 299992 296682
rect 299940 296618 299992 296624
rect 299952 277409 299980 296618
rect 299662 277400 299718 277409
rect 299662 277335 299718 277344
rect 299938 277400 299994 277409
rect 299938 277335 299994 277344
rect 299676 267782 299704 277335
rect 299664 267776 299716 267782
rect 299664 267718 299716 267724
rect 299848 267776 299900 267782
rect 299848 267718 299900 267724
rect 299860 259418 299888 267718
rect 299848 259412 299900 259418
rect 299848 259354 299900 259360
rect 300032 259412 300084 259418
rect 300032 259354 300084 259360
rect 299952 240174 299980 240205
rect 300044 240174 300072 259354
rect 299940 240168 299992 240174
rect 299860 240116 299940 240122
rect 299860 240110 299992 240116
rect 300032 240168 300084 240174
rect 300032 240110 300084 240116
rect 299860 240094 299980 240110
rect 299860 222306 299888 240094
rect 299860 222278 299980 222306
rect 299952 212548 299980 222278
rect 299860 212520 299980 212548
rect 299860 202994 299888 212520
rect 299860 202966 299980 202994
rect 299952 193338 299980 202966
rect 299952 193310 300072 193338
rect 300044 191842 300072 193310
rect 299860 191814 300072 191842
rect 299860 188494 299888 191814
rect 299848 188488 299900 188494
rect 299848 188430 299900 188436
rect 299848 183592 299900 183598
rect 299848 183534 299900 183540
rect 299860 182170 299888 183534
rect 299848 182164 299900 182170
rect 299848 182106 299900 182112
rect 299940 182164 299992 182170
rect 299940 182106 299992 182112
rect 299952 159390 299980 182106
rect 299756 159384 299808 159390
rect 299756 159326 299808 159332
rect 299940 159384 299992 159390
rect 299940 159326 299992 159332
rect 299768 144922 299796 159326
rect 299768 144894 299888 144922
rect 299860 132818 299888 144894
rect 299768 132790 299888 132818
rect 299768 132530 299796 132790
rect 299756 132524 299808 132530
rect 299756 132466 299808 132472
rect 299848 132524 299900 132530
rect 299848 132466 299900 132472
rect 299860 118794 299888 132466
rect 299848 118788 299900 118794
rect 299848 118730 299900 118736
rect 299848 118652 299900 118658
rect 299848 118594 299900 118600
rect 299860 113150 299888 118594
rect 299848 113144 299900 113150
rect 299848 113086 299900 113092
rect 299940 113144 299992 113150
rect 299940 113086 299992 113092
rect 299952 85610 299980 113086
rect 299848 85604 299900 85610
rect 299848 85546 299900 85552
rect 299940 85604 299992 85610
rect 299940 85546 299992 85552
rect 299860 77314 299888 85546
rect 299756 77308 299808 77314
rect 299756 77250 299808 77256
rect 299848 77308 299900 77314
rect 299848 77250 299900 77256
rect 299768 71074 299796 77250
rect 299768 71046 299980 71074
rect 299952 67538 299980 71046
rect 299860 67510 299980 67538
rect 299860 58002 299888 67510
rect 299756 57996 299808 58002
rect 299756 57938 299808 57944
rect 299848 57996 299900 58002
rect 299848 57938 299900 57944
rect 299768 42090 299796 57938
rect 299756 42084 299808 42090
rect 299756 42026 299808 42032
rect 300124 42084 300176 42090
rect 300124 42026 300176 42032
rect 300136 29322 300164 42026
rect 299952 29294 300164 29322
rect 299952 27606 299980 29294
rect 299756 27600 299808 27606
rect 299756 27542 299808 27548
rect 299940 27600 299992 27606
rect 299940 27542 299992 27548
rect 299768 26246 299796 27542
rect 299756 26240 299808 26246
rect 299756 26182 299808 26188
rect 299756 16652 299808 16658
rect 299756 16594 299808 16600
rect 299768 13530 299796 16594
rect 299756 13524 299808 13530
rect 299756 13466 299808 13472
rect 299572 12368 299624 12374
rect 299572 12310 299624 12316
rect 299480 6860 299532 6866
rect 299480 6802 299532 6808
rect 298376 6792 298428 6798
rect 298376 6734 298428 6740
rect 298100 6656 298152 6662
rect 298100 6598 298152 6604
rect 297916 4140 297968 4146
rect 297916 4082 297968 4088
rect 298112 4078 298140 6598
rect 300872 6118 300900 335582
rect 300964 12442 300992 340054
rect 301240 335646 301268 340054
rect 301228 335640 301280 335646
rect 301228 335582 301280 335588
rect 301700 330546 301728 340054
rect 302240 335708 302292 335714
rect 302240 335650 302292 335656
rect 301136 330540 301188 330546
rect 301136 330482 301188 330488
rect 301688 330540 301740 330546
rect 301688 330482 301740 330488
rect 301148 325689 301176 330482
rect 301134 325680 301190 325689
rect 301134 325615 301190 325624
rect 301318 325680 301374 325689
rect 301318 325615 301374 325624
rect 301332 316062 301360 325615
rect 301136 316056 301188 316062
rect 301136 315998 301188 316004
rect 301320 316056 301372 316062
rect 301320 315998 301372 316004
rect 301148 307834 301176 315998
rect 301136 307828 301188 307834
rect 301136 307770 301188 307776
rect 301228 307692 301280 307698
rect 301228 307634 301280 307640
rect 301240 306377 301268 307634
rect 301226 306368 301282 306377
rect 301226 306303 301282 306312
rect 301410 306368 301466 306377
rect 301410 306303 301466 306312
rect 301424 296750 301452 306303
rect 301044 296744 301096 296750
rect 301042 296712 301044 296721
rect 301412 296744 301464 296750
rect 301096 296712 301098 296721
rect 301412 296686 301464 296692
rect 301042 296647 301098 296656
rect 301134 296576 301190 296585
rect 301134 296511 301190 296520
rect 301148 283778 301176 296511
rect 301148 283750 301268 283778
rect 301240 278798 301268 283750
rect 301044 278792 301096 278798
rect 301044 278734 301096 278740
rect 301228 278792 301280 278798
rect 301228 278734 301280 278740
rect 301056 273290 301084 278734
rect 301044 273284 301096 273290
rect 301044 273226 301096 273232
rect 301136 273216 301188 273222
rect 301136 273158 301188 273164
rect 301148 270502 301176 273158
rect 301136 270496 301188 270502
rect 301136 270438 301188 270444
rect 301228 270496 301280 270502
rect 301228 270438 301280 270444
rect 301240 246242 301268 270438
rect 301056 246214 301268 246242
rect 301056 241505 301084 246214
rect 301042 241496 301098 241505
rect 301042 241431 301098 241440
rect 301134 241360 301190 241369
rect 301134 241295 301190 241304
rect 301148 231946 301176 241295
rect 301136 231940 301188 231946
rect 301136 231882 301188 231888
rect 301044 231804 301096 231810
rect 301044 231746 301096 231752
rect 301056 222193 301084 231746
rect 301042 222184 301098 222193
rect 301042 222119 301098 222128
rect 301134 222048 301190 222057
rect 301134 221983 301190 221992
rect 301148 212634 301176 221983
rect 301136 212628 301188 212634
rect 301136 212570 301188 212576
rect 301044 212492 301096 212498
rect 301044 212434 301096 212440
rect 301056 202881 301084 212434
rect 301042 202872 301098 202881
rect 301042 202807 301098 202816
rect 301134 202736 301190 202745
rect 301134 202671 301190 202680
rect 301148 196602 301176 202671
rect 301148 196574 301268 196602
rect 301240 183598 301268 196574
rect 301044 183592 301096 183598
rect 301044 183534 301096 183540
rect 301228 183592 301280 183598
rect 301228 183534 301280 183540
rect 301056 176730 301084 183534
rect 301044 176724 301096 176730
rect 301044 176666 301096 176672
rect 301136 176588 301188 176594
rect 301136 176530 301188 176536
rect 301148 169266 301176 176530
rect 301148 169238 301268 169266
rect 301240 164257 301268 169238
rect 301042 164248 301098 164257
rect 301042 164183 301098 164192
rect 301226 164248 301282 164257
rect 301226 164183 301282 164192
rect 301056 154494 301084 164183
rect 301044 154488 301096 154494
rect 301044 154430 301096 154436
rect 301228 154488 301280 154494
rect 301228 154430 301280 154436
rect 301240 144945 301268 154430
rect 301042 144936 301098 144945
rect 301042 144871 301098 144880
rect 301226 144936 301282 144945
rect 301226 144871 301282 144880
rect 301056 138038 301084 144871
rect 301044 138032 301096 138038
rect 301044 137974 301096 137980
rect 301136 137964 301188 137970
rect 301136 137906 301188 137912
rect 301148 130506 301176 137906
rect 301148 130478 301268 130506
rect 301240 125633 301268 130478
rect 301042 125624 301098 125633
rect 301042 125559 301098 125568
rect 301226 125624 301282 125633
rect 301226 125559 301282 125568
rect 301056 113286 301084 125559
rect 301044 113280 301096 113286
rect 301044 113222 301096 113228
rect 301136 113212 301188 113218
rect 301136 113154 301188 113160
rect 301148 85610 301176 113154
rect 301136 85604 301188 85610
rect 301136 85546 301188 85552
rect 301228 85604 301280 85610
rect 301228 85546 301280 85552
rect 301240 77382 301268 85546
rect 301228 77376 301280 77382
rect 301228 77318 301280 77324
rect 301228 75880 301280 75886
rect 301228 75822 301280 75828
rect 301240 66298 301268 75822
rect 301044 66292 301096 66298
rect 301044 66234 301096 66240
rect 301228 66292 301280 66298
rect 301228 66234 301280 66240
rect 301056 57934 301084 66234
rect 301044 57928 301096 57934
rect 301044 57870 301096 57876
rect 301044 51808 301096 51814
rect 301044 51750 301096 51756
rect 301056 46918 301084 51750
rect 301044 46912 301096 46918
rect 301044 46854 301096 46860
rect 301320 46912 301372 46918
rect 301320 46854 301372 46860
rect 301332 45558 301360 46854
rect 301320 45552 301372 45558
rect 301320 45494 301372 45500
rect 301320 35964 301372 35970
rect 301320 35906 301372 35912
rect 301332 29016 301360 35906
rect 301332 28988 301452 29016
rect 301424 28778 301452 28988
rect 301240 28750 301452 28778
rect 301240 27606 301268 28750
rect 301136 27600 301188 27606
rect 301136 27542 301188 27548
rect 301228 27600 301280 27606
rect 301228 27542 301280 27548
rect 301148 13598 301176 27542
rect 301136 13592 301188 13598
rect 301136 13534 301188 13540
rect 300952 12436 301004 12442
rect 300952 12378 301004 12384
rect 300860 6112 300912 6118
rect 300860 6054 300912 6060
rect 302252 6050 302280 335650
rect 302344 11694 302372 340054
rect 302712 335714 302740 340054
rect 302700 335708 302752 335714
rect 302700 335650 302752 335656
rect 303080 334762 303108 340054
rect 303160 337952 303212 337958
rect 303160 337894 303212 337900
rect 302608 334756 302660 334762
rect 302608 334698 302660 334704
rect 303068 334756 303120 334762
rect 303068 334698 303120 334704
rect 302620 328438 302648 334698
rect 303172 334642 303200 337894
rect 303620 335640 303672 335646
rect 303620 335582 303672 335588
rect 302896 334614 303200 334642
rect 302608 328432 302660 328438
rect 302608 328374 302660 328380
rect 302608 318844 302660 318850
rect 302608 318786 302660 318792
rect 302620 311982 302648 318786
rect 302608 311976 302660 311982
rect 302608 311918 302660 311924
rect 302516 311840 302568 311846
rect 302516 311782 302568 311788
rect 302528 299538 302556 311782
rect 302516 299532 302568 299538
rect 302516 299474 302568 299480
rect 302608 299532 302660 299538
rect 302608 299474 302660 299480
rect 302620 296682 302648 299474
rect 302608 296676 302660 296682
rect 302608 296618 302660 296624
rect 302700 296676 302752 296682
rect 302700 296618 302752 296624
rect 302712 270586 302740 296618
rect 302620 270558 302740 270586
rect 302620 249801 302648 270558
rect 302422 249792 302478 249801
rect 302422 249727 302478 249736
rect 302606 249792 302662 249801
rect 302606 249727 302662 249736
rect 302436 240174 302464 249727
rect 302424 240168 302476 240174
rect 302424 240110 302476 240116
rect 302700 240168 302752 240174
rect 302700 240110 302752 240116
rect 302712 232014 302740 240110
rect 302700 232008 302752 232014
rect 302700 231950 302752 231956
rect 302608 230512 302660 230518
rect 302608 230454 302660 230460
rect 302620 222306 302648 230454
rect 302620 222278 302740 222306
rect 302712 212650 302740 222278
rect 302712 212622 302832 212650
rect 302804 212378 302832 212622
rect 302620 212350 302832 212378
rect 302620 202994 302648 212350
rect 302620 202966 302740 202994
rect 302712 193322 302740 202966
rect 302700 193316 302752 193322
rect 302700 193258 302752 193264
rect 302516 193180 302568 193186
rect 302516 193122 302568 193128
rect 302528 183666 302556 193122
rect 302516 183660 302568 183666
rect 302516 183602 302568 183608
rect 302608 183592 302660 183598
rect 302608 183534 302660 183540
rect 302620 176798 302648 183534
rect 302608 176792 302660 176798
rect 302608 176734 302660 176740
rect 302516 176656 302568 176662
rect 302516 176598 302568 176604
rect 302528 169590 302556 176598
rect 302516 169584 302568 169590
rect 302516 169526 302568 169532
rect 302792 169584 302844 169590
rect 302792 169526 302844 169532
rect 302804 162897 302832 169526
rect 302606 162888 302662 162897
rect 302606 162823 302608 162832
rect 302660 162823 302662 162832
rect 302790 162888 302846 162897
rect 302790 162823 302846 162832
rect 302608 162794 302660 162800
rect 302516 153264 302568 153270
rect 302516 153206 302568 153212
rect 302528 153134 302556 153206
rect 302516 153128 302568 153134
rect 302516 153070 302568 153076
rect 302792 153128 302844 153134
rect 302792 153070 302844 153076
rect 302804 143585 302832 153070
rect 302606 143576 302662 143585
rect 302424 143540 302476 143546
rect 302606 143511 302608 143520
rect 302424 143482 302476 143488
rect 302660 143511 302662 143520
rect 302790 143576 302846 143585
rect 302790 143511 302846 143520
rect 302608 143482 302660 143488
rect 302436 132530 302464 143482
rect 302424 132524 302476 132530
rect 302424 132466 302476 132472
rect 302608 132524 302660 132530
rect 302608 132466 302660 132472
rect 302620 104854 302648 132466
rect 302608 104848 302660 104854
rect 302608 104790 302660 104796
rect 302608 95260 302660 95266
rect 302608 95202 302660 95208
rect 302620 77314 302648 95202
rect 302516 77308 302568 77314
rect 302516 77250 302568 77256
rect 302608 77308 302660 77314
rect 302608 77250 302660 77256
rect 302528 67726 302556 77250
rect 302516 67720 302568 67726
rect 302516 67662 302568 67668
rect 302424 67652 302476 67658
rect 302424 67594 302476 67600
rect 302436 58002 302464 67594
rect 302424 57996 302476 58002
rect 302424 57938 302476 57944
rect 302516 57996 302568 58002
rect 302516 57938 302568 57944
rect 302528 46918 302556 57938
rect 302516 46912 302568 46918
rect 302516 46854 302568 46860
rect 302608 46912 302660 46918
rect 302608 46854 302660 46860
rect 302620 19378 302648 46854
rect 302790 29064 302846 29073
rect 302790 28999 302846 29008
rect 302804 28801 302832 28999
rect 302790 28792 302846 28801
rect 302790 28727 302846 28736
rect 302516 19372 302568 19378
rect 302516 19314 302568 19320
rect 302608 19372 302660 19378
rect 302608 19314 302660 19320
rect 302528 13666 302556 19314
rect 302516 13660 302568 13666
rect 302516 13602 302568 13608
rect 302332 11688 302384 11694
rect 302332 11630 302384 11636
rect 302240 6044 302292 6050
rect 302240 5986 302292 5992
rect 301412 4412 301464 4418
rect 301412 4354 301464 4360
rect 300308 4140 300360 4146
rect 300308 4082 300360 4088
rect 298100 4072 298152 4078
rect 297364 4004 297416 4010
rect 297836 3998 297956 4026
rect 298100 4014 298152 4020
rect 297364 3946 297416 3952
rect 297928 480 297956 3998
rect 299112 3392 299164 3398
rect 299112 3334 299164 3340
rect 299124 480 299152 3334
rect 300320 480 300348 4082
rect 301424 480 301452 4354
rect 302608 4072 302660 4078
rect 302608 4014 302660 4020
rect 302620 480 302648 4014
rect 302896 3398 302924 334614
rect 303632 5982 303660 335582
rect 303724 11626 303752 340054
rect 304184 335646 304212 340054
rect 304172 335640 304224 335646
rect 304172 335582 304224 335588
rect 304644 328506 304672 340054
rect 305000 335640 305052 335646
rect 305000 335582 305052 335588
rect 303896 328500 303948 328506
rect 303896 328442 303948 328448
rect 304632 328500 304684 328506
rect 304632 328442 304684 328448
rect 303908 311930 303936 328442
rect 303816 311902 303936 311930
rect 303816 311794 303844 311902
rect 303816 311766 303936 311794
rect 303908 292618 303936 311766
rect 303816 292590 303936 292618
rect 303816 292482 303844 292590
rect 303816 292454 303936 292482
rect 303908 176746 303936 292454
rect 303816 176718 303936 176746
rect 303816 176610 303844 176718
rect 303816 176582 303936 176610
rect 303908 138122 303936 176582
rect 303816 138094 303936 138122
rect 303816 137986 303844 138094
rect 303816 137958 303936 137986
rect 303908 118810 303936 137958
rect 303816 118782 303936 118810
rect 303816 118674 303844 118782
rect 303816 118646 303936 118674
rect 303908 80102 303936 118646
rect 303896 80096 303948 80102
rect 303896 80038 303948 80044
rect 303896 79960 303948 79966
rect 303896 79902 303948 79908
rect 303908 77246 303936 79902
rect 303896 77240 303948 77246
rect 303896 77182 303948 77188
rect 303988 77240 304040 77246
rect 303988 77182 304040 77188
rect 304000 58002 304028 77182
rect 303896 57996 303948 58002
rect 303896 57938 303948 57944
rect 303988 57996 304040 58002
rect 303988 57938 304040 57944
rect 303908 51762 303936 57938
rect 303816 51734 303936 51762
rect 303816 40186 303844 51734
rect 303804 40180 303856 40186
rect 303804 40122 303856 40128
rect 303896 32428 303948 32434
rect 303896 32370 303948 32376
rect 303908 13802 303936 32370
rect 303896 13796 303948 13802
rect 303896 13738 303948 13744
rect 303712 11620 303764 11626
rect 303712 11562 303764 11568
rect 303620 5976 303672 5982
rect 303620 5918 303672 5924
rect 305012 5914 305040 335582
rect 305104 11558 305132 340054
rect 305656 335646 305684 340054
rect 306196 338020 306248 338026
rect 306196 337962 306248 337968
rect 305644 335640 305696 335646
rect 305644 335582 305696 335588
rect 305092 11552 305144 11558
rect 305092 11494 305144 11500
rect 305000 5908 305052 5914
rect 305000 5850 305052 5856
rect 305000 4344 305052 4350
rect 305000 4286 305052 4292
rect 302884 3392 302936 3398
rect 302884 3334 302936 3340
rect 303804 3324 303856 3330
rect 303804 3266 303856 3272
rect 303816 480 303844 3266
rect 305012 480 305040 4286
rect 306208 480 306236 337962
rect 306392 333418 306420 340068
rect 306668 340054 306866 340082
rect 307036 340054 307418 340082
rect 307878 340054 307984 340082
rect 306392 333390 306604 333418
rect 306472 331084 306524 331090
rect 306472 331026 306524 331032
rect 306288 157548 306340 157554
rect 306288 157490 306340 157496
rect 306300 157457 306328 157490
rect 306286 157448 306342 157457
rect 306286 157383 306342 157392
rect 306288 87100 306340 87106
rect 306288 87042 306340 87048
rect 306300 87009 306328 87042
rect 306286 87000 306342 87009
rect 306286 86935 306342 86944
rect 306378 75984 306434 75993
rect 306378 75919 306380 75928
rect 306432 75919 306434 75928
rect 306380 75890 306432 75896
rect 306378 40216 306434 40225
rect 306378 40151 306380 40160
rect 306432 40151 306434 40160
rect 306380 40122 306432 40128
rect 306380 28824 306432 28830
rect 306378 28792 306380 28801
rect 306432 28792 306434 28801
rect 306378 28727 306434 28736
rect 306378 17096 306434 17105
rect 306378 17031 306380 17040
rect 306432 17031 306434 17040
rect 306380 17002 306432 17008
rect 306484 11490 306512 331026
rect 306576 13734 306604 333390
rect 306668 331090 306696 340054
rect 307036 331242 307064 340054
rect 307760 337748 307812 337754
rect 307760 337690 307812 337696
rect 307772 337657 307800 337690
rect 307758 337648 307814 337657
rect 307758 337583 307814 337592
rect 307760 335640 307812 335646
rect 307760 335582 307812 335588
rect 306760 331214 307064 331242
rect 306656 331084 306708 331090
rect 306656 331026 306708 331032
rect 306760 317490 306788 331214
rect 306748 317484 306800 317490
rect 306748 317426 306800 317432
rect 306748 316056 306800 316062
rect 306748 315998 306800 316004
rect 306760 307834 306788 315998
rect 306748 307828 306800 307834
rect 306748 307770 306800 307776
rect 306932 307692 306984 307698
rect 306932 307634 306984 307640
rect 306944 306354 306972 307634
rect 306852 306326 306972 306354
rect 306852 299538 306880 306326
rect 306840 299532 306892 299538
rect 306840 299474 306892 299480
rect 306840 296744 306892 296750
rect 306840 296686 306892 296692
rect 306852 292670 306880 296686
rect 306840 292664 306892 292670
rect 306840 292606 306892 292612
rect 306748 292528 306800 292534
rect 306748 292470 306800 292476
rect 306760 287065 306788 292470
rect 306746 287056 306802 287065
rect 306746 286991 306802 287000
rect 307022 287056 307078 287065
rect 307022 286991 307078 287000
rect 307036 277506 307064 286991
rect 307024 277500 307076 277506
rect 307024 277442 307076 277448
rect 306840 277432 306892 277438
rect 306840 277374 306892 277380
rect 306852 262954 306880 277374
rect 306840 262948 306892 262954
rect 306840 262890 306892 262896
rect 306932 249824 306984 249830
rect 306930 249792 306932 249801
rect 306984 249792 306986 249801
rect 306930 249727 306986 249736
rect 307114 249792 307170 249801
rect 307114 249727 307170 249736
rect 307128 240174 307156 249727
rect 306932 240168 306984 240174
rect 306932 240110 306984 240116
rect 307116 240168 307168 240174
rect 307116 240110 307168 240116
rect 306944 231878 306972 240110
rect 306932 231872 306984 231878
rect 306932 231814 306984 231820
rect 306748 231804 306800 231810
rect 306748 231746 306800 231752
rect 306760 222222 306788 231746
rect 306748 222216 306800 222222
rect 306748 222158 306800 222164
rect 306932 222216 306984 222222
rect 306932 222158 306984 222164
rect 306944 212634 306972 222158
rect 306932 212628 306984 212634
rect 306932 212570 306984 212576
rect 306748 212492 306800 212498
rect 306748 212434 306800 212440
rect 306760 202910 306788 212434
rect 306748 202904 306800 202910
rect 306748 202846 306800 202852
rect 306932 202904 306984 202910
rect 306932 202846 306984 202852
rect 306944 193338 306972 202846
rect 306944 193310 307064 193338
rect 307036 191842 307064 193310
rect 306852 191814 307064 191842
rect 306852 188494 306880 191814
rect 306840 188488 306892 188494
rect 306840 188430 306892 188436
rect 306840 183592 306892 183598
rect 306840 183534 306892 183540
rect 306852 176798 306880 183534
rect 306840 176792 306892 176798
rect 306840 176734 306892 176740
rect 306748 176656 306800 176662
rect 306748 176598 306800 176604
rect 306760 169590 306788 176598
rect 306748 169584 306800 169590
rect 306748 169526 306800 169532
rect 307024 169584 307076 169590
rect 307024 169526 307076 169532
rect 307036 162897 307064 169526
rect 306838 162888 306894 162897
rect 306748 162852 306800 162858
rect 306838 162823 306840 162832
rect 306748 162794 306800 162800
rect 306892 162823 306894 162832
rect 307022 162888 307078 162897
rect 307022 162823 307078 162832
rect 306840 162794 306892 162800
rect 306760 149546 306788 162794
rect 307576 157480 307628 157486
rect 307574 157448 307576 157457
rect 307628 157448 307630 157457
rect 307574 157383 307630 157392
rect 306760 149518 306880 149546
rect 306852 138122 306880 149518
rect 306852 138094 306972 138122
rect 306944 137850 306972 138094
rect 306760 137822 306972 137850
rect 306760 132462 306788 137822
rect 306748 132456 306800 132462
rect 306748 132398 306800 132404
rect 306840 129940 306892 129946
rect 306840 129882 306892 129888
rect 306852 121446 306880 129882
rect 306840 121440 306892 121446
rect 306840 121382 306892 121388
rect 306840 111852 306892 111858
rect 306840 111794 306892 111800
rect 306852 92614 306880 111794
rect 306840 92608 306892 92614
rect 306840 92550 306892 92556
rect 306748 92540 306800 92546
rect 306748 92482 306800 92488
rect 306760 85610 306788 92482
rect 306748 85604 306800 85610
rect 306748 85546 306800 85552
rect 306840 85604 306892 85610
rect 306840 85546 306892 85552
rect 306852 84182 306880 85546
rect 306840 84176 306892 84182
rect 306840 84118 306892 84124
rect 306748 75812 306800 75818
rect 306748 75754 306800 75760
rect 306760 66298 306788 75754
rect 306656 66292 306708 66298
rect 306656 66234 306708 66240
rect 306748 66292 306800 66298
rect 306748 66234 306800 66240
rect 306668 60042 306696 66234
rect 306656 60036 306708 60042
rect 306656 59978 306708 59984
rect 307024 52012 307076 52018
rect 307024 51954 307076 51960
rect 307036 45558 307064 51954
rect 307024 45552 307076 45558
rect 307024 45494 307076 45500
rect 307024 35964 307076 35970
rect 307024 35906 307076 35912
rect 307036 30546 307064 35906
rect 306944 30518 307064 30546
rect 306944 27606 306972 30518
rect 306932 27600 306984 27606
rect 306932 27542 306984 27548
rect 306840 27532 306892 27538
rect 306840 27474 306892 27480
rect 306852 19258 306880 27474
rect 306852 19230 306972 19258
rect 306564 13728 306616 13734
rect 306564 13670 306616 13676
rect 306472 11484 306524 11490
rect 306472 11426 306524 11432
rect 306944 9722 306972 19230
rect 307574 16552 307630 16561
rect 307574 16487 307630 16496
rect 307588 11286 307616 16487
rect 307576 11280 307628 11286
rect 307576 11222 307628 11228
rect 306656 9716 306708 9722
rect 306656 9658 306708 9664
rect 306932 9716 306984 9722
rect 306932 9658 306984 9664
rect 306668 5846 306696 9658
rect 306656 5840 306708 5846
rect 306656 5782 306708 5788
rect 307772 5778 307800 335582
rect 307956 13054 307984 340054
rect 308048 340054 308338 340082
rect 308600 340054 308890 340082
rect 309244 340054 309350 340082
rect 309428 340054 309810 340082
rect 310072 340054 310362 340082
rect 310624 340054 310822 340082
rect 311084 340054 311282 340082
rect 311544 340054 311834 340082
rect 312004 340054 312294 340082
rect 307944 13048 307996 13054
rect 307944 12990 307996 12996
rect 308048 11422 308076 340054
rect 308600 335646 308628 340054
rect 308588 335640 308640 335646
rect 308588 335582 308640 335588
rect 309140 335640 309192 335646
rect 309140 335582 309192 335588
rect 308036 11416 308088 11422
rect 308036 11358 308088 11364
rect 307760 5772 307812 5778
rect 307760 5714 307812 5720
rect 309152 5710 309180 335582
rect 309244 9450 309272 340054
rect 309428 11354 309456 340054
rect 309784 337340 309836 337346
rect 309784 337282 309836 337288
rect 309416 11348 309468 11354
rect 309416 11290 309468 11296
rect 309232 9444 309284 9450
rect 309232 9386 309284 9392
rect 309140 5704 309192 5710
rect 309140 5646 309192 5652
rect 308588 4276 308640 4282
rect 308588 4218 308640 4224
rect 307390 3360 307446 3369
rect 307390 3295 307446 3304
rect 307404 480 307432 3295
rect 308600 480 308628 4218
rect 309796 4078 309824 337282
rect 310072 335646 310100 340054
rect 310060 335640 310112 335646
rect 310060 335582 310112 335588
rect 310520 332104 310572 332110
rect 310520 332046 310572 332052
rect 310532 5642 310560 332046
rect 310624 9518 310652 340054
rect 311084 331242 311112 340054
rect 311544 332110 311572 340054
rect 311532 332104 311584 332110
rect 311532 332046 311584 332052
rect 310808 331214 311112 331242
rect 310808 321638 310836 331214
rect 310796 321632 310848 321638
rect 310796 321574 310848 321580
rect 310888 321496 310940 321502
rect 310888 321438 310940 321444
rect 310900 311982 310928 321438
rect 310888 311976 310940 311982
rect 310888 311918 310940 311924
rect 310704 307896 310756 307902
rect 310704 307838 310756 307844
rect 310716 307766 310744 307838
rect 310704 307760 310756 307766
rect 310704 307702 310756 307708
rect 310888 298172 310940 298178
rect 310888 298114 310940 298120
rect 310900 293078 310928 298114
rect 310888 293072 310940 293078
rect 310888 293014 310940 293020
rect 310888 282804 310940 282810
rect 310888 282746 310940 282752
rect 310900 278730 310928 282746
rect 310888 278724 310940 278730
rect 310888 278666 310940 278672
rect 310888 263492 310940 263498
rect 310888 263434 310940 263440
rect 310900 256086 310928 263434
rect 310888 256080 310940 256086
rect 310888 256022 310940 256028
rect 310704 251320 310756 251326
rect 310704 251262 310756 251268
rect 310716 251190 310744 251262
rect 310704 251184 310756 251190
rect 310704 251126 310756 251132
rect 310888 241528 310940 241534
rect 310888 241470 310940 241476
rect 310900 234734 310928 241470
rect 310888 234728 310940 234734
rect 310888 234670 310940 234676
rect 310796 234592 310848 234598
rect 310796 234534 310848 234540
rect 310808 231810 310836 234534
rect 310796 231804 310848 231810
rect 310796 231746 310848 231752
rect 310888 222216 310940 222222
rect 310888 222158 310940 222164
rect 310900 215422 310928 222158
rect 310888 215416 310940 215422
rect 310888 215358 310940 215364
rect 310796 215280 310848 215286
rect 310796 215222 310848 215228
rect 310808 212498 310836 215222
rect 310796 212492 310848 212498
rect 310796 212434 310848 212440
rect 310888 202904 310940 202910
rect 310888 202846 310940 202852
rect 310900 196110 310928 202846
rect 310888 196104 310940 196110
rect 310888 196046 310940 196052
rect 310796 195968 310848 195974
rect 310796 195910 310848 195916
rect 310808 193225 310836 195910
rect 310794 193216 310850 193225
rect 310794 193151 310850 193160
rect 311070 193216 311126 193225
rect 311070 193151 311126 193160
rect 311084 183598 311112 193151
rect 310888 183592 310940 183598
rect 310888 183534 310940 183540
rect 311072 183592 311124 183598
rect 311072 183534 311124 183540
rect 310900 176798 310928 183534
rect 310888 176792 310940 176798
rect 310888 176734 310940 176740
rect 310796 176656 310848 176662
rect 310796 176598 310848 176604
rect 310808 167074 310836 176598
rect 310796 167068 310848 167074
rect 310796 167010 310848 167016
rect 310888 166932 310940 166938
rect 310888 166874 310940 166880
rect 310900 153377 310928 166874
rect 310886 153368 310942 153377
rect 310886 153303 310942 153312
rect 310794 153232 310850 153241
rect 310794 153167 310796 153176
rect 310848 153167 310850 153176
rect 310796 153138 310848 153144
rect 310796 147620 310848 147626
rect 310796 147562 310848 147568
rect 310808 143562 310836 147562
rect 310808 143534 310928 143562
rect 310900 138718 310928 143534
rect 310888 138712 310940 138718
rect 310888 138654 310940 138660
rect 310796 128308 310848 128314
rect 310796 128250 310848 128256
rect 310808 125610 310836 128250
rect 310808 125582 310928 125610
rect 310900 125526 310928 125582
rect 310888 125520 310940 125526
rect 310888 125462 310940 125468
rect 310888 114640 310940 114646
rect 310808 114588 310888 114594
rect 310808 114582 310940 114588
rect 310808 114566 310928 114582
rect 310808 114510 310836 114566
rect 310796 114504 310848 114510
rect 310796 114446 310848 114452
rect 310888 104916 310940 104922
rect 310888 104858 310940 104864
rect 310900 99482 310928 104858
rect 310888 99476 310940 99482
rect 310888 99418 310940 99424
rect 310888 99340 310940 99346
rect 310888 99282 310940 99288
rect 310900 95282 310928 99282
rect 310808 95254 310928 95282
rect 310808 95198 310836 95254
rect 310796 95192 310848 95198
rect 310796 95134 310848 95140
rect 310796 85604 310848 85610
rect 310796 85546 310848 85552
rect 310808 76242 310836 85546
rect 310808 76214 310928 76242
rect 310900 75970 310928 76214
rect 310808 75942 310928 75970
rect 311254 75984 311310 75993
rect 310808 75886 310836 75942
rect 311254 75919 311256 75928
rect 311308 75919 311310 75928
rect 311256 75890 311308 75896
rect 310796 75880 310848 75886
rect 310796 75822 310848 75828
rect 310796 66360 310848 66366
rect 310796 66302 310848 66308
rect 310808 66230 310836 66302
rect 310796 66224 310848 66230
rect 310796 66166 310848 66172
rect 311072 60036 311124 60042
rect 311072 59978 311124 59984
rect 311084 45694 311112 59978
rect 310888 45688 310940 45694
rect 310888 45630 310940 45636
rect 311072 45688 311124 45694
rect 311072 45630 311124 45636
rect 310900 45558 310928 45630
rect 310888 45552 310940 45558
rect 310888 45494 310940 45500
rect 311072 45552 311124 45558
rect 311072 45494 311124 45500
rect 311084 27690 311112 45494
rect 310900 27662 311112 27690
rect 310900 22114 310928 27662
rect 310900 22086 311020 22114
rect 310992 16726 311020 22086
rect 310980 16720 311032 16726
rect 310980 16662 311032 16668
rect 310796 16652 310848 16658
rect 310796 16594 310848 16600
rect 310808 16561 310836 16594
rect 310794 16552 310850 16561
rect 310794 16487 310850 16496
rect 312004 9586 312032 340054
rect 312544 337272 312596 337278
rect 312544 337214 312596 337220
rect 311992 9580 312044 9586
rect 311992 9522 312044 9528
rect 310612 9512 310664 9518
rect 310612 9454 310664 9460
rect 310520 5636 310572 5642
rect 310520 5578 310572 5584
rect 312176 4208 312228 4214
rect 312176 4150 312228 4156
rect 309784 4072 309836 4078
rect 309784 4014 309836 4020
rect 310980 3392 311032 3398
rect 310980 3334 311032 3340
rect 309784 3188 309836 3194
rect 309784 3130 309836 3136
rect 309796 480 309824 3130
rect 310992 480 311020 3334
rect 312188 480 312216 4150
rect 312556 3058 312584 337214
rect 312740 337142 312768 340068
rect 312728 337136 312780 337142
rect 312728 337078 312780 337084
rect 313292 5574 313320 340068
rect 313384 340054 313766 340082
rect 313384 9654 313412 340054
rect 314212 337210 314240 340068
rect 314778 340054 314884 340082
rect 314660 338088 314712 338094
rect 314660 338030 314712 338036
rect 314200 337204 314252 337210
rect 314200 337146 314252 337152
rect 313372 9648 313424 9654
rect 313372 9590 313424 9596
rect 313280 5568 313332 5574
rect 313280 5510 313332 5516
rect 314672 4865 314700 338030
rect 314856 12986 314884 340054
rect 314948 340054 315238 340082
rect 315408 340054 315698 340082
rect 314844 12980 314896 12986
rect 314844 12922 314896 12928
rect 314948 8906 314976 340054
rect 315408 338094 315436 340054
rect 316132 338156 316184 338162
rect 316132 338098 316184 338104
rect 315396 338088 315448 338094
rect 315396 338030 315448 338036
rect 316040 337340 316092 337346
rect 316040 337282 316092 337288
rect 315948 157480 316000 157486
rect 315946 157448 315948 157457
rect 316000 157448 316002 157457
rect 315946 157383 316002 157392
rect 315948 40180 316000 40186
rect 315948 40122 316000 40128
rect 315960 40089 315988 40122
rect 315946 40080 316002 40089
rect 315946 40015 316002 40024
rect 315946 28928 316002 28937
rect 315946 28863 316002 28872
rect 315960 28830 315988 28863
rect 315948 28824 316000 28830
rect 315948 28766 316000 28772
rect 315948 17060 316000 17066
rect 315948 17002 316000 17008
rect 315960 16697 315988 17002
rect 315946 16688 316002 16697
rect 315946 16623 316002 16632
rect 314936 8900 314988 8906
rect 314936 8842 314988 8848
rect 314658 4856 314714 4865
rect 314658 4791 314714 4800
rect 316052 4758 316080 337282
rect 316144 8838 316172 338098
rect 316236 12918 316264 340068
rect 316328 340054 316710 340082
rect 316880 340054 317170 340082
rect 317616 340054 317722 340082
rect 317892 340054 318182 340082
rect 318352 340054 318642 340082
rect 318996 340054 319194 340082
rect 319272 340054 319654 340082
rect 319824 340054 320114 340082
rect 320284 340054 320666 340082
rect 320744 340054 321126 340082
rect 316328 338162 316356 340054
rect 316316 338156 316368 338162
rect 316316 338098 316368 338104
rect 316880 337346 316908 340054
rect 317328 337748 317380 337754
rect 317328 337690 317380 337696
rect 317340 337657 317368 337690
rect 317326 337648 317382 337657
rect 317326 337583 317382 337592
rect 316868 337340 316920 337346
rect 316868 337282 316920 337288
rect 317420 337340 317472 337346
rect 317420 337282 317472 337288
rect 316684 337136 316736 337142
rect 316684 337078 316736 337084
rect 316224 12912 316276 12918
rect 316224 12854 316276 12860
rect 316132 8832 316184 8838
rect 316132 8774 316184 8780
rect 316040 4752 316092 4758
rect 316040 4694 316092 4700
rect 313372 4072 313424 4078
rect 313372 4014 313424 4020
rect 312544 3052 312596 3058
rect 312544 2994 312596 3000
rect 313384 480 313412 4014
rect 314568 4004 314620 4010
rect 314568 3946 314620 3952
rect 314580 480 314608 3946
rect 316696 3262 316724 337078
rect 317326 157720 317382 157729
rect 317326 157655 317382 157664
rect 317340 157457 317368 157655
rect 317326 157448 317382 157457
rect 317326 157383 317382 157392
rect 317326 29336 317382 29345
rect 317326 29271 317382 29280
rect 317340 28937 317368 29271
rect 317326 28928 317382 28937
rect 317326 28863 317382 28872
rect 317432 4690 317460 337282
rect 317512 306400 317564 306406
rect 317512 306342 317564 306348
rect 317524 219434 317552 306342
rect 317512 219428 317564 219434
rect 317512 219370 317564 219376
rect 317512 209840 317564 209846
rect 317512 209782 317564 209788
rect 317524 200122 317552 209782
rect 317512 200116 317564 200122
rect 317512 200058 317564 200064
rect 317512 190528 317564 190534
rect 317512 190470 317564 190476
rect 317524 180810 317552 190470
rect 317512 180804 317564 180810
rect 317512 180746 317564 180752
rect 317512 142180 317564 142186
rect 317512 142122 317564 142128
rect 317524 137970 317552 142122
rect 317512 137964 317564 137970
rect 317512 137906 317564 137912
rect 317512 55276 317564 55282
rect 317512 55218 317564 55224
rect 317524 45558 317552 55218
rect 317512 45552 317564 45558
rect 317512 45494 317564 45500
rect 317512 31816 317564 31822
rect 317512 31758 317564 31764
rect 317524 8770 317552 31758
rect 317616 12850 317644 340054
rect 317892 337770 317920 340054
rect 317708 337742 317920 337770
rect 317708 306406 317736 337742
rect 318352 337346 318380 340054
rect 318800 338156 318852 338162
rect 318800 338098 318852 338104
rect 318340 337340 318392 337346
rect 318340 337282 318392 337288
rect 317696 306400 317748 306406
rect 317696 306342 317748 306348
rect 317696 219428 317748 219434
rect 317696 219370 317748 219376
rect 317708 209846 317736 219370
rect 317696 209840 317748 209846
rect 317696 209782 317748 209788
rect 317696 200116 317748 200122
rect 317696 200058 317748 200064
rect 317708 190534 317736 200058
rect 317696 190528 317748 190534
rect 317696 190470 317748 190476
rect 317696 180804 317748 180810
rect 317696 180746 317748 180752
rect 317708 142186 317736 180746
rect 317696 142180 317748 142186
rect 317696 142122 317748 142128
rect 317788 137964 317840 137970
rect 317788 137906 317840 137912
rect 317800 128330 317828 137906
rect 317708 128302 317828 128330
rect 317708 99770 317736 128302
rect 317708 99742 317828 99770
rect 317800 89758 317828 99742
rect 317788 89752 317840 89758
rect 317788 89694 317840 89700
rect 317880 89616 317932 89622
rect 317880 89558 317932 89564
rect 317892 85542 317920 89558
rect 317880 85536 317932 85542
rect 317880 85478 317932 85484
rect 317696 75948 317748 75954
rect 317696 75890 317748 75896
rect 317708 55282 317736 75890
rect 317696 55276 317748 55282
rect 317696 55218 317748 55224
rect 317696 45552 317748 45558
rect 317696 45494 317748 45500
rect 317708 31822 317736 45494
rect 317696 31816 317748 31822
rect 317696 31758 317748 31764
rect 317604 12844 317656 12850
rect 317604 12786 317656 12792
rect 317512 8764 317564 8770
rect 317512 8706 317564 8712
rect 318708 4752 318760 4758
rect 318708 4694 318760 4700
rect 317420 4684 317472 4690
rect 317420 4626 317472 4632
rect 318720 3466 318748 4694
rect 318812 4622 318840 338098
rect 318892 337340 318944 337346
rect 318892 337282 318944 337288
rect 318904 8702 318932 337282
rect 318996 12782 319024 340054
rect 319272 337346 319300 340054
rect 319824 338162 319852 340054
rect 319812 338156 319864 338162
rect 319812 338098 319864 338104
rect 319260 337340 319312 337346
rect 319260 337282 319312 337288
rect 320180 337340 320232 337346
rect 320180 337282 320232 337288
rect 319444 337000 319496 337006
rect 319444 336942 319496 336948
rect 318984 12776 319036 12782
rect 318984 12718 319036 12724
rect 318892 8696 318944 8702
rect 318892 8638 318944 8644
rect 318800 4616 318852 4622
rect 318800 4558 318852 4564
rect 318708 3460 318760 3466
rect 318708 3402 318760 3408
rect 316684 3256 316736 3262
rect 316684 3198 316736 3204
rect 318064 3256 318116 3262
rect 318064 3198 318116 3204
rect 315764 3052 315816 3058
rect 315764 2994 315816 3000
rect 315776 480 315804 2994
rect 316960 2984 317012 2990
rect 316960 2926 317012 2932
rect 316972 480 317000 2926
rect 318076 480 318104 3198
rect 319456 3126 319484 336942
rect 320192 8634 320220 337282
rect 320284 12714 320312 340054
rect 320744 337346 320772 340054
rect 320732 337340 320784 337346
rect 320732 337282 320784 337288
rect 321468 337204 321520 337210
rect 321468 337146 321520 337152
rect 320272 12708 320324 12714
rect 320272 12650 320324 12656
rect 320180 8628 320232 8634
rect 320180 8570 320232 8576
rect 321480 4808 321508 337146
rect 321204 4780 321508 4808
rect 320364 4548 320416 4554
rect 320364 4490 320416 4496
rect 320376 3534 320404 4490
rect 321204 3534 321232 4780
rect 321572 4706 321600 340068
rect 321756 340054 322138 340082
rect 322216 340054 322598 340082
rect 322952 340054 323058 340082
rect 323136 340054 323518 340082
rect 323688 340054 324070 340082
rect 324332 340054 324530 340082
rect 324700 340054 324990 340082
rect 325160 340054 325542 340082
rect 325712 340054 326002 340082
rect 326080 340054 326462 340082
rect 321652 335640 321704 335646
rect 321652 335582 321704 335588
rect 321664 8566 321692 335582
rect 321756 12646 321784 340054
rect 322216 335646 322244 340054
rect 322204 335640 322256 335646
rect 322204 335582 322256 335588
rect 321744 12640 321796 12646
rect 321744 12582 321796 12588
rect 321652 8560 321704 8566
rect 321652 8502 321704 8508
rect 321652 5092 321704 5098
rect 321652 5034 321704 5040
rect 321664 4962 321692 5034
rect 321652 4956 321704 4962
rect 321652 4898 321704 4904
rect 321388 4678 321600 4706
rect 321388 4622 321416 4678
rect 321376 4616 321428 4622
rect 321376 4558 321428 4564
rect 322756 4616 322808 4622
rect 322756 4558 322808 4564
rect 320364 3528 320416 3534
rect 320364 3470 320416 3476
rect 320456 3528 320508 3534
rect 320456 3470 320508 3476
rect 321192 3528 321244 3534
rect 321192 3470 321244 3476
rect 321652 3528 321704 3534
rect 321652 3470 321704 3476
rect 319444 3120 319496 3126
rect 319444 3062 319496 3068
rect 319260 2916 319312 2922
rect 319260 2858 319312 2864
rect 319272 480 319300 2858
rect 320468 480 320496 3470
rect 321664 480 321692 3470
rect 322768 3466 322796 4558
rect 322952 4486 322980 340054
rect 323032 85604 323084 85610
rect 323032 85546 323084 85552
rect 323044 75954 323072 85546
rect 323032 75948 323084 75954
rect 323032 75890 323084 75896
rect 323136 12578 323164 340054
rect 323688 328506 323716 340054
rect 323308 328500 323360 328506
rect 323308 328442 323360 328448
rect 323676 328500 323728 328506
rect 323676 328442 323728 328448
rect 323320 311982 323348 328442
rect 323308 311976 323360 311982
rect 323308 311918 323360 311924
rect 323216 311908 323268 311914
rect 323216 311850 323268 311856
rect 323228 304314 323256 311850
rect 323228 304286 323440 304314
rect 323412 302138 323440 304286
rect 323320 302110 323440 302138
rect 323320 299470 323348 302110
rect 323308 299464 323360 299470
rect 323308 299406 323360 299412
rect 323492 288448 323544 288454
rect 323492 288390 323544 288396
rect 323504 282826 323532 288390
rect 323412 282798 323532 282826
rect 323412 280158 323440 282798
rect 323308 280152 323360 280158
rect 323308 280094 323360 280100
rect 323400 280152 323452 280158
rect 323400 280094 323452 280100
rect 323320 273986 323348 280094
rect 323320 273958 323440 273986
rect 323412 252754 323440 273958
rect 323400 252748 323452 252754
rect 323400 252690 323452 252696
rect 323400 241528 323452 241534
rect 323400 241470 323452 241476
rect 323412 234734 323440 241470
rect 323400 234728 323452 234734
rect 323400 234670 323452 234676
rect 323400 231804 323452 231810
rect 323400 231746 323452 231752
rect 323412 217546 323440 231746
rect 323412 217518 323532 217546
rect 323504 211177 323532 217518
rect 323306 211168 323362 211177
rect 323306 211103 323362 211112
rect 323490 211168 323546 211177
rect 323490 211103 323546 211112
rect 323320 205698 323348 211103
rect 323308 205692 323360 205698
rect 323308 205634 323360 205640
rect 323400 205556 323452 205562
rect 323400 205498 323452 205504
rect 323412 198098 323440 205498
rect 323412 198070 323532 198098
rect 323504 193254 323532 198070
rect 323308 193248 323360 193254
rect 323306 193216 323308 193225
rect 323492 193248 323544 193254
rect 323360 193216 323362 193225
rect 323306 193151 323362 193160
rect 323490 193216 323492 193225
rect 323544 193216 323546 193225
rect 323490 193151 323546 193160
rect 323504 186266 323532 193151
rect 323412 186238 323532 186266
rect 323412 178786 323440 186238
rect 323412 178758 323532 178786
rect 323504 173942 323532 178758
rect 323308 173936 323360 173942
rect 323308 173878 323360 173884
rect 323492 173936 323544 173942
rect 323492 173878 323544 173884
rect 323320 169402 323348 173878
rect 323320 169374 323440 169402
rect 323412 157570 323440 169374
rect 323412 157542 323532 157570
rect 323504 155394 323532 157542
rect 323412 155366 323532 155394
rect 323412 144906 323440 155366
rect 323308 144900 323360 144906
rect 323308 144842 323360 144848
rect 323400 144900 323452 144906
rect 323400 144842 323452 144848
rect 323320 143546 323348 144842
rect 323308 143540 323360 143546
rect 323308 143482 323360 143488
rect 323492 143540 323544 143546
rect 323492 143482 323544 143488
rect 323504 128330 323532 143482
rect 323412 128302 323532 128330
rect 323412 125594 323440 128302
rect 323216 125588 323268 125594
rect 323216 125530 323268 125536
rect 323400 125588 323452 125594
rect 323400 125530 323452 125536
rect 323228 118674 323256 125530
rect 323228 118646 323348 118674
rect 323320 109698 323348 118646
rect 323320 109670 323532 109698
rect 323504 106162 323532 109670
rect 323412 106134 323532 106162
rect 323412 104854 323440 106134
rect 323400 104848 323452 104854
rect 323400 104790 323452 104796
rect 323400 95260 323452 95266
rect 323400 95202 323452 95208
rect 323412 85610 323440 95202
rect 323400 85604 323452 85610
rect 323400 85546 323452 85552
rect 323308 75948 323360 75954
rect 323308 75890 323360 75896
rect 323320 61470 323348 75890
rect 323308 61464 323360 61470
rect 323308 61406 323360 61412
rect 323308 48340 323360 48346
rect 323308 48282 323360 48288
rect 323320 38690 323348 48282
rect 323308 38684 323360 38690
rect 323308 38626 323360 38632
rect 323400 38548 323452 38554
rect 323400 38490 323452 38496
rect 323412 28966 323440 38490
rect 323308 28960 323360 28966
rect 323308 28902 323360 28908
rect 323400 28960 323452 28966
rect 323400 28902 323452 28908
rect 323124 12572 323176 12578
rect 323124 12514 323176 12520
rect 323320 8498 323348 28902
rect 323308 8492 323360 8498
rect 323308 8434 323360 8440
rect 324332 4894 324360 340054
rect 324700 335730 324728 340054
rect 324424 335702 324728 335730
rect 324424 7614 324452 335702
rect 325160 328506 325188 340054
rect 324688 328500 324740 328506
rect 324688 328442 324740 328448
rect 325148 328500 325200 328506
rect 325148 328442 325200 328448
rect 324700 311930 324728 328442
rect 324608 311902 324728 311930
rect 324608 304314 324636 311902
rect 324516 304286 324636 304314
rect 324516 302138 324544 304286
rect 324516 302110 324728 302138
rect 324700 299470 324728 302110
rect 324688 299464 324740 299470
rect 324688 299406 324740 299412
rect 324688 289876 324740 289882
rect 324688 289818 324740 289824
rect 324700 282962 324728 289818
rect 324700 282934 324820 282962
rect 324792 282826 324820 282934
rect 324608 282798 324820 282826
rect 324608 280106 324636 282798
rect 324516 280078 324636 280106
rect 324516 278730 324544 280078
rect 324504 278724 324556 278730
rect 324504 278666 324556 278672
rect 324596 269136 324648 269142
rect 324596 269078 324648 269084
rect 324608 260846 324636 269078
rect 324596 260840 324648 260846
rect 324596 260782 324648 260788
rect 324688 260772 324740 260778
rect 324688 260714 324740 260720
rect 324700 249898 324728 260714
rect 324596 249892 324648 249898
rect 324596 249834 324648 249840
rect 324688 249892 324740 249898
rect 324688 249834 324740 249840
rect 324608 240174 324636 249834
rect 324596 240168 324648 240174
rect 324596 240110 324648 240116
rect 324688 240168 324740 240174
rect 324688 240110 324740 240116
rect 324700 239986 324728 240110
rect 324608 239958 324728 239986
rect 324608 231810 324636 239958
rect 324596 231804 324648 231810
rect 324596 231746 324648 231752
rect 324780 231804 324832 231810
rect 324780 231746 324832 231752
rect 324792 212566 324820 231746
rect 324688 212560 324740 212566
rect 324688 212502 324740 212508
rect 324780 212560 324832 212566
rect 324780 212502 324832 212508
rect 324700 202910 324728 212502
rect 324596 202904 324648 202910
rect 324596 202846 324648 202852
rect 324688 202904 324740 202910
rect 324688 202846 324740 202852
rect 324608 193254 324636 202846
rect 324596 193248 324648 193254
rect 324596 193190 324648 193196
rect 324688 193248 324740 193254
rect 324688 193190 324740 193196
rect 324700 191826 324728 193190
rect 324688 191820 324740 191826
rect 324688 191762 324740 191768
rect 324872 191820 324924 191826
rect 324872 191762 324924 191768
rect 324884 182209 324912 191762
rect 324594 182200 324650 182209
rect 324594 182135 324650 182144
rect 324870 182200 324926 182209
rect 324870 182135 324926 182144
rect 324608 172530 324636 182135
rect 324608 172514 324728 172530
rect 324608 172508 324740 172514
rect 324608 172502 324688 172508
rect 324688 172450 324740 172456
rect 324700 172419 324728 172450
rect 324596 162920 324648 162926
rect 324596 162862 324648 162868
rect 324608 157570 324636 162862
rect 324516 157542 324636 157570
rect 324516 157298 324544 157542
rect 324516 157270 324636 157298
rect 324608 144906 324636 157270
rect 324596 144900 324648 144906
rect 324596 144842 324648 144848
rect 324780 144900 324832 144906
rect 324780 144842 324832 144848
rect 324792 139890 324820 144842
rect 324700 139862 324820 139890
rect 324700 135250 324728 139862
rect 324596 135244 324648 135250
rect 324596 135186 324648 135192
rect 324688 135244 324740 135250
rect 324688 135186 324740 135192
rect 324608 125594 324636 135186
rect 324596 125588 324648 125594
rect 324596 125530 324648 125536
rect 324780 125588 324832 125594
rect 324780 125530 324832 125536
rect 324792 120630 324820 125530
rect 324780 120624 324832 120630
rect 324780 120566 324832 120572
rect 324596 113212 324648 113218
rect 324596 113154 324648 113160
rect 324608 109750 324636 113154
rect 324596 109744 324648 109750
rect 324596 109686 324648 109692
rect 324596 109608 324648 109614
rect 324596 109550 324648 109556
rect 324608 104854 324636 109550
rect 324596 104848 324648 104854
rect 324596 104790 324648 104796
rect 324596 95260 324648 95266
rect 324596 95202 324648 95208
rect 324608 86970 324636 95202
rect 324596 86964 324648 86970
rect 324596 86906 324648 86912
rect 324688 86896 324740 86902
rect 324688 86838 324740 86844
rect 324700 66314 324728 86838
rect 324700 66286 324912 66314
rect 324884 64870 324912 66286
rect 324872 64864 324924 64870
rect 324872 64806 324924 64812
rect 324964 64864 325016 64870
rect 324964 64806 325016 64812
rect 324976 48226 325004 64806
rect 324700 48198 325004 48226
rect 324700 28966 324728 48198
rect 324596 28960 324648 28966
rect 324596 28902 324648 28908
rect 324688 28960 324740 28966
rect 324688 28902 324740 28908
rect 324608 8430 324636 28902
rect 324596 8424 324648 8430
rect 324596 8366 324648 8372
rect 324412 7608 324464 7614
rect 324412 7550 324464 7556
rect 324320 4888 324372 4894
rect 324320 4830 324372 4836
rect 325712 4826 325740 340054
rect 326080 335594 326108 340054
rect 325804 335566 326108 335594
rect 325804 7682 325832 335566
rect 326540 333334 326568 340190
rect 327092 340054 327474 340082
rect 327644 340054 327934 340082
rect 328486 340054 328684 340082
rect 325976 333328 326028 333334
rect 325976 333270 326028 333276
rect 326528 333328 326580 333334
rect 326528 333270 326580 333276
rect 325988 317422 326016 333270
rect 325976 317416 326028 317422
rect 325976 317358 326028 317364
rect 325884 307828 325936 307834
rect 325884 307770 325936 307776
rect 325896 299470 325924 307770
rect 325884 299464 325936 299470
rect 325884 299406 325936 299412
rect 325976 299396 326028 299402
rect 325976 299338 326028 299344
rect 325988 298110 326016 299338
rect 325976 298104 326028 298110
rect 325976 298046 326028 298052
rect 325976 288448 326028 288454
rect 325976 288390 326028 288396
rect 325988 263702 326016 288390
rect 325976 263696 326028 263702
rect 325976 263638 326028 263644
rect 325884 263560 325936 263566
rect 325884 263502 325936 263508
rect 325896 251190 325924 263502
rect 325884 251184 325936 251190
rect 325884 251126 325936 251132
rect 325884 249824 325936 249830
rect 325882 249792 325884 249801
rect 325936 249792 325938 249801
rect 325882 249727 325938 249736
rect 326158 249792 326214 249801
rect 326158 249727 326214 249736
rect 326172 240174 326200 249727
rect 325976 240168 326028 240174
rect 325976 240110 326028 240116
rect 326160 240168 326212 240174
rect 326160 240110 326212 240116
rect 325988 227338 326016 240110
rect 325988 227310 326108 227338
rect 326080 220862 326108 227310
rect 325884 220856 325936 220862
rect 325884 220798 325936 220804
rect 326068 220856 326120 220862
rect 326068 220798 326120 220804
rect 325896 212566 325924 220798
rect 325884 212560 325936 212566
rect 325884 212502 325936 212508
rect 325976 212560 326028 212566
rect 325976 212502 326028 212508
rect 325988 202910 326016 212502
rect 325884 202904 325936 202910
rect 325882 202872 325884 202881
rect 325976 202904 326028 202910
rect 325936 202872 325938 202881
rect 325976 202846 326028 202852
rect 325882 202807 325938 202816
rect 325974 202736 326030 202745
rect 325974 202671 326030 202680
rect 325988 186454 326016 202671
rect 325976 186448 326028 186454
rect 325976 186390 326028 186396
rect 325884 186312 325936 186318
rect 325884 186254 325936 186260
rect 325896 173942 325924 186254
rect 325884 173936 325936 173942
rect 325884 173878 325936 173884
rect 325976 173936 326028 173942
rect 325976 173878 326028 173884
rect 325988 164234 326016 173878
rect 325896 164206 326016 164234
rect 325896 162840 325924 164206
rect 325896 162812 326016 162840
rect 325988 157282 326016 162812
rect 325976 157276 326028 157282
rect 325976 157218 326028 157224
rect 325976 157140 326028 157146
rect 325976 157082 326028 157088
rect 325988 149818 326016 157082
rect 325988 149790 326108 149818
rect 326080 144945 326108 149790
rect 325882 144936 325938 144945
rect 325882 144871 325884 144880
rect 325936 144871 325938 144880
rect 326066 144936 326122 144945
rect 326066 144871 326068 144880
rect 325884 144842 325936 144848
rect 326120 144871 326122 144880
rect 326068 144842 326120 144848
rect 326080 137714 326108 144842
rect 325988 137686 326108 137714
rect 325988 128450 326016 137686
rect 325976 128444 326028 128450
rect 325976 128386 326028 128392
rect 325884 128308 325936 128314
rect 325884 128250 325936 128256
rect 325896 125594 325924 128250
rect 325884 125588 325936 125594
rect 325884 125530 325936 125536
rect 326068 125588 326120 125594
rect 326068 125530 326120 125536
rect 326080 118454 326108 125530
rect 326068 118448 326120 118454
rect 326068 118390 326120 118396
rect 326068 118312 326120 118318
rect 326068 118254 326120 118260
rect 326080 115818 326108 118254
rect 325988 115790 326108 115818
rect 325988 95266 326016 115790
rect 325884 95260 325936 95266
rect 325884 95202 325936 95208
rect 325976 95260 326028 95266
rect 325976 95202 326028 95208
rect 325896 85610 325924 95202
rect 325884 85604 325936 85610
rect 325884 85546 325936 85552
rect 325976 85604 326028 85610
rect 325976 85546 326028 85552
rect 325988 67658 326016 85546
rect 325884 67652 325936 67658
rect 325884 67594 325936 67600
rect 325976 67652 326028 67658
rect 325976 67594 326028 67600
rect 325896 66230 325924 67594
rect 325884 66224 325936 66230
rect 325884 66166 325936 66172
rect 326068 48204 326120 48210
rect 326068 48146 326120 48152
rect 326080 46900 326108 48146
rect 325988 46872 326108 46900
rect 325988 37330 326016 46872
rect 325976 37324 326028 37330
rect 325976 37266 326028 37272
rect 326068 37324 326120 37330
rect 326068 37266 326120 37272
rect 326080 29034 326108 37266
rect 325976 29028 326028 29034
rect 325976 28970 326028 28976
rect 326068 29028 326120 29034
rect 326068 28970 326120 28976
rect 325988 19310 326016 28970
rect 325976 19304 326028 19310
rect 325976 19246 326028 19252
rect 325976 19168 326028 19174
rect 325976 19110 326028 19116
rect 325988 8974 326016 19110
rect 325976 8968 326028 8974
rect 325976 8910 326028 8916
rect 325792 7676 325844 7682
rect 325792 7618 325844 7624
rect 327092 5098 327120 340054
rect 327644 336734 327672 340054
rect 327724 336864 327776 336870
rect 327724 336806 327776 336812
rect 327632 336728 327684 336734
rect 327632 336670 327684 336676
rect 327264 327140 327316 327146
rect 327264 327082 327316 327088
rect 327276 309126 327304 327082
rect 327172 309120 327224 309126
rect 327172 309062 327224 309068
rect 327264 309120 327316 309126
rect 327264 309062 327316 309068
rect 327184 301730 327212 309062
rect 327184 301702 327304 301730
rect 327276 298110 327304 301702
rect 327264 298104 327316 298110
rect 327264 298046 327316 298052
rect 327172 288448 327224 288454
rect 327170 288416 327172 288425
rect 327224 288416 327226 288425
rect 327170 288351 327226 288360
rect 327538 288416 327594 288425
rect 327538 288351 327594 288360
rect 327552 278798 327580 288351
rect 327356 278792 327408 278798
rect 327356 278734 327408 278740
rect 327540 278792 327592 278798
rect 327540 278734 327592 278740
rect 327368 275210 327396 278734
rect 327276 275182 327396 275210
rect 327276 270502 327304 275182
rect 327264 270496 327316 270502
rect 327264 270438 327316 270444
rect 327356 270496 327408 270502
rect 327356 270438 327408 270444
rect 327368 249966 327396 270438
rect 327356 249960 327408 249966
rect 327356 249902 327408 249908
rect 327172 249892 327224 249898
rect 327172 249834 327224 249840
rect 327184 249762 327212 249834
rect 327172 249756 327224 249762
rect 327172 249698 327224 249704
rect 327172 240236 327224 240242
rect 327172 240178 327224 240184
rect 327184 240106 327212 240178
rect 327172 240100 327224 240106
rect 327172 240042 327224 240048
rect 327172 230580 327224 230586
rect 327172 230522 327224 230528
rect 327184 230489 327212 230522
rect 327170 230480 327226 230489
rect 327170 230415 327226 230424
rect 327538 230480 327594 230489
rect 327538 230415 327594 230424
rect 327552 220862 327580 230415
rect 327356 220856 327408 220862
rect 327356 220798 327408 220804
rect 327540 220856 327592 220862
rect 327540 220798 327592 220804
rect 327368 217274 327396 220798
rect 327276 217246 327396 217274
rect 327276 212537 327304 217246
rect 327262 212528 327318 212537
rect 327262 212463 327318 212472
rect 327354 212392 327410 212401
rect 327354 212327 327410 212336
rect 327368 197962 327396 212327
rect 327276 197934 327396 197962
rect 327276 188442 327304 197934
rect 327184 188414 327304 188442
rect 327184 183569 327212 188414
rect 327170 183560 327226 183569
rect 327170 183495 327226 183504
rect 327354 183560 327410 183569
rect 327354 183495 327410 183504
rect 327368 182170 327396 183495
rect 327356 182164 327408 182170
rect 327356 182106 327408 182112
rect 327540 182164 327592 182170
rect 327540 182106 327592 182112
rect 327552 172553 327580 182106
rect 327262 172544 327318 172553
rect 327262 172479 327318 172488
rect 327538 172544 327594 172553
rect 327538 172479 327594 172488
rect 327276 166410 327304 172479
rect 327184 166382 327304 166410
rect 327184 162858 327212 166382
rect 327172 162852 327224 162858
rect 327172 162794 327224 162800
rect 327448 162852 327500 162858
rect 327448 162794 327500 162800
rect 327460 153241 327488 162794
rect 327262 153232 327318 153241
rect 327262 153167 327318 153176
rect 327446 153232 327502 153241
rect 327446 153167 327502 153176
rect 327276 149818 327304 153167
rect 327276 149790 327396 149818
rect 327368 144945 327396 149790
rect 327170 144936 327226 144945
rect 327354 144936 327410 144945
rect 327170 144871 327172 144880
rect 327224 144871 327226 144880
rect 327264 144900 327316 144906
rect 327172 144842 327224 144848
rect 327354 144871 327410 144880
rect 327264 144842 327316 144848
rect 327276 143546 327304 144842
rect 327264 143540 327316 143546
rect 327264 143482 327316 143488
rect 327264 135244 327316 135250
rect 327264 135186 327316 135192
rect 327276 133906 327304 135186
rect 327276 133878 327396 133906
rect 327368 125633 327396 133878
rect 327170 125624 327226 125633
rect 327170 125559 327172 125568
rect 327224 125559 327226 125568
rect 327354 125624 327410 125633
rect 327354 125559 327410 125568
rect 327172 125530 327224 125536
rect 327264 125520 327316 125526
rect 327264 125462 327316 125468
rect 327276 119354 327304 125462
rect 327184 119326 327304 119354
rect 327184 103494 327212 119326
rect 327172 103488 327224 103494
rect 327172 103430 327224 103436
rect 327172 98728 327224 98734
rect 327172 98670 327224 98676
rect 327184 86970 327212 98670
rect 327172 86964 327224 86970
rect 327172 86906 327224 86912
rect 327264 86964 327316 86970
rect 327264 86906 327316 86912
rect 327276 72298 327304 86906
rect 327184 72270 327304 72298
rect 327184 66230 327212 72270
rect 327172 66224 327224 66230
rect 327172 66166 327224 66172
rect 327264 56636 327316 56642
rect 327264 56578 327316 56584
rect 327276 46918 327304 56578
rect 327264 46912 327316 46918
rect 327264 46854 327316 46860
rect 327264 37324 327316 37330
rect 327264 37266 327316 37272
rect 327276 31822 327304 37266
rect 327264 31816 327316 31822
rect 327264 31758 327316 31764
rect 327264 31612 327316 31618
rect 327264 31554 327316 31560
rect 327276 19310 327304 31554
rect 327264 19304 327316 19310
rect 327264 19246 327316 19252
rect 327264 19168 327316 19174
rect 327264 19110 327316 19116
rect 327276 7002 327304 19110
rect 327264 6996 327316 7002
rect 327264 6938 327316 6944
rect 327080 5092 327132 5098
rect 327080 5034 327132 5040
rect 327080 4956 327132 4962
rect 327080 4898 327132 4904
rect 326344 4888 326396 4894
rect 326344 4830 326396 4836
rect 325700 4820 325752 4826
rect 325700 4762 325752 4768
rect 323308 4752 323360 4758
rect 323308 4694 323360 4700
rect 322940 4480 322992 4486
rect 322940 4422 322992 4428
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 322756 3460 322808 3466
rect 322756 3402 322808 3408
rect 322860 480 322888 3538
rect 323320 3058 323348 4694
rect 325148 4480 325200 4486
rect 325148 4422 325200 4428
rect 325160 3670 325188 4422
rect 325148 3664 325200 3670
rect 325148 3606 325200 3612
rect 325240 3664 325292 3670
rect 325240 3606 325292 3612
rect 324044 3460 324096 3466
rect 324044 3402 324096 3408
rect 323308 3052 323360 3058
rect 323308 2994 323360 3000
rect 324056 480 324084 3402
rect 325252 480 325280 3606
rect 326356 2922 326384 4830
rect 326436 3732 326488 3738
rect 326436 3674 326488 3680
rect 326344 2916 326396 2922
rect 326344 2858 326396 2864
rect 326448 480 326476 3674
rect 327092 3602 327120 4898
rect 327080 3596 327132 3602
rect 327080 3538 327132 3544
rect 327736 3126 327764 336806
rect 328552 331356 328604 331362
rect 328552 331298 328604 331304
rect 328274 110800 328330 110809
rect 328458 110800 328514 110809
rect 328330 110758 328458 110786
rect 328274 110735 328330 110744
rect 328458 110735 328514 110744
rect 328564 7750 328592 331298
rect 328656 9042 328684 340054
rect 328748 340054 328946 340082
rect 329024 340054 329406 340082
rect 329958 340054 330064 340082
rect 328644 9036 328696 9042
rect 328644 8978 328696 8984
rect 328552 7744 328604 7750
rect 328552 7686 328604 7692
rect 328748 5030 328776 340054
rect 329024 331362 329052 340054
rect 329840 335640 329892 335646
rect 329840 335582 329892 335588
rect 329012 331356 329064 331362
rect 329012 331298 329064 331304
rect 329852 5098 329880 335582
rect 329932 224256 329984 224262
rect 329932 224198 329984 224204
rect 329944 219473 329972 224198
rect 329930 219464 329986 219473
rect 329930 219399 329986 219408
rect 329932 182164 329984 182170
rect 329932 182106 329984 182112
rect 329944 172553 329972 182106
rect 329930 172544 329986 172553
rect 329930 172479 329986 172488
rect 329932 144356 329984 144362
rect 329932 144298 329984 144304
rect 329944 137970 329972 144298
rect 329932 137964 329984 137970
rect 329932 137906 329984 137912
rect 330036 9110 330064 340054
rect 330128 340054 330418 340082
rect 330128 335646 330156 340054
rect 330116 335640 330168 335646
rect 330116 335582 330168 335588
rect 330496 328506 330524 340190
rect 331324 340054 331430 340082
rect 331508 340054 331890 340082
rect 331968 340054 332350 340082
rect 332796 340054 332902 340082
rect 333072 340054 333362 340082
rect 333440 340054 333822 340082
rect 334176 340054 334374 340082
rect 334544 340054 334834 340082
rect 334912 340054 335294 340082
rect 335464 340054 335846 340082
rect 336016 340054 336306 340082
rect 331324 333282 331352 340054
rect 331324 333254 331444 333282
rect 331220 332172 331272 332178
rect 331220 332114 331272 332120
rect 330208 328500 330260 328506
rect 330208 328442 330260 328448
rect 330484 328500 330536 328506
rect 330484 328442 330536 328448
rect 330220 328386 330248 328442
rect 330128 328358 330248 328386
rect 330128 327078 330156 328358
rect 330116 327072 330168 327078
rect 330116 327014 330168 327020
rect 330208 318844 330260 318850
rect 330208 318786 330260 318792
rect 330220 316033 330248 318786
rect 330206 316024 330262 316033
rect 330206 315959 330262 315968
rect 330390 316024 330446 316033
rect 330390 315959 330446 315968
rect 330404 306406 330432 315959
rect 330208 306400 330260 306406
rect 330208 306342 330260 306348
rect 330392 306400 330444 306406
rect 330392 306342 330444 306348
rect 330220 302326 330248 306342
rect 330208 302320 330260 302326
rect 330208 302262 330260 302268
rect 330116 302184 330168 302190
rect 330116 302126 330168 302132
rect 330128 298058 330156 302126
rect 330206 298072 330262 298081
rect 330128 298030 330206 298058
rect 330206 298007 330262 298016
rect 330390 298072 330446 298081
rect 330390 298007 330446 298016
rect 330404 296698 330432 298007
rect 330312 296670 330432 296698
rect 330312 288454 330340 296670
rect 330300 288448 330352 288454
rect 330300 288390 330352 288396
rect 330300 287088 330352 287094
rect 330300 287030 330352 287036
rect 330312 277438 330340 287030
rect 330116 277432 330168 277438
rect 330116 277374 330168 277380
rect 330300 277432 330352 277438
rect 330300 277374 330352 277380
rect 330128 277302 330156 277374
rect 330116 277296 330168 277302
rect 330116 277238 330168 277244
rect 330116 263220 330168 263226
rect 330116 263162 330168 263168
rect 330128 259418 330156 263162
rect 330116 259412 330168 259418
rect 330116 259354 330168 259360
rect 330208 259412 330260 259418
rect 330208 259354 330260 259360
rect 330220 258058 330248 259354
rect 330208 258052 330260 258058
rect 330208 257994 330260 258000
rect 330392 258052 330444 258058
rect 330392 257994 330444 258000
rect 330404 248441 330432 257994
rect 330206 248432 330262 248441
rect 330206 248367 330262 248376
rect 330390 248432 330446 248441
rect 330390 248367 330446 248376
rect 330220 245018 330248 248367
rect 330128 244990 330248 245018
rect 330128 240106 330156 244990
rect 330116 240100 330168 240106
rect 330116 240042 330168 240048
rect 330208 240100 330260 240106
rect 330208 240042 330260 240048
rect 330220 238746 330248 240042
rect 330208 238740 330260 238746
rect 330208 238682 330260 238688
rect 330392 238672 330444 238678
rect 330392 238614 330444 238620
rect 330404 229129 330432 238614
rect 330206 229120 330262 229129
rect 330206 229055 330262 229064
rect 330390 229120 330446 229129
rect 330390 229055 330446 229064
rect 330220 224262 330248 229055
rect 330208 224256 330260 224262
rect 330208 224198 330260 224204
rect 330114 219464 330170 219473
rect 330114 219399 330116 219408
rect 330168 219399 330170 219408
rect 330116 219370 330168 219376
rect 330116 209840 330168 209846
rect 330168 209788 330248 209794
rect 330116 209782 330248 209788
rect 330128 209778 330248 209782
rect 330128 209772 330260 209778
rect 330128 209766 330208 209772
rect 330208 209714 330260 209720
rect 330220 209683 330248 209714
rect 330116 202836 330168 202842
rect 330116 202778 330168 202784
rect 330128 186386 330156 202778
rect 330116 186380 330168 186386
rect 330116 186322 330168 186328
rect 330116 186244 330168 186250
rect 330116 186186 330168 186192
rect 330128 183569 330156 186186
rect 330114 183560 330170 183569
rect 330114 183495 330170 183504
rect 330114 183424 330170 183433
rect 330114 183359 330170 183368
rect 330128 182170 330156 183359
rect 330116 182164 330168 182170
rect 330116 182106 330168 182112
rect 330206 172544 330262 172553
rect 330206 172479 330262 172488
rect 330220 164354 330248 172479
rect 330116 164348 330168 164354
rect 330116 164290 330168 164296
rect 330208 164348 330260 164354
rect 330208 164290 330260 164296
rect 330128 157978 330156 164290
rect 330482 157992 330538 158001
rect 330128 157950 330432 157978
rect 330404 144362 330432 157950
rect 330482 157927 330538 157936
rect 330496 157729 330524 157927
rect 330482 157720 330538 157729
rect 330482 157655 330538 157664
rect 330392 144356 330444 144362
rect 330392 144298 330444 144304
rect 330208 137964 330260 137970
rect 330208 137906 330260 137912
rect 330220 121446 330248 137906
rect 330208 121440 330260 121446
rect 330208 121382 330260 121388
rect 330576 121440 330628 121446
rect 330576 121382 330628 121388
rect 330588 120086 330616 121382
rect 330576 120080 330628 120086
rect 330576 120022 330628 120028
rect 330576 111784 330628 111790
rect 330576 111726 330628 111732
rect 330588 106758 330616 111726
rect 330576 106752 330628 106758
rect 330576 106694 330628 106700
rect 330208 102196 330260 102202
rect 330208 102138 330260 102144
rect 330220 97306 330248 102138
rect 330208 97300 330260 97306
rect 330208 97242 330260 97248
rect 330300 82952 330352 82958
rect 330300 82894 330352 82900
rect 330312 75970 330340 82894
rect 330220 75942 330340 75970
rect 330220 75886 330248 75942
rect 330208 75880 330260 75886
rect 330208 75822 330260 75828
rect 330208 69964 330260 69970
rect 330208 69906 330260 69912
rect 330220 66178 330248 69906
rect 330220 66150 330340 66178
rect 330312 60602 330340 66150
rect 330220 60574 330340 60602
rect 330220 48362 330248 60574
rect 330128 48334 330248 48362
rect 330128 46918 330156 48334
rect 330116 46912 330168 46918
rect 330116 46854 330168 46860
rect 330116 37324 330168 37330
rect 330116 37266 330168 37272
rect 330128 28937 330156 37266
rect 330482 29336 330538 29345
rect 330482 29271 330538 29280
rect 330496 29073 330524 29271
rect 330482 29064 330538 29073
rect 330482 28999 330538 29008
rect 330114 28928 330170 28937
rect 330114 28863 330170 28872
rect 330206 28792 330262 28801
rect 330206 28727 330262 28736
rect 330220 9654 330248 28727
rect 330208 9648 330260 9654
rect 330208 9590 330260 9596
rect 330024 9104 330076 9110
rect 330024 9046 330076 9052
rect 331232 5166 331260 332114
rect 331312 331764 331364 331770
rect 331312 331706 331364 331712
rect 331324 7886 331352 331706
rect 331416 8362 331444 333254
rect 331508 332178 331536 340054
rect 331496 332172 331548 332178
rect 331496 332114 331548 332120
rect 331968 331770 331996 340054
rect 332692 335708 332744 335714
rect 332692 335650 332744 335656
rect 332600 335640 332652 335646
rect 332600 335582 332652 335588
rect 331956 331764 332008 331770
rect 331956 331706 332008 331712
rect 331404 8356 331456 8362
rect 331404 8298 331456 8304
rect 331312 7880 331364 7886
rect 331312 7822 331364 7828
rect 332612 5234 332640 335582
rect 332704 7954 332732 335650
rect 332796 9178 332824 340054
rect 333072 335646 333100 340054
rect 333244 336932 333296 336938
rect 333244 336874 333296 336880
rect 333060 335640 333112 335646
rect 333060 335582 333112 335588
rect 332784 9172 332836 9178
rect 332784 9114 332836 9120
rect 332692 7948 332744 7954
rect 332692 7890 332744 7896
rect 332600 5228 332652 5234
rect 332600 5170 332652 5176
rect 331220 5160 331272 5166
rect 331220 5102 331272 5108
rect 329840 5092 329892 5098
rect 329840 5034 329892 5040
rect 328736 5024 328788 5030
rect 328736 4966 328788 4972
rect 328460 4820 328512 4826
rect 328460 4762 328512 4768
rect 328472 3738 328500 4762
rect 333256 4146 333284 336874
rect 333440 335714 333468 340054
rect 333428 335708 333480 335714
rect 333428 335650 333480 335656
rect 334072 335708 334124 335714
rect 334072 335650 334124 335656
rect 333980 335640 334032 335646
rect 333980 335582 334032 335588
rect 333612 5024 333664 5030
rect 333612 4966 333664 4972
rect 332416 4140 332468 4146
rect 332416 4082 332468 4088
rect 333244 4140 333296 4146
rect 333244 4082 333296 4088
rect 328460 3732 328512 3738
rect 328460 3674 328512 3680
rect 331220 3732 331272 3738
rect 331220 3674 331272 3680
rect 327724 3120 327776 3126
rect 327724 3062 327776 3068
rect 328828 3120 328880 3126
rect 328828 3062 328880 3068
rect 327632 3052 327684 3058
rect 327632 2994 327684 3000
rect 327644 480 327672 2994
rect 328840 480 328868 3062
rect 330024 2848 330076 2854
rect 330024 2790 330076 2796
rect 330036 480 330064 2790
rect 331232 480 331260 3674
rect 332428 480 332456 4082
rect 333624 480 333652 4966
rect 333992 4690 334020 335582
rect 334084 8022 334112 335650
rect 334176 9246 334204 340054
rect 334544 335646 334572 340054
rect 334912 335714 334940 340054
rect 335268 337136 335320 337142
rect 335268 337078 335320 337084
rect 334900 335708 334952 335714
rect 334900 335650 334952 335656
rect 334532 335640 334584 335646
rect 334532 335582 334584 335588
rect 334164 9240 334216 9246
rect 334164 9182 334216 9188
rect 334072 8016 334124 8022
rect 334072 7958 334124 7964
rect 333980 4684 334032 4690
rect 333980 4626 334032 4632
rect 335280 4146 335308 337078
rect 335360 335640 335412 335646
rect 335360 335582 335412 335588
rect 335372 4554 335400 335582
rect 335464 6594 335492 340054
rect 336016 335646 336044 340054
rect 336096 337680 336148 337686
rect 336096 337622 336148 337628
rect 336004 335640 336056 335646
rect 336004 335582 336056 335588
rect 336108 334506 336136 337622
rect 336752 334558 336780 340068
rect 336844 340054 337318 340082
rect 336016 334478 336136 334506
rect 336740 334552 336792 334558
rect 336740 334494 336792 334500
rect 335452 6588 335504 6594
rect 335452 6530 335504 6536
rect 335360 4548 335412 4554
rect 335360 4490 335412 4496
rect 334716 4140 334768 4146
rect 334716 4082 334768 4088
rect 335268 4140 335320 4146
rect 335268 4082 335320 4088
rect 334728 480 334756 4082
rect 335820 3800 335872 3806
rect 336016 3754 336044 334478
rect 336844 331294 336872 340054
rect 337764 338162 337792 340068
rect 338238 340054 338344 340082
rect 337384 338156 337436 338162
rect 337384 338098 337436 338104
rect 337752 338156 337804 338162
rect 337752 338098 337804 338104
rect 337396 336734 337424 338098
rect 337384 336728 337436 336734
rect 337384 336670 337436 336676
rect 338120 335640 338172 335646
rect 338120 335582 338172 335588
rect 336924 334552 336976 334558
rect 336924 334494 336976 334500
rect 336832 331288 336884 331294
rect 336832 331230 336884 331236
rect 336832 331152 336884 331158
rect 336832 331094 336884 331100
rect 336740 254652 336792 254658
rect 336740 254594 336792 254600
rect 336752 249937 336780 254594
rect 336738 249928 336794 249937
rect 336738 249863 336794 249872
rect 336738 183560 336794 183569
rect 336738 183495 336794 183504
rect 336752 173942 336780 183495
rect 336740 173936 336792 173942
rect 336740 173878 336792 173884
rect 336740 33856 336792 33862
rect 336740 33798 336792 33804
rect 336752 19378 336780 33798
rect 336740 19372 336792 19378
rect 336740 19314 336792 19320
rect 336646 17096 336702 17105
rect 336646 17031 336702 17040
rect 336660 16697 336688 17031
rect 336646 16688 336702 16697
rect 336646 16623 336702 16632
rect 336844 6730 336872 331094
rect 336936 202842 336964 334494
rect 337384 328432 337436 328438
rect 337384 328374 337436 328380
rect 337396 321638 337424 328374
rect 337384 321632 337436 321638
rect 337384 321574 337436 321580
rect 337384 318844 337436 318850
rect 337384 318786 337436 318792
rect 337396 311914 337424 318786
rect 337200 311908 337252 311914
rect 337200 311850 337252 311856
rect 337384 311908 337436 311914
rect 337384 311850 337436 311856
rect 337212 307766 337240 311850
rect 337200 307760 337252 307766
rect 337200 307702 337252 307708
rect 337016 298240 337068 298246
rect 337016 298182 337068 298188
rect 337028 298110 337056 298182
rect 337016 298104 337068 298110
rect 337016 298046 337068 298052
rect 337200 292460 337252 292466
rect 337200 292402 337252 292408
rect 337212 288402 337240 292402
rect 337120 288374 337240 288402
rect 337120 282946 337148 288374
rect 337108 282940 337160 282946
rect 337108 282882 337160 282888
rect 337108 278792 337160 278798
rect 337108 278734 337160 278740
rect 337120 273290 337148 278734
rect 337108 273284 337160 273290
rect 337108 273226 337160 273232
rect 337200 273148 337252 273154
rect 337200 273090 337252 273096
rect 337212 269090 337240 273090
rect 337120 269062 337240 269090
rect 337120 263634 337148 269062
rect 337108 263628 337160 263634
rect 337108 263570 337160 263576
rect 337108 259480 337160 259486
rect 337108 259422 337160 259428
rect 337120 254658 337148 259422
rect 337108 254652 337160 254658
rect 337108 254594 337160 254600
rect 337106 249928 337162 249937
rect 337106 249863 337162 249872
rect 337120 249801 337148 249863
rect 337106 249792 337162 249801
rect 337106 249727 337162 249736
rect 337290 249792 337346 249801
rect 337290 249727 337346 249736
rect 337120 240174 337148 240205
rect 337304 240174 337332 249727
rect 337108 240168 337160 240174
rect 337028 240116 337108 240122
rect 337028 240110 337160 240116
rect 337292 240168 337344 240174
rect 337292 240110 337344 240116
rect 337028 240094 337148 240110
rect 337028 230586 337056 240094
rect 337016 230580 337068 230586
rect 337016 230522 337068 230528
rect 337200 230580 337252 230586
rect 337200 230522 337252 230528
rect 337212 230489 337240 230522
rect 337198 230480 337254 230489
rect 337198 230415 337254 230424
rect 337382 230480 337438 230489
rect 337382 230415 337438 230424
rect 337396 220930 337424 230415
rect 337108 220924 337160 220930
rect 337108 220866 337160 220872
rect 337384 220924 337436 220930
rect 337384 220866 337436 220872
rect 337120 220794 337148 220866
rect 337108 220788 337160 220794
rect 337108 220730 337160 220736
rect 337292 220788 337344 220794
rect 337292 220730 337344 220736
rect 337304 215234 337332 220730
rect 337212 215206 337332 215234
rect 337212 205578 337240 215206
rect 337120 205550 337240 205578
rect 337120 202881 337148 205550
rect 337106 202872 337162 202881
rect 336924 202836 336976 202842
rect 337106 202807 337162 202816
rect 337382 202872 337438 202881
rect 337382 202807 337438 202816
rect 336924 202778 336976 202784
rect 337396 193254 337424 202807
rect 336924 193248 336976 193254
rect 336924 193190 336976 193196
rect 337200 193248 337252 193254
rect 337200 193190 337252 193196
rect 337384 193248 337436 193254
rect 337384 193190 337436 193196
rect 336936 183569 336964 193190
rect 337212 186266 337240 193190
rect 337120 186238 337240 186266
rect 336922 183560 336978 183569
rect 337120 183530 337148 186238
rect 336922 183495 336978 183504
rect 337108 183524 337160 183530
rect 337108 183466 337160 183472
rect 337200 178764 337252 178770
rect 337200 178706 337252 178712
rect 336924 173936 336976 173942
rect 336924 173878 336976 173884
rect 336936 86970 336964 173878
rect 337212 168994 337240 178706
rect 337120 168966 337240 168994
rect 337120 157418 337148 168966
rect 337108 157412 337160 157418
rect 337108 157354 337160 157360
rect 337200 157276 337252 157282
rect 337200 157218 337252 157224
rect 337212 153202 337240 157218
rect 337200 153196 337252 153202
rect 337200 153138 337252 153144
rect 337108 143608 337160 143614
rect 337108 143550 337160 143556
rect 337120 138038 337148 143550
rect 337108 138032 337160 138038
rect 337108 137974 337160 137980
rect 337200 137964 337252 137970
rect 337200 137906 337252 137912
rect 337212 133890 337240 137906
rect 337200 133884 337252 133890
rect 337200 133826 337252 133832
rect 337292 124228 337344 124234
rect 337292 124170 337344 124176
rect 337304 118726 337332 124170
rect 337108 118720 337160 118726
rect 337108 118662 337160 118668
rect 337292 118720 337344 118726
rect 337292 118662 337344 118668
rect 337120 109018 337148 118662
rect 337120 108990 337332 109018
rect 337304 104854 337332 108990
rect 337292 104848 337344 104854
rect 337292 104790 337344 104796
rect 337200 95260 337252 95266
rect 337200 95202 337252 95208
rect 336924 86964 336976 86970
rect 336924 86906 336976 86912
rect 336924 86828 336976 86834
rect 336924 86770 336976 86776
rect 336936 66230 336964 86770
rect 336924 66224 336976 66230
rect 337212 66201 337240 95202
rect 336924 66166 336976 66172
rect 337198 66192 337254 66201
rect 337198 66127 337254 66136
rect 337290 56672 337346 56681
rect 336924 56636 336976 56642
rect 337290 56607 337346 56616
rect 336924 56578 336976 56584
rect 336936 46918 336964 56578
rect 337304 56574 337332 56607
rect 337292 56568 337344 56574
rect 337292 56510 337344 56516
rect 337108 46980 337160 46986
rect 337108 46922 337160 46928
rect 336924 46912 336976 46918
rect 336924 46854 336976 46860
rect 337120 46866 337148 46922
rect 337120 46838 337240 46866
rect 337212 41426 337240 46838
rect 337028 41398 337240 41426
rect 337028 37346 337056 41398
rect 336924 37324 336976 37330
rect 337028 37318 337240 37346
rect 336924 37266 336976 37272
rect 336936 33862 336964 37266
rect 337212 37262 337240 37318
rect 337200 37256 337252 37262
rect 337200 37198 337252 37204
rect 336924 33856 336976 33862
rect 336924 33798 336976 33804
rect 337108 27668 337160 27674
rect 337108 27610 337160 27616
rect 336924 19372 336976 19378
rect 336924 19314 336976 19320
rect 336936 9654 336964 19314
rect 337120 11218 337148 27610
rect 337108 11212 337160 11218
rect 337108 11154 337160 11160
rect 336924 9648 336976 9654
rect 336924 9590 336976 9596
rect 336832 6724 336884 6730
rect 336832 6666 336884 6672
rect 337108 5092 337160 5098
rect 337108 5034 337160 5040
rect 335872 3748 336044 3754
rect 335820 3742 336044 3748
rect 335832 3726 336044 3742
rect 336004 3188 336056 3194
rect 336004 3130 336056 3136
rect 336016 2990 336044 3130
rect 336188 3052 336240 3058
rect 336188 2994 336240 3000
rect 336004 2984 336056 2990
rect 336004 2926 336056 2932
rect 336200 2922 336228 2994
rect 335912 2916 335964 2922
rect 335912 2858 335964 2864
rect 336188 2916 336240 2922
rect 336188 2858 336240 2864
rect 335924 480 335952 2858
rect 337120 480 337148 5034
rect 338132 4486 338160 335582
rect 338316 8158 338344 340054
rect 338408 340054 338790 340082
rect 338960 340054 339250 340082
rect 339604 340054 339710 340082
rect 338304 8152 338356 8158
rect 338304 8094 338356 8100
rect 338408 6662 338436 340054
rect 338764 336932 338816 336938
rect 338764 336874 338816 336880
rect 338396 6656 338448 6662
rect 338396 6598 338448 6604
rect 338120 4480 338172 4486
rect 338120 4422 338172 4428
rect 338776 4146 338804 336874
rect 338960 335646 338988 340054
rect 338948 335640 339000 335646
rect 338948 335582 339000 335588
rect 339500 182164 339552 182170
rect 339500 182106 339552 182112
rect 339512 172553 339540 182106
rect 339498 172544 339554 172553
rect 339498 172479 339554 172488
rect 339500 104848 339552 104854
rect 339500 104790 339552 104796
rect 339512 103494 339540 104790
rect 339500 103488 339552 103494
rect 339500 103430 339552 103436
rect 339500 95260 339552 95266
rect 339500 95202 339552 95208
rect 339512 85610 339540 95202
rect 339500 85604 339552 85610
rect 339500 85546 339552 85552
rect 339604 8226 339632 340054
rect 340248 336802 340276 340068
rect 340708 338162 340736 340068
rect 340984 340054 341182 340082
rect 340328 338156 340380 338162
rect 340328 338098 340380 338104
rect 340696 338156 340748 338162
rect 340696 338098 340748 338104
rect 340236 336796 340288 336802
rect 340236 336738 340288 336744
rect 340340 336734 340368 338098
rect 340788 336932 340840 336938
rect 340788 336874 340840 336880
rect 340328 336728 340380 336734
rect 340328 336670 340380 336676
rect 339776 318844 339828 318850
rect 339776 318786 339828 318792
rect 339788 311930 339816 318786
rect 339696 311902 339816 311930
rect 339696 311846 339724 311902
rect 339684 311840 339736 311846
rect 339684 311782 339736 311788
rect 339868 311840 339920 311846
rect 339868 311782 339920 311788
rect 339880 309126 339908 311782
rect 339868 309120 339920 309126
rect 339868 309062 339920 309068
rect 339868 299940 339920 299946
rect 339868 299882 339920 299888
rect 339880 282946 339908 299882
rect 339684 282940 339736 282946
rect 339684 282882 339736 282888
rect 339868 282940 339920 282946
rect 339868 282882 339920 282888
rect 339696 282826 339724 282882
rect 339696 282798 339816 282826
rect 339788 273306 339816 282798
rect 339788 273278 339908 273306
rect 339880 263634 339908 273278
rect 339684 263628 339736 263634
rect 339684 263570 339736 263576
rect 339868 263628 339920 263634
rect 339868 263570 339920 263576
rect 339696 263514 339724 263570
rect 339696 263486 339816 263514
rect 339788 253994 339816 263486
rect 339788 253966 339908 253994
rect 339880 244322 339908 253966
rect 339684 244316 339736 244322
rect 339684 244258 339736 244264
rect 339868 244316 339920 244322
rect 339868 244258 339920 244264
rect 339696 244202 339724 244258
rect 339696 244174 339816 244202
rect 339788 234682 339816 244174
rect 339788 234654 339908 234682
rect 339880 225010 339908 234654
rect 339684 225004 339736 225010
rect 339684 224946 339736 224952
rect 339868 225004 339920 225010
rect 339868 224946 339920 224952
rect 339696 224890 339724 224946
rect 339696 224862 339816 224890
rect 339788 215370 339816 224862
rect 339788 215342 339908 215370
rect 339880 205698 339908 215342
rect 339684 205692 339736 205698
rect 339684 205634 339736 205640
rect 339868 205692 339920 205698
rect 339868 205634 339920 205640
rect 339696 205578 339724 205634
rect 339696 205550 339816 205578
rect 339788 196058 339816 205550
rect 339788 196030 339908 196058
rect 339880 183054 339908 196030
rect 339684 183048 339736 183054
rect 339684 182990 339736 182996
rect 339868 183048 339920 183054
rect 339868 182990 339920 182996
rect 339696 182170 339724 182990
rect 339684 182164 339736 182170
rect 339684 182106 339736 182112
rect 339866 172544 339922 172553
rect 339866 172479 339922 172488
rect 339880 166954 339908 172479
rect 339788 166926 339908 166954
rect 339788 157434 339816 166926
rect 339788 157406 339908 157434
rect 339880 144945 339908 157406
rect 339682 144936 339738 144945
rect 339682 144871 339738 144880
rect 339866 144936 339922 144945
rect 339866 144871 339922 144880
rect 339696 140026 339724 144871
rect 339696 139998 339908 140026
rect 339880 128382 339908 139998
rect 339684 128376 339736 128382
rect 339868 128376 339920 128382
rect 339736 128324 339868 128330
rect 339684 128318 339920 128324
rect 339696 128302 339908 128318
rect 339880 118794 339908 128302
rect 339868 118788 339920 118794
rect 339868 118730 339920 118736
rect 339776 116000 339828 116006
rect 339776 115942 339828 115948
rect 339788 104854 339816 115942
rect 339776 104848 339828 104854
rect 339776 104790 339828 104796
rect 339868 85604 339920 85610
rect 339868 85546 339920 85552
rect 339880 79914 339908 85546
rect 339788 79886 339908 79914
rect 339788 60738 339816 79886
rect 339696 60722 339816 60738
rect 339684 60716 339816 60722
rect 339736 60710 339816 60716
rect 339868 60716 339920 60722
rect 339684 60658 339736 60664
rect 339868 60658 339920 60664
rect 339880 57934 339908 60658
rect 339868 57928 339920 57934
rect 339868 57870 339920 57876
rect 339776 48340 339828 48346
rect 339776 48282 339828 48288
rect 339788 41426 339816 48282
rect 339696 41398 339816 41426
rect 339696 41290 339724 41398
rect 339696 41262 339816 41290
rect 339788 12458 339816 41262
rect 339696 12430 339816 12458
rect 339592 8220 339644 8226
rect 339592 8162 339644 8168
rect 339696 6526 339724 12430
rect 339684 6520 339736 6526
rect 339684 6462 339736 6468
rect 340800 4146 340828 336874
rect 340880 135244 340932 135250
rect 340880 135186 340932 135192
rect 340892 125633 340920 135186
rect 340878 125624 340934 125633
rect 340878 125559 340934 125568
rect 340984 8294 341012 340054
rect 341628 337550 341656 340068
rect 341720 340054 342194 340082
rect 342364 340054 342654 340082
rect 341616 337544 341668 337550
rect 341616 337486 341668 337492
rect 341720 335594 341748 340054
rect 341800 337272 341852 337278
rect 341800 337214 341852 337220
rect 341168 335566 341748 335594
rect 341168 331226 341196 335566
rect 341812 335458 341840 337214
rect 341536 335430 341840 335458
rect 341156 331220 341208 331226
rect 341156 331162 341208 331168
rect 341340 331220 341392 331226
rect 341340 331162 341392 331168
rect 341352 328438 341380 331162
rect 341340 328432 341392 328438
rect 341340 328374 341392 328380
rect 341432 318844 341484 318850
rect 341432 318786 341484 318792
rect 341444 311914 341472 318786
rect 341248 311908 341300 311914
rect 341248 311850 341300 311856
rect 341432 311908 341484 311914
rect 341432 311850 341484 311856
rect 341260 309126 341288 311850
rect 341248 309120 341300 309126
rect 341248 309062 341300 309068
rect 341156 299532 341208 299538
rect 341156 299474 341208 299480
rect 341168 299418 341196 299474
rect 341246 299432 341302 299441
rect 341168 299390 341246 299418
rect 341246 299367 341302 299376
rect 341246 289912 341302 289921
rect 341246 289847 341302 289856
rect 341260 289814 341288 289847
rect 341248 289808 341300 289814
rect 341248 289750 341300 289756
rect 341156 280220 341208 280226
rect 341156 280162 341208 280168
rect 341168 280106 341196 280162
rect 341246 280120 341302 280129
rect 341168 280078 341246 280106
rect 341246 280055 341302 280064
rect 341246 270600 341302 270609
rect 341246 270535 341302 270544
rect 341260 270502 341288 270535
rect 341248 270496 341300 270502
rect 341248 270438 341300 270444
rect 341156 260908 341208 260914
rect 341156 260850 341208 260856
rect 341168 260794 341196 260850
rect 341246 260808 341302 260817
rect 341168 260766 341246 260794
rect 341246 260743 341302 260752
rect 341246 251288 341302 251297
rect 341246 251223 341302 251232
rect 341260 244390 341288 251223
rect 341248 244384 341300 244390
rect 341248 244326 341300 244332
rect 341156 244248 341208 244254
rect 341156 244190 341208 244196
rect 341168 240145 341196 244190
rect 341154 240136 341210 240145
rect 341154 240071 341210 240080
rect 341430 240136 341486 240145
rect 341430 240071 341486 240080
rect 341444 230518 341472 240071
rect 341248 230512 341300 230518
rect 341248 230454 341300 230460
rect 341432 230512 341484 230518
rect 341432 230454 341484 230460
rect 341260 225078 341288 230454
rect 341248 225072 341300 225078
rect 341248 225014 341300 225020
rect 341156 224936 341208 224942
rect 341156 224878 341208 224884
rect 341168 220794 341196 224878
rect 341156 220788 341208 220794
rect 341156 220730 341208 220736
rect 341156 215280 341208 215286
rect 341156 215222 341208 215228
rect 341168 211154 341196 215222
rect 341168 211126 341288 211154
rect 341260 202910 341288 211126
rect 341156 202904 341208 202910
rect 341154 202872 341156 202881
rect 341248 202904 341300 202910
rect 341208 202872 341210 202881
rect 341248 202846 341300 202852
rect 341430 202872 341486 202881
rect 341154 202807 341210 202816
rect 341430 202807 341486 202816
rect 341444 193254 341472 202807
rect 341248 193248 341300 193254
rect 341248 193190 341300 193196
rect 341432 193248 341484 193254
rect 341432 193190 341484 193196
rect 341260 186266 341288 193190
rect 341168 186238 341288 186266
rect 341168 182170 341196 186238
rect 341156 182164 341208 182170
rect 341156 182106 341208 182112
rect 341432 182164 341484 182170
rect 341432 182106 341484 182112
rect 341444 164234 341472 182106
rect 341260 164206 341472 164234
rect 341260 159390 341288 164206
rect 341064 159384 341116 159390
rect 341064 159326 341116 159332
rect 341248 159384 341300 159390
rect 341248 159326 341300 159332
rect 341076 154578 341104 159326
rect 341076 154562 341288 154578
rect 341064 154556 341300 154562
rect 341116 154550 341248 154556
rect 341064 154498 341116 154504
rect 341248 154498 341300 154504
rect 341076 144945 341104 154498
rect 341260 154467 341288 154498
rect 341062 144936 341118 144945
rect 341062 144871 341118 144880
rect 341246 144936 341302 144945
rect 341246 144871 341302 144880
rect 341260 144786 341288 144871
rect 341260 144758 341472 144786
rect 341444 135289 341472 144758
rect 341246 135280 341302 135289
rect 341246 135215 341248 135224
rect 341300 135215 341302 135224
rect 341430 135280 341486 135289
rect 341430 135215 341486 135224
rect 341248 135186 341300 135192
rect 341062 125624 341118 125633
rect 341062 125559 341064 125568
rect 341116 125559 341118 125568
rect 341064 125530 341116 125536
rect 341156 118652 341208 118658
rect 341156 118594 341208 118600
rect 341168 115954 341196 118594
rect 341168 115938 341288 115954
rect 341168 115932 341300 115938
rect 341168 115926 341248 115932
rect 341248 115874 341300 115880
rect 341432 115932 341484 115938
rect 341432 115874 341484 115880
rect 341260 115843 341288 115874
rect 341444 106321 341472 115874
rect 341246 106312 341302 106321
rect 341246 106247 341302 106256
rect 341430 106312 341486 106321
rect 341430 106247 341486 106256
rect 341260 89706 341288 106247
rect 341168 89678 341288 89706
rect 341168 86970 341196 89678
rect 341156 86964 341208 86970
rect 341156 86906 341208 86912
rect 341064 77308 341116 77314
rect 341064 77250 341116 77256
rect 341076 77178 341104 77250
rect 341064 77172 341116 77178
rect 341064 77114 341116 77120
rect 341156 70304 341208 70310
rect 341156 70246 341208 70252
rect 341168 60722 341196 70246
rect 341156 60716 341208 60722
rect 341156 60658 341208 60664
rect 341340 60716 341392 60722
rect 341340 60658 341392 60664
rect 341352 53122 341380 60658
rect 341260 53094 341380 53122
rect 341260 48521 341288 53094
rect 341246 48512 341302 48521
rect 341246 48447 341302 48456
rect 341430 48376 341486 48385
rect 341430 48311 341486 48320
rect 341444 46918 341472 48311
rect 341432 46912 341484 46918
rect 341432 46854 341484 46860
rect 341248 37324 341300 37330
rect 341248 37266 341300 37272
rect 341260 27742 341288 37266
rect 341248 27736 341300 27742
rect 341248 27678 341300 27684
rect 341156 27668 341208 27674
rect 341156 27610 341208 27616
rect 341168 26246 341196 27610
rect 341156 26240 341208 26246
rect 341156 26182 341208 26188
rect 341248 9716 341300 9722
rect 341248 9658 341300 9664
rect 340972 8288 341024 8294
rect 340972 8230 341024 8236
rect 341260 6458 341288 9658
rect 341248 6452 341300 6458
rect 341248 6394 341300 6400
rect 338764 4140 338816 4146
rect 338764 4082 338816 4088
rect 339500 4140 339552 4146
rect 339500 4082 339552 4088
rect 340788 4140 340840 4146
rect 340788 4082 340840 4088
rect 338304 3732 338356 3738
rect 338304 3674 338356 3680
rect 338316 480 338344 3674
rect 339512 480 339540 4082
rect 341536 3806 341564 335430
rect 342364 6186 342392 340054
rect 342720 337544 342772 337550
rect 342718 337512 342720 337521
rect 342772 337512 342774 337521
rect 342718 337447 342774 337456
rect 342904 337204 342956 337210
rect 342904 337146 342956 337152
rect 342352 6180 342404 6186
rect 342352 6122 342404 6128
rect 342916 3874 342944 337146
rect 343100 336802 343128 340068
rect 343088 336796 343140 336802
rect 343088 336738 343140 336744
rect 343652 6390 343680 340068
rect 344112 337482 344140 340068
rect 344572 337686 344600 340068
rect 345138 340054 345244 340082
rect 344560 337680 344612 337686
rect 344560 337622 344612 337628
rect 344284 337544 344336 337550
rect 344284 337486 344336 337492
rect 344100 337476 344152 337482
rect 344100 337418 344152 337424
rect 343640 6384 343692 6390
rect 343640 6326 343692 6332
rect 342904 3868 342956 3874
rect 342904 3810 342956 3816
rect 343088 3868 343140 3874
rect 343088 3810 343140 3816
rect 341524 3800 341576 3806
rect 341524 3742 341576 3748
rect 341892 3800 341944 3806
rect 341892 3742 341944 3748
rect 341524 3392 341576 3398
rect 340984 3340 341524 3346
rect 340984 3334 341576 3340
rect 340984 3318 341564 3334
rect 340696 3188 340748 3194
rect 340696 3130 340748 3136
rect 340708 480 340736 3130
rect 340984 2922 341012 3318
rect 340972 2916 341024 2922
rect 340972 2858 341024 2864
rect 341904 480 341932 3742
rect 343100 480 343128 3810
rect 344296 3330 344324 337486
rect 344376 336864 344428 336870
rect 344376 336806 344428 336812
rect 344284 3324 344336 3330
rect 344284 3266 344336 3272
rect 344284 2916 344336 2922
rect 344284 2858 344336 2864
rect 344296 480 344324 2858
rect 344388 2854 344416 336806
rect 345216 6254 345244 340054
rect 345584 337618 345612 340068
rect 345676 340054 346058 340082
rect 345572 337612 345624 337618
rect 345572 337554 345624 337560
rect 345676 336818 345704 340054
rect 345756 337612 345808 337618
rect 345756 337554 345808 337560
rect 345768 337521 345796 337554
rect 345754 337512 345810 337521
rect 345754 337447 345810 337456
rect 345940 336932 345992 336938
rect 345584 336802 345704 336818
rect 345572 336796 345704 336802
rect 345624 336790 345704 336796
rect 345860 336892 345940 336920
rect 345572 336738 345624 336744
rect 345860 331242 345888 336892
rect 345940 336874 345992 336880
rect 345676 331214 345888 331242
rect 345204 6248 345256 6254
rect 345204 6190 345256 6196
rect 345676 4146 345704 331214
rect 346306 87136 346362 87145
rect 346306 87071 346362 87080
rect 346320 87009 346348 87071
rect 346306 87000 346362 87009
rect 346306 86935 346362 86944
rect 346596 5302 346624 340068
rect 347056 337890 347084 340068
rect 347044 337884 347096 337890
rect 347044 337826 347096 337832
rect 347516 337482 347544 340068
rect 347976 340054 348082 340082
rect 347504 337476 347556 337482
rect 347504 337418 347556 337424
rect 347780 110560 347832 110566
rect 347778 110528 347780 110537
rect 347832 110528 347834 110537
rect 347778 110463 347834 110472
rect 347780 87032 347832 87038
rect 347778 87000 347780 87009
rect 347832 87000 347834 87009
rect 347778 86935 347834 86944
rect 347780 29096 347832 29102
rect 347778 29064 347780 29073
rect 347832 29064 347834 29073
rect 347778 28999 347834 29008
rect 347778 16960 347834 16969
rect 347778 16895 347780 16904
rect 347832 16895 347834 16904
rect 347780 16866 347832 16872
rect 347976 5370 348004 340054
rect 348528 338706 348556 340068
rect 348516 338700 348568 338706
rect 348516 338642 348568 338648
rect 348424 337884 348476 337890
rect 348424 337826 348476 337832
rect 347964 5364 348016 5370
rect 347964 5306 348016 5312
rect 346584 5296 346636 5302
rect 346584 5238 346636 5244
rect 345664 4140 345716 4146
rect 345664 4082 345716 4088
rect 347872 4140 347924 4146
rect 347872 4082 347924 4088
rect 345756 3256 345808 3262
rect 345492 3204 345756 3210
rect 345492 3198 345808 3204
rect 345492 3182 345796 3198
rect 346676 3188 346728 3194
rect 344376 2848 344428 2854
rect 344376 2790 344428 2796
rect 345492 480 345520 3182
rect 346676 3130 346728 3136
rect 346688 480 346716 3130
rect 347884 480 347912 4082
rect 348436 3330 348464 337826
rect 348988 337278 349016 340068
rect 349356 340054 349554 340082
rect 349068 337476 349120 337482
rect 349068 337418 349120 337424
rect 348976 337272 349028 337278
rect 348976 337214 349028 337220
rect 349080 4146 349108 337418
rect 349356 5438 349384 340054
rect 350000 337686 350028 340068
rect 350184 340054 350474 340082
rect 350644 340054 351026 340082
rect 349988 337680 350040 337686
rect 349988 337622 350040 337628
rect 350184 337618 350212 340054
rect 350172 337612 350224 337618
rect 350172 337554 350224 337560
rect 350644 6322 350672 340054
rect 351184 337612 351236 337618
rect 351184 337554 351236 337560
rect 350632 6316 350684 6322
rect 350632 6258 350684 6264
rect 349344 5432 349396 5438
rect 349344 5374 349396 5380
rect 351196 4146 351224 337554
rect 351472 336802 351500 340068
rect 351932 337822 351960 340068
rect 352116 340054 352498 340082
rect 351920 337816 351972 337822
rect 351920 337758 351972 337764
rect 351828 337544 351880 337550
rect 351828 337486 351880 337492
rect 351460 336796 351512 336802
rect 351460 336738 351512 336744
rect 351840 4146 351868 337486
rect 352116 5506 352144 340054
rect 352944 337958 352972 340068
rect 352932 337952 352984 337958
rect 352932 337894 352984 337900
rect 353404 337006 353432 340068
rect 353496 340054 353970 340082
rect 353392 337000 353444 337006
rect 353392 336942 353444 336948
rect 352564 336796 352616 336802
rect 352564 336738 352616 336744
rect 352104 5500 352156 5506
rect 352104 5442 352156 5448
rect 349068 4140 349120 4146
rect 349068 4082 349120 4088
rect 351184 4140 351236 4146
rect 351184 4082 351236 4088
rect 351368 4140 351420 4146
rect 351368 4082 351420 4088
rect 351828 4140 351880 4146
rect 351828 4082 351880 4088
rect 348424 3324 348476 3330
rect 348424 3266 348476 3272
rect 349068 3324 349120 3330
rect 349068 3266 349120 3272
rect 349080 480 349108 3266
rect 350264 3256 350316 3262
rect 350264 3198 350316 3204
rect 350276 480 350304 3198
rect 351380 480 351408 4082
rect 352576 3074 352604 336738
rect 352656 16924 352708 16930
rect 352656 16866 352708 16872
rect 352668 16697 352696 16866
rect 352654 16688 352710 16697
rect 352654 16623 352710 16632
rect 353496 4418 353524 340054
rect 354416 338094 354444 340068
rect 354404 338088 354456 338094
rect 354404 338030 354456 338036
rect 354876 337686 354904 340068
rect 354968 340054 355442 340082
rect 354864 337680 354916 337686
rect 354864 337622 354916 337628
rect 353484 4412 353536 4418
rect 353484 4354 353536 4360
rect 354968 4350 354996 340054
rect 355888 338026 355916 340068
rect 356256 340054 356362 340082
rect 356624 340054 356914 340082
rect 355876 338020 355928 338026
rect 355876 337962 355928 337968
rect 355324 337952 355376 337958
rect 355324 337894 355376 337900
rect 354956 4344 355008 4350
rect 354956 4286 355008 4292
rect 354956 4140 355008 4146
rect 354956 4082 355008 4088
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 352484 3046 352604 3074
rect 352484 2990 352512 3046
rect 352472 2984 352524 2990
rect 352472 2926 352524 2932
rect 352564 2984 352616 2990
rect 352564 2926 352616 2932
rect 352576 480 352604 2926
rect 353772 480 353800 3334
rect 354968 480 354996 4082
rect 355336 3262 355364 337894
rect 355968 337204 356020 337210
rect 355968 337146 356020 337152
rect 355980 4146 356008 337146
rect 356152 332852 356204 332858
rect 356152 332794 356204 332800
rect 356164 4282 356192 332794
rect 356152 4276 356204 4282
rect 356152 4218 356204 4224
rect 355968 4140 356020 4146
rect 355968 4082 356020 4088
rect 356256 3369 356284 340054
rect 356624 332858 356652 340054
rect 356704 337748 356756 337754
rect 356704 337690 356756 337696
rect 356612 332852 356664 332858
rect 356612 332794 356664 332800
rect 356242 3360 356298 3369
rect 356242 3295 356298 3304
rect 355324 3256 355376 3262
rect 355324 3198 355376 3204
rect 356716 2922 356744 337690
rect 357360 336870 357388 340068
rect 357348 336864 357400 336870
rect 357348 336806 357400 336812
rect 357820 336802 357848 340068
rect 358004 340054 358386 340082
rect 357808 336796 357860 336802
rect 357808 336738 357860 336744
rect 358004 335322 358032 340054
rect 358084 338088 358136 338094
rect 358084 338030 358136 338036
rect 357912 335294 358032 335322
rect 357912 326534 357940 335294
rect 357624 326528 357676 326534
rect 357624 326470 357676 326476
rect 357900 326528 357952 326534
rect 357900 326470 357952 326476
rect 357636 325689 357664 326470
rect 357438 325680 357494 325689
rect 357438 325615 357494 325624
rect 357622 325680 357678 325689
rect 357622 325615 357678 325624
rect 357452 316062 357480 325615
rect 357636 316062 357664 316093
rect 357440 316056 357492 316062
rect 357440 315998 357492 316004
rect 357624 316056 357676 316062
rect 357676 316004 357756 316010
rect 357624 315998 357756 316004
rect 357636 315982 357756 315998
rect 357728 302954 357756 315982
rect 357544 302926 357756 302954
rect 357544 299418 357572 302926
rect 357544 299390 357664 299418
rect 357636 288454 357664 299390
rect 357440 288448 357492 288454
rect 357440 288390 357492 288396
rect 357624 288448 357676 288454
rect 357624 288390 357676 288396
rect 357452 287065 357480 288390
rect 357438 287056 357494 287065
rect 357438 286991 357494 287000
rect 357806 287056 357862 287065
rect 357806 286991 357862 287000
rect 357728 277438 357756 277469
rect 357820 277438 357848 286991
rect 357716 277432 357768 277438
rect 357808 277432 357860 277438
rect 357768 277380 357808 277386
rect 357860 277380 357940 277386
rect 357716 277374 357940 277380
rect 357728 277358 357940 277374
rect 357912 272610 357940 277358
rect 357440 272604 357492 272610
rect 357440 272546 357492 272552
rect 357900 272604 357952 272610
rect 357900 272546 357952 272552
rect 357452 263616 357480 272546
rect 357452 263588 357664 263616
rect 357636 263514 357664 263588
rect 357544 263486 357664 263514
rect 357544 253910 357572 263486
rect 357532 253904 357584 253910
rect 357532 253846 357584 253852
rect 357716 253904 357768 253910
rect 357716 253846 357768 253852
rect 357728 251190 357756 253846
rect 357624 251184 357676 251190
rect 357624 251126 357676 251132
rect 357716 251184 357768 251190
rect 357716 251126 357768 251132
rect 357636 231878 357664 251126
rect 357624 231872 357676 231878
rect 357624 231814 357676 231820
rect 357716 231872 357768 231878
rect 357716 231814 357768 231820
rect 357728 224890 357756 231814
rect 357636 224862 357756 224890
rect 357636 215370 357664 224862
rect 357544 215342 357664 215370
rect 357544 215286 357572 215342
rect 357532 215280 357584 215286
rect 357532 215222 357584 215228
rect 357716 215280 357768 215286
rect 357716 215222 357768 215228
rect 357728 212514 357756 215222
rect 357636 212486 357756 212514
rect 357636 193254 357664 212486
rect 357624 193248 357676 193254
rect 357624 193190 357676 193196
rect 357716 193248 357768 193254
rect 357716 193190 357768 193196
rect 357728 182209 357756 193190
rect 357530 182200 357586 182209
rect 357530 182135 357586 182144
rect 357714 182200 357770 182209
rect 357714 182135 357770 182144
rect 357544 172530 357572 182135
rect 357544 172502 357756 172530
rect 357728 162874 357756 172502
rect 357636 162846 357756 162874
rect 357636 147642 357664 162846
rect 357544 147614 357664 147642
rect 357544 138020 357572 147614
rect 357452 137992 357572 138020
rect 357452 135250 357480 137992
rect 357440 135244 357492 135250
rect 357440 135186 357492 135192
rect 357532 128240 357584 128246
rect 357532 128182 357584 128188
rect 357544 125594 357572 128182
rect 357532 125588 357584 125594
rect 357532 125530 357584 125536
rect 357624 125520 357676 125526
rect 357624 125462 357676 125468
rect 357346 110800 357402 110809
rect 357346 110735 357402 110744
rect 357360 110566 357388 110735
rect 357348 110560 357400 110566
rect 357348 110502 357400 110508
rect 357636 96642 357664 125462
rect 357636 96614 357756 96642
rect 357346 87272 357402 87281
rect 357346 87207 357402 87216
rect 357360 87038 357388 87207
rect 357348 87032 357400 87038
rect 357348 86974 357400 86980
rect 357728 80170 357756 96614
rect 357716 80164 357768 80170
rect 357716 80106 357768 80112
rect 357624 80096 357676 80102
rect 357624 80038 357676 80044
rect 357636 70514 357664 80038
rect 357624 70508 357676 70514
rect 357624 70450 357676 70456
rect 357624 66292 357676 66298
rect 357624 66234 357676 66240
rect 357636 60738 357664 66234
rect 357636 60710 357756 60738
rect 357728 48362 357756 60710
rect 357636 48334 357756 48362
rect 357636 42242 357664 48334
rect 357544 42214 357664 42242
rect 357544 37330 357572 42214
rect 357532 37324 357584 37330
rect 357532 37266 357584 37272
rect 357716 37324 357768 37330
rect 357716 37266 357768 37272
rect 357728 37210 357756 37266
rect 357544 37182 357756 37210
rect 357346 29336 357402 29345
rect 357346 29271 357402 29280
rect 357360 29102 357388 29271
rect 357348 29096 357400 29102
rect 357348 29038 357400 29044
rect 357544 28914 357572 37182
rect 357544 28886 357756 28914
rect 357728 4214 357756 28886
rect 357716 4208 357768 4214
rect 357716 4150 357768 4156
rect 358096 4146 358124 338030
rect 358728 337680 358780 337686
rect 358728 337622 358780 337628
rect 358740 325786 358768 337622
rect 358636 325780 358688 325786
rect 358636 325722 358688 325728
rect 358728 325780 358780 325786
rect 358728 325722 358780 325728
rect 358648 325650 358676 325722
rect 358544 325644 358596 325650
rect 358544 325586 358596 325592
rect 358636 325644 358688 325650
rect 358636 325586 358688 325592
rect 358556 316169 358584 325586
rect 358542 316160 358598 316169
rect 358542 316095 358598 316104
rect 358542 316024 358598 316033
rect 358542 315959 358598 315968
rect 358556 306406 358584 315959
rect 358544 306400 358596 306406
rect 358544 306342 358596 306348
rect 358728 306400 358780 306406
rect 358728 306342 358780 306348
rect 358740 298246 358768 306342
rect 358728 298240 358780 298246
rect 358728 298182 358780 298188
rect 358636 298172 358688 298178
rect 358636 298114 358688 298120
rect 358648 288454 358676 298114
rect 358636 288448 358688 288454
rect 358636 288390 358688 288396
rect 358728 288448 358780 288454
rect 358728 288390 358780 288396
rect 358740 261225 358768 288390
rect 358726 261216 358782 261225
rect 358726 261151 358782 261160
rect 358726 260944 358782 260953
rect 358726 260879 358782 260888
rect 358740 259457 358768 260879
rect 358542 259448 358598 259457
rect 358542 259383 358598 259392
rect 358726 259448 358782 259457
rect 358726 259383 358782 259392
rect 358556 249830 358584 259383
rect 358544 249824 358596 249830
rect 358544 249766 358596 249772
rect 358728 249824 358780 249830
rect 358728 249766 358780 249772
rect 358740 241670 358768 249766
rect 358728 241664 358780 241670
rect 358728 241606 358780 241612
rect 358728 241528 358780 241534
rect 358728 241470 358780 241476
rect 358740 240145 358768 241470
rect 358542 240136 358598 240145
rect 358542 240071 358598 240080
rect 358726 240136 358782 240145
rect 358726 240071 358782 240080
rect 358556 230518 358584 240071
rect 358544 230512 358596 230518
rect 358544 230454 358596 230460
rect 358728 230512 358780 230518
rect 358728 230454 358780 230460
rect 358740 222358 358768 230454
rect 358728 222352 358780 222358
rect 358728 222294 358780 222300
rect 358728 222216 358780 222222
rect 358728 222158 358780 222164
rect 358740 220833 358768 222158
rect 358542 220824 358598 220833
rect 358542 220759 358598 220768
rect 358726 220824 358782 220833
rect 358726 220759 358782 220768
rect 358556 211206 358584 220759
rect 358544 211200 358596 211206
rect 358544 211142 358596 211148
rect 358636 211200 358688 211206
rect 358636 211142 358688 211148
rect 358648 202910 358676 211142
rect 358636 202904 358688 202910
rect 358636 202846 358688 202852
rect 358728 202904 358780 202910
rect 358728 202846 358780 202852
rect 358740 201482 358768 202846
rect 358728 201476 358780 201482
rect 358728 201418 358780 201424
rect 358636 191888 358688 191894
rect 358636 191830 358688 191836
rect 358648 183598 358676 191830
rect 358636 183592 358688 183598
rect 358636 183534 358688 183540
rect 358728 183592 358780 183598
rect 358728 183534 358780 183540
rect 358740 182170 358768 183534
rect 358544 182164 358596 182170
rect 358544 182106 358596 182112
rect 358728 182164 358780 182170
rect 358728 182106 358780 182112
rect 358556 172553 358584 182106
rect 358542 172544 358598 172553
rect 358542 172479 358598 172488
rect 358726 172544 358782 172553
rect 358726 172479 358782 172488
rect 358740 162858 358768 172479
rect 358636 162852 358688 162858
rect 358636 162794 358688 162800
rect 358728 162852 358780 162858
rect 358728 162794 358780 162800
rect 358648 144922 358676 162794
rect 358648 144894 358768 144922
rect 358740 143546 358768 144894
rect 358728 143540 358780 143546
rect 358728 143482 358780 143488
rect 358728 133952 358780 133958
rect 358728 133894 358780 133900
rect 358740 124166 358768 133894
rect 358728 124160 358780 124166
rect 358728 124102 358780 124108
rect 358728 114572 358780 114578
rect 358728 114514 358780 114520
rect 358740 106350 358768 114514
rect 358728 106344 358780 106350
rect 358728 106286 358780 106292
rect 358728 104984 358780 104990
rect 358728 104926 358780 104932
rect 358740 104854 358768 104926
rect 358728 104848 358780 104854
rect 358728 104790 358780 104796
rect 358636 95260 358688 95266
rect 358636 95202 358688 95208
rect 358648 85649 358676 95202
rect 358634 85640 358690 85649
rect 358634 85575 358690 85584
rect 358728 75948 358780 75954
rect 358728 75890 358780 75896
rect 358740 66178 358768 75890
rect 358648 66150 358768 66178
rect 358648 48346 358676 66150
rect 358636 48340 358688 48346
rect 358636 48282 358688 48288
rect 358728 48340 358780 48346
rect 358728 48282 358780 48288
rect 358740 46918 358768 48282
rect 358728 46912 358780 46918
rect 358728 46854 358780 46860
rect 358636 37324 358688 37330
rect 358636 37266 358688 37272
rect 358648 29034 358676 37266
rect 358636 29028 358688 29034
rect 358636 28970 358688 28976
rect 358728 29028 358780 29034
rect 358728 28970 358780 28976
rect 358740 27606 358768 28970
rect 358728 27600 358780 27606
rect 358728 27542 358780 27548
rect 358544 9716 358596 9722
rect 358544 9658 358596 9664
rect 358084 4140 358136 4146
rect 358084 4082 358136 4088
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 356704 2916 356756 2922
rect 356704 2858 356756 2864
rect 356152 2848 356204 2854
rect 356152 2790 356204 2796
rect 356796 2848 356848 2854
rect 357072 2848 357124 2854
rect 356848 2796 357072 2802
rect 356796 2790 357124 2796
rect 356164 480 356192 2790
rect 356808 2774 357112 2790
rect 357360 480 357388 3198
rect 358556 480 358584 9658
rect 358832 4010 358860 340068
rect 358924 340054 359306 340082
rect 359476 340054 359766 340082
rect 358820 4004 358872 4010
rect 358820 3946 358872 3952
rect 358924 3670 358952 340054
rect 359476 337362 359504 340054
rect 359200 337334 359504 337362
rect 359200 318918 359228 337334
rect 359464 337272 359516 337278
rect 359464 337214 359516 337220
rect 359188 318912 359240 318918
rect 359188 318854 359240 318860
rect 359096 318844 359148 318850
rect 359096 318786 359148 318792
rect 359108 311896 359136 318786
rect 359108 311868 359228 311896
rect 359200 299690 359228 311868
rect 359108 299662 359228 299690
rect 359108 298110 359136 299662
rect 359096 298104 359148 298110
rect 359096 298046 359148 298052
rect 359188 298104 359240 298110
rect 359188 298046 359240 298052
rect 359200 282826 359228 298046
rect 359108 282798 359228 282826
rect 359108 273306 359136 282798
rect 359016 273278 359136 273306
rect 359016 273222 359044 273278
rect 359004 273216 359056 273222
rect 359004 273158 359056 273164
rect 359188 273216 359240 273222
rect 359188 273158 359240 273164
rect 359200 260914 359228 273158
rect 359096 260908 359148 260914
rect 359096 260850 359148 260856
rect 359188 260908 359240 260914
rect 359188 260850 359240 260856
rect 359108 253994 359136 260850
rect 359016 253966 359136 253994
rect 359016 253910 359044 253966
rect 359004 253904 359056 253910
rect 359004 253846 359056 253852
rect 359188 253904 359240 253910
rect 359188 253846 359240 253852
rect 359200 241534 359228 253846
rect 359096 241528 359148 241534
rect 359096 241470 359148 241476
rect 359188 241528 359240 241534
rect 359188 241470 359240 241476
rect 359108 231878 359136 241470
rect 359096 231872 359148 231878
rect 359096 231814 359148 231820
rect 359188 231872 359240 231878
rect 359188 231814 359240 231820
rect 359200 224890 359228 231814
rect 359108 224862 359228 224890
rect 359108 215370 359136 224862
rect 359016 215342 359136 215370
rect 359016 215286 359044 215342
rect 359004 215280 359056 215286
rect 359004 215222 359056 215228
rect 359188 215280 359240 215286
rect 359188 215222 359240 215228
rect 359200 202910 359228 215222
rect 359096 202904 359148 202910
rect 359096 202846 359148 202852
rect 359188 202904 359240 202910
rect 359188 202846 359240 202852
rect 359108 193254 359136 202846
rect 359096 193248 359148 193254
rect 359096 193190 359148 193196
rect 359188 193248 359240 193254
rect 359188 193190 359240 193196
rect 359200 182209 359228 193190
rect 359002 182200 359058 182209
rect 359002 182135 359058 182144
rect 359186 182200 359242 182209
rect 359186 182135 359242 182144
rect 359016 179382 359044 182135
rect 359004 179376 359056 179382
rect 359004 179318 359056 179324
rect 359096 169788 359148 169794
rect 359096 169730 359148 169736
rect 359108 162874 359136 169730
rect 359016 162858 359136 162874
rect 359004 162852 359148 162858
rect 359056 162846 359096 162852
rect 359004 162794 359056 162800
rect 359096 162794 359148 162800
rect 359108 161430 359136 162794
rect 359096 161424 359148 161430
rect 359096 161366 359148 161372
rect 359188 151836 359240 151842
rect 359188 151778 359240 151784
rect 359200 144906 359228 151778
rect 359188 144900 359240 144906
rect 359188 144842 359240 144848
rect 359280 144900 359332 144906
rect 359280 144842 359332 144848
rect 359292 139890 359320 144842
rect 359200 139862 359320 139890
rect 359200 128330 359228 139862
rect 359108 128302 359228 128330
rect 359108 118708 359136 128302
rect 359108 118680 359228 118708
rect 359200 118538 359228 118680
rect 359108 118510 359228 118538
rect 359108 96642 359136 118510
rect 359108 96614 359228 96642
rect 359002 85368 359058 85377
rect 359002 85303 359058 85312
rect 359016 75954 359044 85303
rect 359004 75948 359056 75954
rect 359004 75890 359056 75896
rect 359200 74594 359228 96614
rect 359096 74588 359148 74594
rect 359096 74530 359148 74536
rect 359188 74588 359240 74594
rect 359188 74530 359240 74536
rect 359108 64870 359136 74530
rect 359096 64864 359148 64870
rect 359096 64806 359148 64812
rect 359096 56568 359148 56574
rect 359096 56510 359148 56516
rect 359108 46918 359136 56510
rect 359096 46912 359148 46918
rect 359096 46854 359148 46860
rect 359188 37324 359240 37330
rect 359188 37266 359240 37272
rect 359200 29102 359228 37266
rect 359188 29096 359240 29102
rect 359188 29038 359240 29044
rect 359188 28960 359240 28966
rect 359188 28902 359240 28908
rect 359200 4758 359228 28902
rect 359188 4752 359240 4758
rect 359188 4694 359240 4700
rect 358912 3664 358964 3670
rect 358912 3606 358964 3612
rect 359476 3126 359504 337214
rect 360304 336938 360332 340068
rect 360764 337754 360792 340068
rect 360948 340054 361238 340082
rect 360752 337748 360804 337754
rect 360752 337690 360804 337696
rect 360292 336932 360344 336938
rect 360292 336874 360344 336880
rect 360948 331242 360976 340054
rect 361776 337346 361804 340068
rect 361868 340054 362250 340082
rect 362328 340054 362710 340082
rect 363156 340054 363262 340082
rect 361764 337340 361816 337346
rect 361764 337282 361816 337288
rect 361672 335640 361724 335646
rect 361672 335582 361724 335588
rect 360304 331226 360976 331242
rect 360292 331220 360976 331226
rect 360344 331214 360476 331220
rect 360292 331162 360344 331168
rect 360528 331214 360976 331220
rect 360476 331162 360528 331168
rect 360488 323626 360516 331162
rect 360488 323598 360608 323626
rect 360580 311914 360608 323598
rect 360200 311908 360252 311914
rect 360200 311850 360252 311856
rect 360568 311908 360620 311914
rect 360568 311850 360620 311856
rect 360212 309126 360240 311850
rect 360200 309120 360252 309126
rect 360200 309062 360252 309068
rect 360292 309120 360344 309126
rect 360292 309062 360344 309068
rect 360304 302138 360332 309062
rect 360304 302110 360516 302138
rect 360488 293298 360516 302110
rect 360396 293270 360516 293298
rect 360396 273306 360424 293270
rect 360396 273278 360516 273306
rect 360488 263634 360516 273278
rect 360292 263628 360344 263634
rect 360292 263570 360344 263576
rect 360476 263628 360528 263634
rect 360476 263570 360528 263576
rect 360304 263514 360332 263570
rect 360304 263486 360424 263514
rect 360396 253994 360424 263486
rect 360396 253966 360516 253994
rect 360488 244322 360516 253966
rect 360292 244316 360344 244322
rect 360292 244258 360344 244264
rect 360476 244316 360528 244322
rect 360476 244258 360528 244264
rect 360304 244202 360332 244258
rect 360304 244174 360424 244202
rect 360396 234682 360424 244174
rect 360396 234654 360516 234682
rect 360488 225010 360516 234654
rect 360292 225004 360344 225010
rect 360292 224946 360344 224952
rect 360476 225004 360528 225010
rect 360476 224946 360528 224952
rect 360304 224890 360332 224946
rect 360304 224862 360424 224890
rect 360396 215370 360424 224862
rect 360396 215342 360516 215370
rect 360488 205698 360516 215342
rect 360292 205692 360344 205698
rect 360292 205634 360344 205640
rect 360476 205692 360528 205698
rect 360476 205634 360528 205640
rect 360304 205578 360332 205634
rect 360304 205550 360424 205578
rect 360396 196058 360424 205550
rect 360396 196030 360516 196058
rect 360488 182481 360516 196030
rect 360474 182472 360530 182481
rect 360474 182407 360530 182416
rect 360290 182200 360346 182209
rect 360290 182135 360346 182144
rect 360304 171086 360332 182135
rect 360292 171080 360344 171086
rect 360292 171022 360344 171028
rect 360476 161492 360528 161498
rect 360476 161434 360528 161440
rect 360488 128382 360516 161434
rect 360292 128376 360344 128382
rect 360476 128376 360528 128382
rect 360344 128324 360424 128330
rect 360292 128318 360424 128324
rect 360476 128318 360528 128324
rect 360304 128302 360424 128318
rect 360396 120714 360424 128302
rect 360396 120686 360608 120714
rect 360580 118674 360608 120686
rect 360488 118646 360608 118674
rect 360488 95305 360516 118646
rect 360474 95296 360530 95305
rect 360474 95231 360530 95240
rect 360382 95160 360438 95169
rect 360382 95095 360438 95104
rect 360396 85542 360424 95095
rect 360384 85536 360436 85542
rect 360384 85478 360436 85484
rect 360200 75948 360252 75954
rect 360200 75890 360252 75896
rect 360212 70258 360240 75890
rect 360212 70230 360332 70258
rect 360304 60722 360332 70230
rect 360292 60716 360344 60722
rect 360292 60658 360344 60664
rect 360476 60716 360528 60722
rect 360476 60658 360528 60664
rect 360488 52850 360516 60658
rect 360396 52822 360516 52850
rect 360396 41426 360424 52822
rect 360304 41410 360424 41426
rect 360292 41404 360424 41410
rect 360344 41398 360424 41404
rect 360476 41404 360528 41410
rect 360292 41346 360344 41352
rect 360476 41346 360528 41352
rect 360488 12458 360516 41346
rect 360304 12430 360516 12458
rect 360304 4894 360332 12430
rect 361684 4962 361712 335582
rect 361672 4956 361724 4962
rect 361672 4898 361724 4904
rect 360292 4888 360344 4894
rect 360292 4830 360344 4836
rect 359740 4004 359792 4010
rect 359740 3946 359792 3952
rect 359464 3120 359516 3126
rect 359464 3062 359516 3068
rect 359752 480 359780 3946
rect 360936 3664 360988 3670
rect 360936 3606 360988 3612
rect 360948 480 360976 3606
rect 361868 3602 361896 340054
rect 362224 336864 362276 336870
rect 362224 336806 362276 336812
rect 362236 335458 362264 336806
rect 362328 335646 362356 340054
rect 362868 337816 362920 337822
rect 362868 337758 362920 337764
rect 362316 335640 362368 335646
rect 362316 335582 362368 335588
rect 362236 335430 362356 335458
rect 362328 318918 362356 335430
rect 362316 318912 362368 318918
rect 362316 318854 362368 318860
rect 362224 318844 362276 318850
rect 362224 318786 362276 318792
rect 362236 312066 362264 318786
rect 362052 312038 362264 312066
rect 362052 306377 362080 312038
rect 362038 306368 362094 306377
rect 362038 306303 362094 306312
rect 362406 306368 362462 306377
rect 362406 306303 362462 306312
rect 362420 296750 362448 306303
rect 362224 296744 362276 296750
rect 362224 296686 362276 296692
rect 362408 296744 362460 296750
rect 362408 296686 362460 296692
rect 362236 277370 362264 296686
rect 362224 277364 362276 277370
rect 362224 277306 362276 277312
rect 362224 263492 362276 263498
rect 362224 263434 362276 263440
rect 362236 259434 362264 263434
rect 362236 259406 362356 259434
rect 362328 253978 362356 259406
rect 362316 253972 362368 253978
rect 362316 253914 362368 253920
rect 362224 253904 362276 253910
rect 362224 253846 362276 253852
rect 362236 241466 362264 253846
rect 362224 241460 362276 241466
rect 362224 241402 362276 241408
rect 362408 230512 362460 230518
rect 362408 230454 362460 230460
rect 362420 222222 362448 230454
rect 362224 222216 362276 222222
rect 362224 222158 362276 222164
rect 362408 222216 362460 222222
rect 362408 222158 362460 222164
rect 362236 220810 362264 222158
rect 362236 220782 362356 220810
rect 362328 215354 362356 220782
rect 362316 215348 362368 215354
rect 362316 215290 362368 215296
rect 362132 211200 362184 211206
rect 362132 211142 362184 211148
rect 362144 202910 362172 211142
rect 362132 202904 362184 202910
rect 362132 202846 362184 202852
rect 362224 202904 362276 202910
rect 362224 202846 362276 202852
rect 362236 198082 362264 202846
rect 362224 198076 362276 198082
rect 362224 198018 362276 198024
rect 362316 193248 362368 193254
rect 362316 193190 362368 193196
rect 362328 182238 362356 193190
rect 362224 182232 362276 182238
rect 362224 182174 362276 182180
rect 362316 182232 362368 182238
rect 362316 182174 362368 182180
rect 362236 172530 362264 182174
rect 362236 172502 362356 172530
rect 362328 171086 362356 172502
rect 362316 171080 362368 171086
rect 362316 171022 362368 171028
rect 362224 161492 362276 161498
rect 362224 161434 362276 161440
rect 362236 161378 362264 161434
rect 362236 161350 362356 161378
rect 362328 156618 362356 161350
rect 362144 156590 362356 156618
rect 362144 144906 362172 156590
rect 362132 144900 362184 144906
rect 362132 144842 362184 144848
rect 362316 144900 362368 144906
rect 362316 144842 362368 144848
rect 362328 143546 362356 144842
rect 362316 143540 362368 143546
rect 362316 143482 362368 143488
rect 362500 143540 362552 143546
rect 362500 143482 362552 143488
rect 362512 133929 362540 143482
rect 362314 133920 362370 133929
rect 362314 133855 362370 133864
rect 362498 133920 362554 133929
rect 362498 133855 362554 133864
rect 362328 120714 362356 133855
rect 362236 120686 362356 120714
rect 362236 109138 362264 120686
rect 362224 109132 362276 109138
rect 362224 109074 362276 109080
rect 362132 108996 362184 109002
rect 362132 108938 362184 108944
rect 362144 100042 362172 108938
rect 362144 100014 362356 100042
rect 362328 95198 362356 100014
rect 362316 95192 362368 95198
rect 362316 95134 362368 95140
rect 362408 85604 362460 85610
rect 362408 85546 362460 85552
rect 362420 75954 362448 85546
rect 362224 75948 362276 75954
rect 362224 75890 362276 75896
rect 362408 75948 362460 75954
rect 362408 75890 362460 75896
rect 362236 74526 362264 75890
rect 362224 74520 362276 74526
rect 362224 74462 362276 74468
rect 362408 74520 362460 74526
rect 362408 74462 362460 74468
rect 362420 64954 362448 74462
rect 362420 64926 362540 64954
rect 362512 64870 362540 64926
rect 362500 64864 362552 64870
rect 362500 64806 362552 64812
rect 362224 55276 362276 55282
rect 362224 55218 362276 55224
rect 362236 41478 362264 55218
rect 362224 41472 362276 41478
rect 362224 41414 362276 41420
rect 362224 38616 362276 38622
rect 362224 38558 362276 38564
rect 362236 27554 362264 38558
rect 362236 27526 362356 27554
rect 362328 18086 362356 27526
rect 362316 18080 362368 18086
rect 362316 18022 362368 18028
rect 362224 8356 362276 8362
rect 362224 8298 362276 8304
rect 362132 4140 362184 4146
rect 362132 4082 362184 4088
rect 361856 3596 361908 3602
rect 361856 3538 361908 3544
rect 362144 480 362172 4082
rect 362236 2786 362264 8298
rect 362880 4146 362908 337758
rect 363052 335640 363104 335646
rect 363052 335582 363104 335588
rect 363064 4826 363092 335582
rect 363052 4820 363104 4826
rect 363052 4762 363104 4768
rect 362868 4140 362920 4146
rect 362868 4082 362920 4088
rect 363156 3534 363184 340054
rect 363708 337278 363736 340068
rect 363800 340054 364182 340082
rect 363696 337272 363748 337278
rect 363696 337214 363748 337220
rect 363604 336796 363656 336802
rect 363604 336738 363656 336744
rect 363328 4140 363380 4146
rect 363328 4082 363380 4088
rect 363144 3528 363196 3534
rect 363144 3470 363196 3476
rect 362224 2780 362276 2786
rect 362224 2722 362276 2728
rect 363340 480 363368 4082
rect 363616 3466 363644 336738
rect 363800 335646 363828 340054
rect 364248 338020 364300 338026
rect 364248 337962 364300 337968
rect 363788 335640 363840 335646
rect 363788 335582 363840 335588
rect 364260 4146 364288 337962
rect 364720 336802 364748 340068
rect 365180 336870 365208 340068
rect 365640 337890 365668 340068
rect 365824 340054 366206 340082
rect 365628 337884 365680 337890
rect 365628 337826 365680 337832
rect 365168 336864 365220 336870
rect 365168 336806 365220 336812
rect 364708 336796 364760 336802
rect 364708 336738 364760 336744
rect 364248 4140 364300 4146
rect 364248 4082 364300 4088
rect 365720 4140 365772 4146
rect 365720 4082 365772 4088
rect 363604 3460 363656 3466
rect 363604 3402 363656 3408
rect 365536 3324 365588 3330
rect 365536 3266 365588 3272
rect 365548 3058 365576 3266
rect 364524 3052 364576 3058
rect 364524 2994 364576 3000
rect 365536 3052 365588 3058
rect 365536 2994 365588 3000
rect 364536 480 364564 2994
rect 365732 480 365760 4082
rect 365824 3942 365852 340054
rect 366652 337142 366680 340068
rect 367126 340054 367232 340082
rect 367008 337612 367060 337618
rect 367008 337554 367060 337560
rect 366916 337340 366968 337346
rect 366916 337282 366968 337288
rect 366640 337136 366692 337142
rect 366640 337078 366692 337084
rect 366822 241496 366878 241505
rect 366822 241431 366878 241440
rect 366836 231946 366864 241431
rect 366824 231940 366876 231946
rect 366824 231882 366876 231888
rect 366822 202872 366878 202881
rect 366822 202807 366878 202816
rect 366836 193322 366864 202807
rect 366824 193316 366876 193322
rect 366824 193258 366876 193264
rect 366824 115864 366876 115870
rect 366824 115806 366876 115812
rect 366836 106321 366864 115806
rect 366822 106312 366878 106321
rect 366822 106247 366878 106256
rect 366928 19310 366956 337282
rect 367020 309126 367048 337554
rect 367008 309120 367060 309126
rect 367008 309062 367060 309068
rect 367008 299532 367060 299538
rect 367008 299474 367060 299480
rect 367020 289814 367048 299474
rect 367008 289808 367060 289814
rect 367008 289750 367060 289756
rect 367008 280220 367060 280226
rect 367008 280162 367060 280168
rect 367020 270502 367048 280162
rect 367008 270496 367060 270502
rect 367008 270438 367060 270444
rect 367008 260908 367060 260914
rect 367008 260850 367060 260856
rect 367020 251190 367048 260850
rect 367008 251184 367060 251190
rect 367008 251126 367060 251132
rect 367008 241528 367060 241534
rect 367006 241496 367008 241505
rect 367060 241496 367062 241505
rect 367006 241431 367062 241440
rect 367008 231940 367060 231946
rect 367008 231882 367060 231888
rect 367020 231810 367048 231882
rect 367008 231804 367060 231810
rect 367008 231746 367060 231752
rect 367008 222216 367060 222222
rect 367008 222158 367060 222164
rect 367020 202881 367048 222158
rect 367006 202872 367062 202881
rect 367006 202807 367062 202816
rect 367008 193316 367060 193322
rect 367008 193258 367060 193264
rect 367020 193186 367048 193258
rect 367008 193180 367060 193186
rect 367008 193122 367060 193128
rect 367008 183592 367060 183598
rect 367008 183534 367060 183540
rect 367020 144906 367048 183534
rect 367008 144900 367060 144906
rect 367008 144842 367060 144848
rect 367008 135312 367060 135318
rect 367008 135254 367060 135260
rect 367020 125594 367048 135254
rect 367008 125588 367060 125594
rect 367008 125530 367060 125536
rect 367008 116000 367060 116006
rect 367008 115942 367060 115948
rect 367020 115870 367048 115942
rect 367008 115864 367060 115870
rect 367008 115806 367060 115812
rect 367006 106312 367062 106321
rect 367006 106247 367062 106256
rect 367020 96937 367048 106247
rect 367006 96928 367062 96937
rect 367006 96863 367062 96872
rect 367006 96656 367062 96665
rect 367006 96591 367008 96600
rect 367060 96591 367062 96600
rect 367008 96562 367060 96568
rect 367008 87032 367060 87038
rect 367008 86974 367060 86980
rect 367020 57934 367048 86974
rect 367100 76220 367152 76226
rect 367100 76162 367152 76168
rect 367112 76129 367140 76162
rect 367098 76120 367154 76129
rect 367098 76055 367154 76064
rect 367008 57928 367060 57934
rect 367008 57870 367060 57876
rect 367008 48340 367060 48346
rect 367008 48282 367060 48288
rect 367020 38622 367048 48282
rect 367008 38616 367060 38622
rect 367008 38558 367060 38564
rect 367098 29200 367154 29209
rect 367098 29135 367154 29144
rect 367008 29096 367060 29102
rect 367112 29073 367140 29135
rect 367008 29038 367060 29044
rect 367098 29064 367154 29073
rect 367020 28966 367048 29038
rect 367098 28999 367154 29008
rect 367008 28960 367060 28966
rect 367008 28902 367060 28908
rect 367008 19372 367060 19378
rect 367008 19314 367060 19320
rect 366916 19304 366968 19310
rect 366916 19246 366968 19252
rect 367020 14414 367048 19314
rect 366824 14408 366876 14414
rect 366824 14350 366876 14356
rect 367008 14408 367060 14414
rect 367008 14350 367060 14356
rect 365812 3936 365864 3942
rect 365812 3878 365864 3884
rect 366836 2802 366864 14350
rect 366916 10124 366968 10130
rect 366916 10066 366968 10072
rect 366928 4146 366956 10066
rect 367204 5030 367232 340054
rect 367664 337074 367692 340068
rect 367940 340054 368138 340082
rect 367652 337068 367704 337074
rect 367652 337010 367704 337016
rect 367940 335646 367968 340054
rect 367284 335640 367336 335646
rect 367284 335582 367336 335588
rect 367928 335640 367980 335646
rect 367928 335582 367980 335588
rect 367192 5024 367244 5030
rect 367192 4966 367244 4972
rect 366916 4140 366968 4146
rect 366916 4082 366968 4088
rect 367296 2922 367324 335582
rect 368204 110696 368256 110702
rect 368204 110638 368256 110644
rect 368216 110537 368244 110638
rect 368202 110528 368258 110537
rect 368202 110463 368258 110472
rect 368584 5098 368612 340068
rect 368676 340054 369150 340082
rect 368572 5092 368624 5098
rect 368572 5034 368624 5040
rect 368676 3738 368704 340054
rect 369124 337136 369176 337142
rect 369124 337078 369176 337084
rect 369136 3874 369164 337078
rect 369596 337006 369624 340068
rect 370056 337958 370084 340068
rect 370148 340054 370622 340082
rect 370044 337952 370096 337958
rect 370044 337894 370096 337900
rect 369768 337408 369820 337414
rect 369768 337350 369820 337356
rect 369584 337000 369636 337006
rect 369584 336942 369636 336948
rect 369780 4146 369808 337350
rect 369216 4140 369268 4146
rect 369216 4082 369268 4088
rect 369768 4140 369820 4146
rect 369768 4082 369820 4088
rect 369124 3868 369176 3874
rect 369124 3810 369176 3816
rect 368664 3732 368716 3738
rect 368664 3674 368716 3680
rect 368020 3460 368072 3466
rect 368020 3402 368072 3408
rect 367284 2916 367336 2922
rect 367284 2858 367336 2864
rect 366836 2774 366956 2802
rect 366928 480 366956 2774
rect 368032 480 368060 3402
rect 369228 480 369256 4082
rect 370148 3806 370176 340054
rect 371068 337142 371096 340068
rect 371528 338094 371556 340068
rect 372080 338162 372108 340068
rect 372068 338156 372120 338162
rect 372068 338098 372120 338104
rect 371516 338088 371568 338094
rect 371516 338030 371568 338036
rect 371148 337952 371200 337958
rect 371148 337894 371200 337900
rect 371056 337136 371108 337142
rect 371056 337078 371108 337084
rect 370504 336796 370556 336802
rect 370504 336738 370556 336744
rect 370412 4140 370464 4146
rect 370412 4082 370464 4088
rect 370136 3800 370188 3806
rect 370136 3742 370188 3748
rect 370424 480 370452 4082
rect 370516 3194 370544 336738
rect 371160 4146 371188 337894
rect 372540 336802 372568 340068
rect 373000 337278 373028 340068
rect 373276 340054 373566 340082
rect 372988 337272 373040 337278
rect 372988 337214 373040 337220
rect 372528 336796 372580 336802
rect 372528 336738 372580 336744
rect 373276 335646 373304 340054
rect 373908 337544 373960 337550
rect 373908 337486 373960 337492
rect 372620 335640 372672 335646
rect 372620 335582 372672 335588
rect 373264 335640 373316 335646
rect 373264 335582 373316 335588
rect 372632 331106 372660 335582
rect 372632 331078 372752 331106
rect 372724 318782 372752 331078
rect 372712 318776 372764 318782
rect 372712 318718 372764 318724
rect 372712 309188 372764 309194
rect 372712 309130 372764 309136
rect 372724 299470 372752 309130
rect 372712 299464 372764 299470
rect 372712 299406 372764 299412
rect 372712 289876 372764 289882
rect 372712 289818 372764 289824
rect 372724 280158 372752 289818
rect 372712 280152 372764 280158
rect 372712 280094 372764 280100
rect 372712 270564 372764 270570
rect 372712 270506 372764 270512
rect 372724 260846 372752 270506
rect 372712 260840 372764 260846
rect 372712 260782 372764 260788
rect 372712 251252 372764 251258
rect 372712 251194 372764 251200
rect 372724 241505 372752 251194
rect 372526 241496 372582 241505
rect 372526 241431 372582 241440
rect 372710 241496 372766 241505
rect 372710 241431 372766 241440
rect 372540 231878 372568 241431
rect 372528 231872 372580 231878
rect 372528 231814 372580 231820
rect 372712 231872 372764 231878
rect 372712 231814 372764 231820
rect 372724 222193 372752 231814
rect 372526 222184 372582 222193
rect 372526 222119 372582 222128
rect 372710 222184 372766 222193
rect 372710 222119 372766 222128
rect 372540 212566 372568 222119
rect 372528 212560 372580 212566
rect 372528 212502 372580 212508
rect 372712 212560 372764 212566
rect 372712 212502 372764 212508
rect 372724 202881 372752 212502
rect 372526 202872 372582 202881
rect 372526 202807 372582 202816
rect 372710 202872 372766 202881
rect 372710 202807 372766 202816
rect 372540 193254 372568 202807
rect 372528 193248 372580 193254
rect 372528 193190 372580 193196
rect 372712 193248 372764 193254
rect 372712 193190 372764 193196
rect 372724 178786 372752 193190
rect 372632 178758 372752 178786
rect 372632 174010 372660 178758
rect 372620 174004 372672 174010
rect 372620 173946 372672 173952
rect 372804 174004 372856 174010
rect 372804 173946 372856 173952
rect 372816 173913 372844 173946
rect 372802 173904 372858 173913
rect 372802 173839 372858 173848
rect 372986 173904 373042 173913
rect 372986 173839 373042 173848
rect 373000 164257 373028 173839
rect 372802 164248 372858 164257
rect 372802 164183 372804 164192
rect 372856 164183 372858 164192
rect 372986 164248 373042 164257
rect 372986 164183 373042 164192
rect 372804 164154 372856 164160
rect 372804 157344 372856 157350
rect 372804 157286 372856 157292
rect 372816 138174 372844 157286
rect 372804 138168 372856 138174
rect 372804 138110 372856 138116
rect 372712 135312 372764 135318
rect 372712 135254 372764 135260
rect 372724 118810 372752 135254
rect 372632 118782 372752 118810
rect 372632 118674 372660 118782
rect 372632 118646 372752 118674
rect 372724 101402 372752 118646
rect 372632 101374 372752 101402
rect 372632 96626 372660 101374
rect 372620 96620 372672 96626
rect 372620 96562 372672 96568
rect 372712 96620 372764 96626
rect 372712 96562 372764 96568
rect 372724 86986 372752 96562
rect 372724 86958 372936 86986
rect 372908 80170 372936 86958
rect 372896 80164 372948 80170
rect 372896 80106 372948 80112
rect 372712 80028 372764 80034
rect 372712 79970 372764 79976
rect 372724 70394 372752 79970
rect 372632 70366 372752 70394
rect 372632 70258 372660 70366
rect 372632 70230 372752 70258
rect 372724 51082 372752 70230
rect 372632 51054 372752 51082
rect 372632 50946 372660 51054
rect 372632 50918 372752 50946
rect 372724 36122 372752 50918
rect 372724 36094 372844 36122
rect 372816 21978 372844 36094
rect 372816 21950 373028 21978
rect 371148 4140 371200 4146
rect 371148 4082 371200 4088
rect 371608 3936 371660 3942
rect 371608 3878 371660 3884
rect 370504 3188 370556 3194
rect 370504 3130 370556 3136
rect 371620 480 371648 3878
rect 372804 3868 372856 3874
rect 372804 3810 372856 3816
rect 372816 480 372844 3810
rect 373000 3126 373028 21950
rect 373920 3874 373948 337486
rect 374012 4078 374040 340068
rect 374472 337482 374500 340068
rect 374748 340054 375038 340082
rect 375498 340054 375696 340082
rect 374460 337476 374512 337482
rect 374460 337418 374512 337424
rect 374748 333198 374776 340054
rect 375288 337544 375340 337550
rect 375288 337486 375340 337492
rect 374092 333192 374144 333198
rect 374092 333134 374144 333140
rect 374736 333192 374788 333198
rect 374736 333134 374788 333140
rect 374000 4072 374052 4078
rect 374000 4014 374052 4020
rect 373908 3868 373960 3874
rect 373908 3810 373960 3816
rect 374000 3800 374052 3806
rect 374000 3742 374052 3748
rect 372988 3120 373040 3126
rect 372988 3062 373040 3068
rect 374012 480 374040 3742
rect 374104 2990 374132 333134
rect 375300 3806 375328 337486
rect 375288 3800 375340 3806
rect 375288 3742 375340 3748
rect 375196 3732 375248 3738
rect 375196 3674 375248 3680
rect 374092 2984 374144 2990
rect 374092 2926 374144 2932
rect 375208 480 375236 3674
rect 375668 3398 375696 340054
rect 375944 337754 375972 340068
rect 376036 340054 376510 340082
rect 375932 337748 375984 337754
rect 375932 337690 375984 337696
rect 376036 336954 376064 340054
rect 375852 336926 376064 336954
rect 375852 321638 375880 336926
rect 376956 336802 376984 340068
rect 377416 337822 377444 340068
rect 377508 340054 377890 340082
rect 377404 337816 377456 337822
rect 377404 337758 377456 337764
rect 376024 336796 376076 336802
rect 376024 336738 376076 336744
rect 376944 336796 376996 336802
rect 376944 336738 376996 336744
rect 375840 321632 375892 321638
rect 375840 321574 375892 321580
rect 375932 321428 375984 321434
rect 375932 321370 375984 321376
rect 375944 289882 375972 321370
rect 375840 289876 375892 289882
rect 375840 289818 375892 289824
rect 375932 289876 375984 289882
rect 375932 289818 375984 289824
rect 375852 280158 375880 289818
rect 375840 280152 375892 280158
rect 375840 280094 375892 280100
rect 375840 270564 375892 270570
rect 375840 270506 375892 270512
rect 375852 260846 375880 270506
rect 375840 260840 375892 260846
rect 375840 260782 375892 260788
rect 375840 251252 375892 251258
rect 375840 251194 375892 251200
rect 375852 241466 375880 251194
rect 375840 241460 375892 241466
rect 375840 241402 375892 241408
rect 375840 231872 375892 231878
rect 375840 231814 375892 231820
rect 375852 222154 375880 231814
rect 375840 222148 375892 222154
rect 375840 222090 375892 222096
rect 375840 212560 375892 212566
rect 375840 212502 375892 212508
rect 375852 202842 375880 212502
rect 375840 202836 375892 202842
rect 375840 202778 375892 202784
rect 375840 193248 375892 193254
rect 375840 193190 375892 193196
rect 375852 183530 375880 193190
rect 375840 183524 375892 183530
rect 375840 183466 375892 183472
rect 375840 173936 375892 173942
rect 375840 173878 375892 173884
rect 375852 164218 375880 173878
rect 375840 164212 375892 164218
rect 375840 164154 375892 164160
rect 375840 154624 375892 154630
rect 375840 154566 375892 154572
rect 375852 144906 375880 154566
rect 375840 144900 375892 144906
rect 375840 144842 375892 144848
rect 375840 135312 375892 135318
rect 375840 135254 375892 135260
rect 375852 118810 375880 135254
rect 375760 118782 375880 118810
rect 375760 118674 375788 118782
rect 375760 118646 375880 118674
rect 375852 106282 375880 118646
rect 375840 106276 375892 106282
rect 375840 106218 375892 106224
rect 375840 97844 375892 97850
rect 375840 97786 375892 97792
rect 375852 80034 375880 97786
rect 375840 80028 375892 80034
rect 375840 79970 375892 79976
rect 375932 79960 375984 79966
rect 375932 79902 375984 79908
rect 375944 60874 375972 79902
rect 375852 60846 375972 60874
rect 375852 60738 375880 60846
rect 375760 60710 375880 60738
rect 375760 60602 375788 60710
rect 375760 60574 375880 60602
rect 375852 41426 375880 60574
rect 375760 41398 375880 41426
rect 375760 41290 375788 41398
rect 375760 41262 375880 41290
rect 375852 22114 375880 41262
rect 375760 22086 375880 22114
rect 375760 21978 375788 22086
rect 375760 21950 375880 21978
rect 375656 3392 375708 3398
rect 375656 3334 375708 3340
rect 375852 2854 375880 21950
rect 376036 3262 376064 336738
rect 377508 335594 377536 340054
rect 378048 337000 378100 337006
rect 378048 336942 378100 336948
rect 377680 336796 377732 336802
rect 377680 336738 377732 336744
rect 377140 335566 377536 335594
rect 377140 321638 377168 335566
rect 377692 331242 377720 336738
rect 377416 331214 377720 331242
rect 377128 321632 377180 321638
rect 377128 321574 377180 321580
rect 377220 321428 377272 321434
rect 377220 321370 377272 321376
rect 377232 289882 377260 321370
rect 377128 289876 377180 289882
rect 377128 289818 377180 289824
rect 377220 289876 377272 289882
rect 377220 289818 377272 289824
rect 377140 280158 377168 289818
rect 377128 280152 377180 280158
rect 377128 280094 377180 280100
rect 377128 270564 377180 270570
rect 377128 270506 377180 270512
rect 377140 260846 377168 270506
rect 377128 260840 377180 260846
rect 377128 260782 377180 260788
rect 377128 251252 377180 251258
rect 377128 251194 377180 251200
rect 377140 241505 377168 251194
rect 376942 241496 376998 241505
rect 376942 241431 376998 241440
rect 377126 241496 377182 241505
rect 377126 241431 377182 241440
rect 376956 231878 376984 241431
rect 376944 231872 376996 231878
rect 376944 231814 376996 231820
rect 377128 231872 377180 231878
rect 377128 231814 377180 231820
rect 377140 222193 377168 231814
rect 376942 222184 376998 222193
rect 376942 222119 376998 222128
rect 377126 222184 377182 222193
rect 377126 222119 377182 222128
rect 376956 212566 376984 222119
rect 376944 212560 376996 212566
rect 376944 212502 376996 212508
rect 377128 212560 377180 212566
rect 377128 212502 377180 212508
rect 377140 202881 377168 212502
rect 376942 202872 376998 202881
rect 376942 202807 376998 202816
rect 377126 202872 377182 202881
rect 377126 202807 377182 202816
rect 376956 193254 376984 202807
rect 376944 193248 376996 193254
rect 376944 193190 376996 193196
rect 377128 193248 377180 193254
rect 377128 193190 377180 193196
rect 377140 183569 377168 193190
rect 376942 183560 376998 183569
rect 376942 183495 376998 183504
rect 377126 183560 377182 183569
rect 377126 183495 377182 183504
rect 376956 173942 376984 183495
rect 376944 173936 376996 173942
rect 376944 173878 376996 173884
rect 377128 173936 377180 173942
rect 377128 173878 377180 173884
rect 377140 164218 377168 173878
rect 376944 164212 376996 164218
rect 376944 164154 376996 164160
rect 377128 164212 377180 164218
rect 377128 164154 377180 164160
rect 376956 154601 376984 164154
rect 376942 154592 376998 154601
rect 376942 154527 376998 154536
rect 377126 154592 377182 154601
rect 377126 154527 377182 154536
rect 377140 144906 377168 154527
rect 376944 144900 376996 144906
rect 376944 144842 376996 144848
rect 377128 144900 377180 144906
rect 377128 144842 377180 144848
rect 376956 135289 376984 144842
rect 376942 135280 376998 135289
rect 376942 135215 376998 135224
rect 377126 135280 377182 135289
rect 377126 135215 377182 135224
rect 377140 118726 377168 135215
rect 377128 118720 377180 118726
rect 377128 118662 377180 118668
rect 377128 118584 377180 118590
rect 377128 118526 377180 118532
rect 377140 115938 377168 118526
rect 377128 115932 377180 115938
rect 377128 115874 377180 115880
rect 376666 110800 376722 110809
rect 376666 110735 376722 110744
rect 376680 110702 376708 110735
rect 376668 110696 376720 110702
rect 376668 110638 376720 110644
rect 377036 106344 377088 106350
rect 377088 106292 377168 106298
rect 377036 106286 377168 106292
rect 377048 106282 377168 106286
rect 377048 106276 377180 106282
rect 377048 106270 377128 106276
rect 377128 106218 377180 106224
rect 377128 99340 377180 99346
rect 377128 99282 377180 99288
rect 376758 87136 376814 87145
rect 376758 87071 376760 87080
rect 376812 87071 376814 87080
rect 376760 87042 376812 87048
rect 377140 80034 377168 99282
rect 377128 80028 377180 80034
rect 377128 79970 377180 79976
rect 377220 79960 377272 79966
rect 377220 79902 377272 79908
rect 376666 76256 376722 76265
rect 376666 76191 376668 76200
rect 376720 76191 376722 76200
rect 376668 76162 376720 76168
rect 377232 60874 377260 79902
rect 377140 60846 377260 60874
rect 377140 60738 377168 60846
rect 377048 60710 377168 60738
rect 377048 60602 377076 60710
rect 377048 60574 377168 60602
rect 377140 41342 377168 60574
rect 377128 41336 377180 41342
rect 377128 41278 377180 41284
rect 377036 38752 377088 38758
rect 377088 38700 377168 38706
rect 377036 38694 377168 38700
rect 377048 38678 377168 38694
rect 377140 32026 377168 38678
rect 377128 32020 377180 32026
rect 377128 31962 377180 31968
rect 377312 32020 377364 32026
rect 377312 31962 377364 31968
rect 377324 29073 377352 31962
rect 377126 29064 377182 29073
rect 377048 29022 377126 29050
rect 377048 22166 377076 29022
rect 377126 28999 377182 29008
rect 377310 29064 377366 29073
rect 377310 28999 377366 29008
rect 377036 22160 377088 22166
rect 377036 22102 377088 22108
rect 377128 22024 377180 22030
rect 377128 21966 377180 21972
rect 377140 17950 377168 21966
rect 377128 17944 377180 17950
rect 377128 17886 377180 17892
rect 376760 8356 376812 8362
rect 376760 8298 376812 8304
rect 376772 4078 376800 8298
rect 376760 4072 376812 4078
rect 376760 4014 376812 4020
rect 377416 3670 377444 331214
rect 378060 4146 378088 336942
rect 378428 336802 378456 340068
rect 378888 337890 378916 340068
rect 379348 338026 379376 340068
rect 379716 340054 379914 340082
rect 379336 338020 379388 338026
rect 379336 337962 379388 337968
rect 378876 337884 378928 337890
rect 378876 337826 378928 337832
rect 378416 336796 378468 336802
rect 378416 336738 378468 336744
rect 377588 4140 377640 4146
rect 377588 4082 377640 4088
rect 378048 4140 378100 4146
rect 378048 4082 378100 4088
rect 378784 4140 378836 4146
rect 378784 4082 378836 4088
rect 377404 3664 377456 3670
rect 377404 3606 377456 3612
rect 376024 3256 376076 3262
rect 376024 3198 376076 3204
rect 376392 3052 376444 3058
rect 376392 2994 376444 3000
rect 375840 2848 375892 2854
rect 375840 2790 375892 2796
rect 376404 480 376432 2994
rect 377600 480 377628 4082
rect 378796 480 378824 4082
rect 379716 3466 379744 340054
rect 380164 337748 380216 337754
rect 380164 337690 380216 337696
rect 380176 4962 380204 337690
rect 380360 337346 380388 340068
rect 380820 337686 380848 340068
rect 381372 337754 381400 340068
rect 381360 337748 381412 337754
rect 381360 337690 381412 337696
rect 381544 337748 381596 337754
rect 381544 337690 381596 337696
rect 380808 337680 380860 337686
rect 380808 337622 380860 337628
rect 380348 337340 380400 337346
rect 380348 337282 380400 337288
rect 380808 336932 380860 336938
rect 380808 336874 380860 336880
rect 380164 4956 380216 4962
rect 380164 4898 380216 4904
rect 380820 3534 380848 336874
rect 381556 5098 381584 337690
rect 381832 337482 381860 340068
rect 382292 338026 382320 340068
rect 382280 338020 382332 338026
rect 382280 337962 382332 337968
rect 382844 337754 382872 340068
rect 382832 337748 382884 337754
rect 382832 337690 382884 337696
rect 383304 337618 383332 340068
rect 383292 337612 383344 337618
rect 383292 337554 383344 337560
rect 383764 337550 383792 340068
rect 383856 340054 384330 340082
rect 383752 337544 383804 337550
rect 383752 337486 383804 337492
rect 381820 337476 381872 337482
rect 381820 337418 381872 337424
rect 382188 337408 382240 337414
rect 382188 337350 382240 337356
rect 381636 336864 381688 336870
rect 381636 336806 381688 336812
rect 381544 5092 381596 5098
rect 381544 5034 381596 5040
rect 379980 3528 380032 3534
rect 379980 3470 380032 3476
rect 380808 3528 380860 3534
rect 380808 3470 380860 3476
rect 381176 3528 381228 3534
rect 381176 3470 381228 3476
rect 379704 3460 379756 3466
rect 379704 3402 379756 3408
rect 379992 480 380020 3470
rect 381188 480 381216 3470
rect 381648 3058 381676 336806
rect 382200 3534 382228 337350
rect 383568 4072 383620 4078
rect 383568 4014 383620 4020
rect 382188 3528 382240 3534
rect 382188 3470 382240 3476
rect 382372 3460 382424 3466
rect 382372 3402 382424 3408
rect 381636 3052 381688 3058
rect 381636 2994 381688 3000
rect 382384 480 382412 3402
rect 383580 480 383608 4014
rect 383856 3738 383884 340054
rect 384304 337680 384356 337686
rect 384304 337622 384356 337628
rect 384316 4078 384344 337622
rect 384776 336870 384804 340068
rect 384948 337748 385000 337754
rect 384948 337690 385000 337696
rect 384764 336864 384816 336870
rect 384764 336806 384816 336812
rect 384304 4072 384356 4078
rect 384304 4014 384356 4020
rect 383844 3732 383896 3738
rect 383844 3674 383896 3680
rect 384960 3346 384988 337690
rect 385236 337006 385264 340068
rect 385328 340054 385802 340082
rect 385224 337000 385276 337006
rect 385224 336942 385276 336948
rect 385132 16856 385184 16862
rect 385130 16824 385132 16833
rect 385184 16824 385186 16833
rect 385130 16759 385186 16768
rect 385328 4146 385356 340054
rect 386248 336938 386276 340068
rect 386708 337414 386736 340068
rect 386696 337408 386748 337414
rect 386696 337350 386748 337356
rect 386800 337226 386828 340190
rect 387720 337686 387748 340068
rect 388180 337754 388208 340068
rect 388444 337884 388496 337890
rect 388444 337826 388496 337832
rect 388168 337748 388220 337754
rect 388168 337690 388220 337696
rect 387708 337680 387760 337686
rect 387708 337622 387760 337628
rect 387064 337476 387116 337482
rect 387064 337418 387116 337424
rect 386616 337198 386828 337226
rect 386236 336932 386288 336938
rect 386236 336874 386288 336880
rect 386236 87100 386288 87106
rect 386236 87042 386288 87048
rect 386420 87100 386472 87106
rect 386420 87042 386472 87048
rect 386248 87009 386276 87042
rect 386432 87009 386460 87042
rect 386234 87000 386290 87009
rect 386234 86935 386290 86944
rect 386418 87000 386474 87009
rect 386418 86935 386474 86944
rect 386418 76528 386474 76537
rect 386418 76463 386474 76472
rect 386432 76265 386460 76463
rect 386418 76256 386474 76265
rect 386418 76191 386474 76200
rect 385316 4140 385368 4146
rect 385316 4082 385368 4088
rect 386616 3466 386644 337198
rect 386604 3460 386656 3466
rect 386604 3402 386656 3408
rect 384684 3318 384988 3346
rect 384684 480 384712 3318
rect 387076 2922 387104 337418
rect 388260 3528 388312 3534
rect 388260 3470 388312 3476
rect 385868 2916 385920 2922
rect 385868 2858 385920 2864
rect 387064 2916 387116 2922
rect 387064 2858 387116 2864
rect 385880 480 385908 2858
rect 387064 2780 387116 2786
rect 387064 2722 387116 2728
rect 387076 480 387104 2722
rect 388272 480 388300 3470
rect 388456 2854 388484 337826
rect 388732 337482 388760 340068
rect 389192 337890 389220 340068
rect 389284 340054 389666 340082
rect 389180 337884 389232 337890
rect 389180 337826 389232 337832
rect 389284 337770 389312 340054
rect 389100 337742 389312 337770
rect 388720 337476 388772 337482
rect 388720 337418 388772 337424
rect 388994 251152 389050 251161
rect 388994 251087 389050 251096
rect 389008 241602 389036 251087
rect 388996 241596 389048 241602
rect 388996 241538 389048 241544
rect 388994 48240 389050 48249
rect 388994 48175 389050 48184
rect 389008 41410 389036 48175
rect 388996 41404 389048 41410
rect 388996 41346 389048 41352
rect 389100 3534 389128 337742
rect 389744 335594 389772 340190
rect 390664 335714 390692 340068
rect 390756 340054 391138 340082
rect 391690 340054 391888 340082
rect 390652 335708 390704 335714
rect 390652 335650 390704 335656
rect 390756 335594 390784 340054
rect 391860 336818 391888 340054
rect 392136 336938 392164 340068
rect 392124 336932 392176 336938
rect 392124 336874 392176 336880
rect 391860 336790 392164 336818
rect 389284 335566 389772 335594
rect 390572 335566 390784 335594
rect 389284 331226 389312 335566
rect 389272 331220 389324 331226
rect 389272 331162 389324 331168
rect 389456 331220 389508 331226
rect 389456 331162 389508 331168
rect 389468 328438 389496 331162
rect 389456 328432 389508 328438
rect 389456 328374 389508 328380
rect 389548 318844 389600 318850
rect 389548 318786 389600 318792
rect 389560 309194 389588 318786
rect 389364 309188 389416 309194
rect 389364 309130 389416 309136
rect 389548 309188 389600 309194
rect 389548 309130 389600 309136
rect 389376 309058 389404 309130
rect 389364 309052 389416 309058
rect 389364 308994 389416 309000
rect 389272 299532 389324 299538
rect 389272 299474 389324 299480
rect 389284 292618 389312 299474
rect 389284 292590 389496 292618
rect 389468 289814 389496 292590
rect 389456 289808 389508 289814
rect 389456 289750 389508 289756
rect 389364 280220 389416 280226
rect 389364 280162 389416 280168
rect 389376 273306 389404 280162
rect 389376 273278 389496 273306
rect 389468 270502 389496 273278
rect 389456 270496 389508 270502
rect 389456 270438 389508 270444
rect 389364 260908 389416 260914
rect 389364 260850 389416 260856
rect 389376 251258 389404 260850
rect 389180 251252 389232 251258
rect 389180 251194 389232 251200
rect 389364 251252 389416 251258
rect 389364 251194 389416 251200
rect 389192 251161 389220 251194
rect 389178 251152 389234 251161
rect 389178 251087 389234 251096
rect 389272 241596 389324 241602
rect 389272 241538 389324 241544
rect 389284 241466 389312 241538
rect 389272 241460 389324 241466
rect 389272 241402 389324 241408
rect 389456 234660 389508 234666
rect 389456 234602 389508 234608
rect 389468 231849 389496 234602
rect 389270 231840 389326 231849
rect 389270 231775 389326 231784
rect 389454 231840 389510 231849
rect 389454 231775 389510 231784
rect 389284 222222 389312 231775
rect 389272 222216 389324 222222
rect 389272 222158 389324 222164
rect 389548 222216 389600 222222
rect 389548 222158 389600 222164
rect 389560 215422 389588 222158
rect 389548 215416 389600 215422
rect 389548 215358 389600 215364
rect 389456 215280 389508 215286
rect 389456 215222 389508 215228
rect 389468 212537 389496 215222
rect 389270 212528 389326 212537
rect 389270 212463 389326 212472
rect 389454 212528 389510 212537
rect 389454 212463 389510 212472
rect 389284 202910 389312 212463
rect 389272 202904 389324 202910
rect 389272 202846 389324 202852
rect 389548 202904 389600 202910
rect 389548 202846 389600 202852
rect 389560 196110 389588 202846
rect 389548 196104 389600 196110
rect 389548 196046 389600 196052
rect 389456 195968 389508 195974
rect 389456 195910 389508 195916
rect 389468 193225 389496 195910
rect 389270 193216 389326 193225
rect 389270 193151 389326 193160
rect 389454 193216 389510 193225
rect 389454 193151 389510 193160
rect 389284 183598 389312 193151
rect 389272 183592 389324 183598
rect 389272 183534 389324 183540
rect 389548 183592 389600 183598
rect 389548 183534 389600 183540
rect 389560 176798 389588 183534
rect 389548 176792 389600 176798
rect 389548 176734 389600 176740
rect 389456 176656 389508 176662
rect 389456 176598 389508 176604
rect 389468 154562 389496 176598
rect 389456 154556 389508 154562
rect 389456 154498 389508 154504
rect 389640 154556 389692 154562
rect 389640 154498 389692 154504
rect 389652 144945 389680 154498
rect 389362 144936 389418 144945
rect 389362 144871 389418 144880
rect 389638 144936 389694 144945
rect 389638 144871 389694 144880
rect 389376 138038 389404 144871
rect 389364 138032 389416 138038
rect 389364 137974 389416 137980
rect 389456 137964 389508 137970
rect 389456 137906 389508 137912
rect 389468 133890 389496 137906
rect 389456 133884 389508 133890
rect 389456 133826 389508 133832
rect 389180 122868 389232 122874
rect 389180 122810 389232 122816
rect 389192 122754 389220 122810
rect 389192 122726 389312 122754
rect 389284 118833 389312 122726
rect 389270 118824 389326 118833
rect 389270 118759 389326 118768
rect 389454 108896 389510 108905
rect 389454 108831 389510 108840
rect 389468 99210 389496 108831
rect 389456 99204 389508 99210
rect 389456 99146 389508 99152
rect 389364 87916 389416 87922
rect 389364 87858 389416 87864
rect 389376 80102 389404 87858
rect 389364 80096 389416 80102
rect 389364 80038 389416 80044
rect 389456 79960 389508 79966
rect 389456 79902 389508 79908
rect 389468 77246 389496 79902
rect 389456 77240 389508 77246
rect 389456 77182 389508 77188
rect 389364 67652 389416 67658
rect 389364 67594 389416 67600
rect 389376 60738 389404 67594
rect 389192 60710 389404 60738
rect 389192 57934 389220 60710
rect 389180 57928 389232 57934
rect 389180 57870 389232 57876
rect 389272 48340 389324 48346
rect 389272 48282 389324 48288
rect 389178 48240 389234 48249
rect 389284 48226 389312 48282
rect 389234 48198 389312 48226
rect 389178 48175 389234 48184
rect 389364 41404 389416 41410
rect 389364 41346 389416 41352
rect 389376 31754 389404 41346
rect 389364 31748 389416 31754
rect 389364 31690 389416 31696
rect 389548 31748 389600 31754
rect 389548 31690 389600 31696
rect 389560 28966 389588 31690
rect 389548 28960 389600 28966
rect 389548 28902 389600 28908
rect 389456 19372 389508 19378
rect 389456 19314 389508 19320
rect 389468 12458 389496 19314
rect 389468 12430 389588 12458
rect 389560 9654 389588 12430
rect 389548 9648 389600 9654
rect 389548 9590 389600 9596
rect 390572 4146 390600 335566
rect 390652 335504 390704 335510
rect 390652 335446 390704 335452
rect 390560 4140 390612 4146
rect 390560 4082 390612 4088
rect 389088 3528 389140 3534
rect 389088 3470 389140 3476
rect 388444 2848 388496 2854
rect 388444 2790 388496 2796
rect 389456 604 389508 610
rect 389456 546 389508 552
rect 389468 480 389496 546
rect 390664 480 390692 335446
rect 392136 12442 392164 336790
rect 393056 331242 393084 340190
rect 393162 340054 393268 340082
rect 393056 331214 393176 331242
rect 392124 12436 392176 12442
rect 392124 12378 392176 12384
rect 393044 12436 393096 12442
rect 393044 12378 393096 12384
rect 391848 4140 391900 4146
rect 391848 4082 391900 4088
rect 391860 480 391888 4082
rect 393056 480 393084 12378
rect 393148 4146 393176 331214
rect 393136 4140 393188 4146
rect 393136 4082 393188 4088
rect 393240 4078 393268 340054
rect 393608 337074 393636 340068
rect 394082 340054 394556 340082
rect 393596 337068 393648 337074
rect 393596 337010 393648 337016
rect 393596 336932 393648 336938
rect 393596 336874 393648 336880
rect 393228 4072 393280 4078
rect 393228 4014 393280 4020
rect 393608 610 393636 336874
rect 394528 3330 394556 340054
rect 394516 3324 394568 3330
rect 394516 3266 394568 3272
rect 394620 3262 394648 340068
rect 395080 336802 395108 340068
rect 395554 340054 395936 340082
rect 395068 336796 395120 336802
rect 395068 336738 395120 336744
rect 395908 87242 395936 340054
rect 396092 336870 396120 340068
rect 396080 336864 396132 336870
rect 396080 336806 396132 336812
rect 396552 336802 396580 340068
rect 397012 337482 397040 340068
rect 397472 338026 397500 340068
rect 397460 338020 397512 338026
rect 397460 337962 397512 337968
rect 398024 337618 398052 340068
rect 398012 337612 398064 337618
rect 398012 337554 398064 337560
rect 397000 337476 397052 337482
rect 397000 337418 397052 337424
rect 398484 337346 398512 340068
rect 398944 337686 398972 340068
rect 399496 337754 399524 340068
rect 399970 340054 400076 340082
rect 399484 337748 399536 337754
rect 399484 337690 399536 337696
rect 398932 337680 398984 337686
rect 398932 337622 398984 337628
rect 399484 337612 399536 337618
rect 399484 337554 399536 337560
rect 398472 337340 398524 337346
rect 398472 337282 398524 337288
rect 397460 337068 397512 337074
rect 397460 337010 397512 337016
rect 395988 336796 396040 336802
rect 395988 336738 396040 336744
rect 396540 336796 396592 336802
rect 396540 336738 396592 336744
rect 396000 87242 396028 336738
rect 395896 87236 395948 87242
rect 395896 87178 395948 87184
rect 395988 87236 396040 87242
rect 395988 87178 396040 87184
rect 395986 87136 396042 87145
rect 395816 87106 395986 87122
rect 395804 87100 395986 87106
rect 395856 87094 395986 87100
rect 395986 87071 396042 87080
rect 395804 87042 395856 87048
rect 395896 87032 395948 87038
rect 395896 86974 395948 86980
rect 395988 87032 396040 87038
rect 395988 86974 396040 86980
rect 395908 17218 395936 86974
rect 395816 17190 395936 17218
rect 396000 17202 396028 86974
rect 396078 76120 396134 76129
rect 396078 76055 396080 76064
rect 396132 76055 396134 76064
rect 396080 76026 396132 76032
rect 396080 40248 396132 40254
rect 396078 40216 396080 40225
rect 396132 40216 396134 40225
rect 396078 40151 396134 40160
rect 395988 17196 396040 17202
rect 395816 14498 395844 17190
rect 395988 17138 396040 17144
rect 395894 17096 395950 17105
rect 395894 17031 395950 17040
rect 395908 16862 395936 17031
rect 395988 16992 396040 16998
rect 395988 16934 396040 16940
rect 395896 16856 395948 16862
rect 395896 16798 395948 16804
rect 395816 14470 395936 14498
rect 395436 4140 395488 4146
rect 395436 4082 395488 4088
rect 394608 3256 394660 3262
rect 394608 3198 394660 3204
rect 393596 604 393648 610
rect 393596 546 393648 552
rect 394240 604 394292 610
rect 394240 546 394292 552
rect 394252 480 394280 546
rect 395448 480 395476 4082
rect 395908 3466 395936 14470
rect 396000 3534 396028 16934
rect 396632 4072 396684 4078
rect 396632 4014 396684 4020
rect 395988 3528 396040 3534
rect 395988 3470 396040 3476
rect 395896 3460 395948 3466
rect 395896 3402 395948 3408
rect 396644 480 396672 4014
rect 397472 610 397500 337010
rect 398104 336864 398156 336870
rect 398104 336806 398156 336812
rect 398116 4146 398144 336806
rect 398196 336796 398248 336802
rect 398196 336738 398248 336744
rect 398104 4140 398156 4146
rect 398104 4082 398156 4088
rect 398208 2990 398236 336738
rect 399390 76120 399446 76129
rect 399390 76055 399392 76064
rect 399444 76055 399446 76064
rect 399392 76026 399444 76032
rect 399024 40248 399076 40254
rect 399022 40216 399024 40225
rect 399076 40216 399078 40225
rect 399022 40151 399078 40160
rect 398746 16688 398802 16697
rect 398930 16688 398986 16697
rect 398802 16646 398930 16674
rect 398746 16623 398802 16632
rect 398930 16623 398986 16632
rect 399496 3806 399524 337554
rect 399484 3800 399536 3806
rect 399484 3742 399536 3748
rect 400048 3670 400076 340054
rect 400416 337958 400444 340068
rect 400404 337952 400456 337958
rect 400404 337894 400456 337900
rect 400128 337748 400180 337754
rect 400128 337690 400180 337696
rect 400140 3738 400168 337690
rect 400968 337414 400996 340068
rect 400956 337408 401008 337414
rect 400956 337350 401008 337356
rect 401428 336938 401456 340068
rect 401888 337210 401916 340068
rect 402440 337754 402468 340068
rect 402808 340054 402914 340082
rect 402428 337748 402480 337754
rect 402428 337690 402480 337696
rect 402244 337408 402296 337414
rect 402244 337350 402296 337356
rect 401876 337204 401928 337210
rect 401876 337146 401928 337152
rect 401416 336932 401468 336938
rect 401416 336874 401468 336880
rect 400128 3732 400180 3738
rect 400128 3674 400180 3680
rect 400036 3664 400088 3670
rect 400036 3606 400088 3612
rect 402256 3602 402284 337350
rect 402244 3596 402296 3602
rect 402244 3538 402296 3544
rect 402808 3534 402836 340054
rect 403360 337754 403388 340068
rect 403926 340054 404308 340082
rect 403624 338020 403676 338026
rect 403624 337962 403676 337968
rect 402888 337748 402940 337754
rect 402888 337690 402940 337696
rect 403348 337748 403400 337754
rect 403348 337690 403400 337696
rect 402900 4010 402928 337690
rect 402888 4004 402940 4010
rect 402888 3946 402940 3952
rect 401324 3528 401376 3534
rect 401324 3470 401376 3476
rect 402796 3528 402848 3534
rect 402796 3470 402848 3476
rect 399024 3324 399076 3330
rect 399024 3266 399076 3272
rect 398196 2984 398248 2990
rect 398196 2926 398248 2932
rect 397460 604 397512 610
rect 397460 546 397512 552
rect 397828 604 397880 610
rect 397828 546 397880 552
rect 397840 480 397868 546
rect 399036 480 399064 3266
rect 400220 3256 400272 3262
rect 400220 3198 400272 3204
rect 400232 480 400260 3198
rect 401336 480 401364 3470
rect 403636 3466 403664 337962
rect 403716 4140 403768 4146
rect 403716 4082 403768 4088
rect 402520 3460 402572 3466
rect 402520 3402 402572 3408
rect 403624 3460 403676 3466
rect 403624 3402 403676 3408
rect 402532 480 402560 3402
rect 403728 480 403756 4082
rect 404280 3398 404308 340054
rect 404372 337822 404400 340068
rect 404832 337890 404860 340068
rect 405398 340054 405688 340082
rect 404820 337884 404872 337890
rect 404820 337826 404872 337832
rect 404360 337816 404412 337822
rect 404360 337758 404412 337764
rect 405004 336932 405056 336938
rect 405004 336874 405056 336880
rect 404268 3392 404320 3398
rect 404268 3334 404320 3340
rect 405016 3330 405044 336874
rect 405004 3324 405056 3330
rect 405004 3266 405056 3272
rect 405660 3126 405688 340054
rect 405844 337550 405872 340068
rect 406304 338094 406332 340068
rect 406870 340054 407068 340082
rect 406292 338088 406344 338094
rect 406292 338030 406344 338036
rect 406384 337680 406436 337686
rect 406384 337622 406436 337628
rect 405832 337544 405884 337550
rect 405832 337486 405884 337492
rect 405924 337476 405976 337482
rect 405924 337418 405976 337424
rect 405648 3120 405700 3126
rect 405648 3062 405700 3068
rect 404912 2984 404964 2990
rect 404912 2926 404964 2932
rect 404924 480 404952 2926
rect 405936 610 405964 337418
rect 406396 3058 406424 337622
rect 407040 3194 407068 340054
rect 407316 337618 407344 340068
rect 407304 337612 407356 337618
rect 407304 337554 407356 337560
rect 407776 337414 407804 340068
rect 408342 340054 408448 340082
rect 408802 340054 409092 340082
rect 407764 337408 407816 337414
rect 407764 337350 407816 337356
rect 408420 5438 408448 340054
rect 408776 337340 408828 337346
rect 408776 337282 408828 337288
rect 408408 5432 408460 5438
rect 408408 5374 408460 5380
rect 408500 3800 408552 3806
rect 408500 3742 408552 3748
rect 407304 3460 407356 3466
rect 407304 3402 407356 3408
rect 407028 3188 407080 3194
rect 407028 3130 407080 3136
rect 406384 3052 406436 3058
rect 406384 2994 406436 3000
rect 405924 604 405976 610
rect 405924 546 405976 552
rect 406108 604 406160 610
rect 406108 546 406160 552
rect 406120 480 406148 546
rect 407316 480 407344 3402
rect 408512 480 408540 3742
rect 408788 2938 408816 337282
rect 409064 336938 409092 340054
rect 409144 337408 409196 337414
rect 409144 337350 409196 337356
rect 409052 336932 409104 336938
rect 409052 336874 409104 336880
rect 409156 3262 409184 337350
rect 409248 337346 409276 340068
rect 409236 337340 409288 337346
rect 409236 337282 409288 337288
rect 409800 3398 409828 340068
rect 410260 337754 410288 340068
rect 410734 340054 411208 340082
rect 410248 337748 410300 337754
rect 410248 337690 410300 337696
rect 411076 337748 411128 337754
rect 411076 337690 411128 337696
rect 411088 3806 411116 337690
rect 411180 4078 411208 340054
rect 411272 337686 411300 340068
rect 411746 340054 412128 340082
rect 412206 340054 412588 340082
rect 412100 337770 412128 340054
rect 412100 337742 412496 337770
rect 411260 337680 411312 337686
rect 411260 337622 411312 337628
rect 412364 337680 412416 337686
rect 412364 337622 412416 337628
rect 412376 5370 412404 337622
rect 412364 5364 412416 5370
rect 412364 5306 412416 5312
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 412468 3942 412496 337742
rect 412456 3936 412508 3942
rect 412456 3878 412508 3884
rect 411076 3800 411128 3806
rect 411076 3742 411128 3748
rect 412560 3738 412588 340054
rect 412744 337006 412772 340068
rect 413218 340054 413600 340082
rect 413284 337952 413336 337958
rect 413284 337894 413336 337900
rect 412732 337000 412784 337006
rect 412732 336942 412784 336948
rect 412088 3732 412140 3738
rect 412088 3674 412140 3680
rect 412548 3732 412600 3738
rect 412548 3674 412600 3680
rect 409788 3392 409840 3398
rect 409788 3334 409840 3340
rect 409144 3256 409196 3262
rect 409144 3198 409196 3204
rect 410892 3052 410944 3058
rect 410892 2994 410944 3000
rect 408788 2910 409736 2938
rect 409708 480 409736 2910
rect 410904 480 410932 2994
rect 412100 480 412128 3674
rect 413192 3664 413244 3670
rect 413192 3606 413244 3612
rect 413204 3346 413232 3606
rect 413296 3534 413324 337894
rect 413572 337736 413600 340054
rect 413664 337958 413692 340068
rect 413652 337952 413704 337958
rect 413652 337894 413704 337900
rect 414216 337754 414244 340068
rect 414676 338026 414704 340068
rect 414664 338020 414716 338026
rect 414664 337962 414716 337968
rect 414204 337748 414256 337754
rect 413572 337708 413968 337736
rect 413836 337000 413888 337006
rect 413836 336942 413888 336948
rect 413848 5302 413876 336942
rect 413836 5296 413888 5302
rect 413836 5238 413888 5244
rect 413940 3874 413968 337708
rect 414204 337690 414256 337696
rect 415136 337142 415164 340068
rect 415596 337754 415624 340068
rect 416148 337822 416176 340068
rect 416136 337816 416188 337822
rect 416136 337758 416188 337764
rect 415308 337748 415360 337754
rect 415308 337690 415360 337696
rect 415584 337748 415636 337754
rect 415584 337690 415636 337696
rect 416504 337748 416556 337754
rect 416504 337690 416556 337696
rect 415124 337136 415176 337142
rect 415124 337078 415176 337084
rect 414018 110664 414074 110673
rect 414018 110599 414020 110608
rect 414072 110599 414074 110608
rect 414020 110570 414072 110576
rect 414020 63776 414072 63782
rect 414018 63744 414020 63753
rect 414072 63744 414074 63753
rect 414018 63679 414074 63688
rect 415320 5234 415348 337690
rect 415308 5228 415360 5234
rect 415308 5170 415360 5176
rect 416516 5166 416544 337690
rect 416504 5160 416556 5166
rect 416504 5102 416556 5108
rect 413928 3868 413980 3874
rect 413928 3810 413980 3816
rect 415676 3596 415728 3602
rect 415676 3538 415728 3544
rect 413284 3528 413336 3534
rect 413284 3470 413336 3476
rect 414480 3528 414532 3534
rect 414480 3470 414532 3476
rect 413204 3318 413324 3346
rect 413296 480 413324 3318
rect 414492 480 414520 3470
rect 415688 480 415716 3538
rect 416608 2922 416636 340068
rect 416688 337816 416740 337822
rect 416688 337758 416740 337764
rect 416700 3670 416728 337758
rect 417068 337754 417096 340068
rect 417424 338088 417476 338094
rect 417424 338030 417476 338036
rect 417056 337748 417108 337754
rect 417056 337690 417108 337696
rect 416964 337204 417016 337210
rect 416964 337146 417016 337152
rect 416688 3664 416740 3670
rect 416688 3606 416740 3612
rect 416872 3324 416924 3330
rect 416872 3266 416924 3272
rect 416596 2916 416648 2922
rect 416596 2858 416648 2864
rect 416884 480 416912 3266
rect 416976 2666 417004 337146
rect 417436 2990 417464 338030
rect 417620 337890 417648 340068
rect 417608 337884 417660 337890
rect 417608 337826 417660 337832
rect 417976 337748 418028 337754
rect 417976 337690 418028 337696
rect 417884 157616 417936 157622
rect 417882 157584 417884 157593
rect 417936 157584 417938 157593
rect 417882 157519 417938 157528
rect 417882 40216 417938 40225
rect 417882 40151 417884 40160
rect 417936 40151 417938 40160
rect 417884 40122 417936 40128
rect 417884 16856 417936 16862
rect 417882 16824 417884 16833
rect 417936 16824 417938 16833
rect 417882 16759 417938 16768
rect 417988 5098 418016 337690
rect 417976 5092 418028 5098
rect 417976 5034 418028 5040
rect 418080 3602 418108 340068
rect 418540 336802 418568 340068
rect 419092 338094 419120 340068
rect 419080 338088 419132 338094
rect 419080 338030 419132 338036
rect 419552 336802 419580 340068
rect 420012 336870 420040 340068
rect 420564 337958 420592 340068
rect 420184 337952 420236 337958
rect 420184 337894 420236 337900
rect 420552 337952 420604 337958
rect 420552 337894 420604 337900
rect 420000 336864 420052 336870
rect 420000 336806 420052 336812
rect 418528 336796 418580 336802
rect 418528 336738 418580 336744
rect 419448 336796 419500 336802
rect 419448 336738 419500 336744
rect 419540 336796 419592 336802
rect 419540 336738 419592 336744
rect 418252 157616 418304 157622
rect 418250 157584 418252 157593
rect 418304 157584 418306 157593
rect 418250 157519 418306 157528
rect 418896 63776 418948 63782
rect 418894 63744 418896 63753
rect 418948 63744 418950 63753
rect 418894 63679 418950 63688
rect 418250 40216 418306 40225
rect 418250 40151 418252 40160
rect 418304 40151 418306 40160
rect 418252 40122 418304 40128
rect 418252 16856 418304 16862
rect 418250 16824 418252 16833
rect 418304 16824 418306 16833
rect 418250 16759 418306 16768
rect 419460 5030 419488 336738
rect 419448 5024 419500 5030
rect 419448 4966 419500 4972
rect 419172 4004 419224 4010
rect 419172 3946 419224 3952
rect 418068 3596 418120 3602
rect 418068 3538 418120 3544
rect 417424 2984 417476 2990
rect 417424 2926 417476 2932
rect 416976 2638 418016 2666
rect 417988 480 418016 2638
rect 419184 480 419212 3946
rect 420196 3330 420224 337894
rect 420276 337816 420328 337822
rect 420276 337758 420328 337764
rect 420288 4010 420316 337758
rect 421024 337346 421052 340068
rect 421196 337476 421248 337482
rect 421196 337418 421248 337424
rect 421012 337340 421064 337346
rect 421012 337282 421064 337288
rect 420736 336864 420788 336870
rect 420736 336806 420788 336812
rect 420748 4962 420776 336806
rect 420828 336796 420880 336802
rect 420828 336738 420880 336744
rect 420736 4956 420788 4962
rect 420736 4898 420788 4904
rect 420276 4004 420328 4010
rect 420276 3946 420328 3952
rect 420840 3534 420868 336738
rect 421208 319002 421236 337418
rect 421484 336802 421512 340068
rect 422036 337822 422064 340068
rect 422024 337816 422076 337822
rect 422024 337758 422076 337764
rect 421564 337136 421616 337142
rect 421564 337078 421616 337084
rect 421472 336796 421524 336802
rect 421472 336738 421524 336744
rect 421208 318974 421328 319002
rect 421300 318866 421328 318974
rect 421208 318838 421328 318866
rect 421208 317422 421236 318838
rect 421196 317416 421248 317422
rect 421196 317358 421248 317364
rect 421196 307828 421248 307834
rect 421196 307770 421248 307776
rect 421208 298110 421236 307770
rect 421196 298104 421248 298110
rect 421196 298046 421248 298052
rect 421196 288448 421248 288454
rect 421196 288390 421248 288396
rect 421208 278769 421236 288390
rect 421194 278760 421250 278769
rect 421194 278695 421250 278704
rect 421378 278760 421434 278769
rect 421378 278695 421434 278704
rect 421392 269142 421420 278695
rect 421196 269136 421248 269142
rect 421196 269078 421248 269084
rect 421380 269136 421432 269142
rect 421380 269078 421432 269084
rect 421208 259457 421236 269078
rect 421194 259448 421250 259457
rect 421194 259383 421250 259392
rect 421378 259448 421434 259457
rect 421378 259383 421434 259392
rect 421392 249830 421420 259383
rect 421196 249824 421248 249830
rect 421196 249766 421248 249772
rect 421380 249824 421432 249830
rect 421380 249766 421432 249772
rect 421208 241777 421236 249766
rect 421194 241768 421250 241777
rect 421194 241703 421250 241712
rect 421194 241632 421250 241641
rect 421194 241567 421250 241576
rect 421208 240145 421236 241567
rect 421194 240136 421250 240145
rect 421194 240071 421250 240080
rect 421378 240136 421434 240145
rect 421378 240071 421434 240080
rect 421392 230518 421420 240071
rect 421196 230512 421248 230518
rect 421196 230454 421248 230460
rect 421380 230512 421432 230518
rect 421380 230454 421432 230460
rect 421208 220833 421236 230454
rect 421194 220824 421250 220833
rect 421194 220759 421250 220768
rect 421378 220824 421434 220833
rect 421378 220759 421434 220768
rect 421392 202910 421420 220759
rect 421196 202904 421248 202910
rect 421196 202846 421248 202852
rect 421380 202904 421432 202910
rect 421380 202846 421432 202852
rect 421208 201482 421236 202846
rect 421104 201476 421156 201482
rect 421104 201418 421156 201424
rect 421196 201476 421248 201482
rect 421196 201418 421248 201424
rect 421116 196625 421144 201418
rect 421102 196616 421158 196625
rect 421102 196551 421158 196560
rect 421194 183696 421250 183705
rect 421194 183631 421250 183640
rect 421208 182170 421236 183631
rect 421196 182164 421248 182170
rect 421196 182106 421248 182112
rect 421380 182164 421432 182170
rect 421380 182106 421432 182112
rect 421392 172553 421420 182106
rect 421194 172544 421250 172553
rect 421194 172479 421250 172488
rect 421378 172544 421434 172553
rect 421378 172479 421434 172488
rect 421208 162858 421236 172479
rect 421196 162852 421248 162858
rect 421196 162794 421248 162800
rect 421196 153264 421248 153270
rect 421196 153206 421248 153212
rect 421208 143546 421236 153206
rect 421196 143540 421248 143546
rect 421196 143482 421248 143488
rect 421196 133952 421248 133958
rect 421196 133894 421248 133900
rect 421208 124166 421236 133894
rect 421196 124160 421248 124166
rect 421196 124102 421248 124108
rect 421196 114572 421248 114578
rect 421196 114514 421248 114520
rect 421208 104854 421236 114514
rect 421196 104848 421248 104854
rect 421196 104790 421248 104796
rect 421196 87032 421248 87038
rect 421196 86974 421248 86980
rect 421208 85542 421236 86974
rect 421196 85536 421248 85542
rect 421196 85478 421248 85484
rect 421012 75948 421064 75954
rect 421012 75890 421064 75896
rect 421024 67697 421052 75890
rect 421010 67688 421066 67697
rect 421010 67623 421066 67632
rect 421194 67688 421250 67697
rect 421194 67623 421250 67632
rect 421208 66230 421236 67623
rect 421196 66224 421248 66230
rect 421196 66166 421248 66172
rect 421104 56704 421156 56710
rect 421104 56646 421156 56652
rect 421116 56574 421144 56646
rect 421104 56568 421156 56574
rect 421104 56510 421156 56516
rect 421012 46980 421064 46986
rect 421012 46922 421064 46928
rect 421024 42090 421052 46922
rect 421012 42084 421064 42090
rect 421012 42026 421064 42032
rect 421012 27668 421064 27674
rect 421012 27610 421064 27616
rect 421024 22778 421052 27610
rect 421012 22772 421064 22778
rect 421012 22714 421064 22720
rect 421472 9716 421524 9722
rect 421472 9658 421524 9664
rect 421484 9602 421512 9658
rect 421392 9574 421512 9602
rect 420828 3528 420880 3534
rect 421392 3505 421420 9574
rect 421576 3670 421604 337078
rect 422496 336802 422524 340068
rect 422208 336796 422260 336802
rect 422208 336738 422260 336744
rect 422484 336796 422536 336802
rect 422484 336738 422536 336744
rect 422220 4894 422248 336738
rect 423416 335594 423444 340190
rect 423508 337278 423536 340068
rect 423496 337272 423548 337278
rect 423496 337214 423548 337220
rect 423968 337210 423996 340068
rect 423956 337204 424008 337210
rect 423956 337146 424008 337152
rect 424428 336802 424456 340068
rect 424692 337612 424744 337618
rect 424692 337554 424744 337560
rect 424324 336796 424376 336802
rect 424324 336738 424376 336744
rect 424416 336796 424468 336802
rect 424416 336738 424468 336744
rect 423416 335566 423628 335594
rect 423496 110628 423548 110634
rect 423496 110570 423548 110576
rect 423508 110537 423536 110570
rect 423494 110528 423550 110537
rect 423494 110463 423550 110472
rect 422208 4888 422260 4894
rect 422208 4830 422260 4836
rect 423600 4826 423628 335566
rect 424140 311908 424192 311914
rect 424140 311850 424192 311856
rect 424152 302258 424180 311850
rect 424140 302252 424192 302258
rect 424140 302194 424192 302200
rect 424048 183592 424100 183598
rect 424048 183534 424100 183540
rect 424060 183462 424088 183534
rect 424048 183456 424100 183462
rect 424048 183398 424100 183404
rect 424232 176588 424284 176594
rect 424232 176530 424284 176536
rect 424244 167006 424272 176530
rect 424232 167000 424284 167006
rect 424232 166942 424284 166948
rect 424140 142860 424192 142866
rect 424140 142802 424192 142808
rect 424152 128382 424180 142802
rect 424140 128376 424192 128382
rect 424140 128318 424192 128324
rect 423588 4820 423640 4826
rect 423588 4762 423640 4768
rect 423956 4004 424008 4010
rect 423956 3946 424008 3952
rect 421564 3664 421616 3670
rect 421564 3606 421616 3612
rect 420828 3470 420880 3476
rect 421378 3496 421434 3505
rect 421378 3431 421434 3440
rect 421562 3496 421618 3505
rect 421562 3431 421618 3440
rect 422760 3460 422812 3466
rect 420184 3324 420236 3330
rect 420184 3266 420236 3272
rect 420368 3052 420420 3058
rect 420368 2994 420420 3000
rect 420380 480 420408 2994
rect 421576 480 421604 3431
rect 422760 3402 422812 3408
rect 422772 480 422800 3402
rect 423968 480 423996 3946
rect 424336 3466 424364 336738
rect 424704 318850 424732 337554
rect 424980 336870 425008 340068
rect 425440 337754 425468 340068
rect 425914 340054 426388 340082
rect 425428 337748 425480 337754
rect 425428 337690 425480 337696
rect 424968 336864 425020 336870
rect 424968 336806 425020 336812
rect 424968 336728 425020 336734
rect 424968 336670 425020 336676
rect 424600 318844 424652 318850
rect 424600 318786 424652 318792
rect 424692 318844 424744 318850
rect 424692 318786 424744 318792
rect 424612 311914 424640 318786
rect 424600 311908 424652 311914
rect 424600 311850 424652 311856
rect 424508 302252 424560 302258
rect 424508 302194 424560 302200
rect 424520 302138 424548 302194
rect 424520 302110 424640 302138
rect 424612 292618 424640 302110
rect 424612 292590 424732 292618
rect 424704 282946 424732 292590
rect 424508 282940 424560 282946
rect 424508 282882 424560 282888
rect 424692 282940 424744 282946
rect 424692 282882 424744 282888
rect 424520 282826 424548 282882
rect 424520 282798 424640 282826
rect 424612 280158 424640 282798
rect 424600 280152 424652 280158
rect 424600 280094 424652 280100
rect 424784 270564 424836 270570
rect 424784 270506 424836 270512
rect 424796 263514 424824 270506
rect 424612 263486 424824 263514
rect 424612 260846 424640 263486
rect 424600 260840 424652 260846
rect 424600 260782 424652 260788
rect 424508 251252 424560 251258
rect 424508 251194 424560 251200
rect 424520 224890 424548 251194
rect 424520 224862 424640 224890
rect 424612 215370 424640 224862
rect 424612 215342 424824 215370
rect 424796 212537 424824 215342
rect 424598 212528 424654 212537
rect 424598 212463 424654 212472
rect 424782 212528 424838 212537
rect 424782 212463 424838 212472
rect 424612 202910 424640 212463
rect 424600 202904 424652 202910
rect 424600 202846 424652 202852
rect 424876 202904 424928 202910
rect 424876 202846 424928 202852
rect 424888 196042 424916 202846
rect 424692 196036 424744 196042
rect 424692 195978 424744 195984
rect 424876 196036 424928 196042
rect 424876 195978 424928 195984
rect 424704 183598 424732 195978
rect 424692 183592 424744 183598
rect 424692 183534 424744 183540
rect 424416 166932 424468 166938
rect 424416 166874 424468 166880
rect 424428 164218 424456 166874
rect 424416 164212 424468 164218
rect 424416 164154 424468 164160
rect 424508 164212 424560 164218
rect 424508 164154 424560 164160
rect 424520 154578 424548 164154
rect 424520 154550 424640 154578
rect 424612 142866 424640 154550
rect 424600 142860 424652 142866
rect 424600 142802 424652 142808
rect 424508 128376 424560 128382
rect 424560 128324 424732 128330
rect 424508 128318 424732 128324
rect 424520 128302 424732 128318
rect 424704 115938 424732 128302
rect 424600 115932 424652 115938
rect 424600 115874 424652 115880
rect 424692 115932 424744 115938
rect 424692 115874 424744 115880
rect 424612 114510 424640 115874
rect 424600 114504 424652 114510
rect 424600 114446 424652 114452
rect 424508 104916 424560 104922
rect 424508 104858 424560 104864
rect 424520 99414 424548 104858
rect 424508 99408 424560 99414
rect 424508 99350 424560 99356
rect 424692 99340 424744 99346
rect 424692 99282 424744 99288
rect 424704 89758 424732 99282
rect 424508 89752 424560 89758
rect 424508 89694 424560 89700
rect 424692 89752 424744 89758
rect 424692 89694 424744 89700
rect 424520 72570 424548 89694
rect 424520 72542 424640 72570
rect 424612 72298 424640 72542
rect 424520 72270 424640 72298
rect 424520 70258 424548 72270
rect 424520 70230 424732 70258
rect 424704 60738 424732 70230
rect 424520 60710 424732 60738
rect 424520 53854 424548 60710
rect 424508 53848 424560 53854
rect 424508 53790 424560 53796
rect 424692 48340 424744 48346
rect 424692 48282 424744 48288
rect 424704 48226 424732 48282
rect 424612 48198 424732 48226
rect 424612 38706 424640 48198
rect 424520 38678 424640 38706
rect 424520 38622 424548 38678
rect 424508 38616 424560 38622
rect 424508 38558 424560 38564
rect 424600 29028 424652 29034
rect 424600 28970 424652 28976
rect 424612 22166 424640 28970
rect 424600 22160 424652 22166
rect 424600 22102 424652 22108
rect 424508 22092 424560 22098
rect 424508 22034 424560 22040
rect 424520 12458 424548 22034
rect 424520 12430 424640 12458
rect 424612 4010 424640 12430
rect 424980 4214 425008 336670
rect 426360 5778 426388 340054
rect 426452 337618 426480 340068
rect 426440 337612 426492 337618
rect 426440 337554 426492 337560
rect 426440 337408 426492 337414
rect 426440 337350 426492 337356
rect 426452 12442 426480 337350
rect 426912 337074 426940 340068
rect 427386 340054 427768 340082
rect 427084 337680 427136 337686
rect 427084 337622 427136 337628
rect 426900 337068 426952 337074
rect 426900 337010 426952 337016
rect 426440 12436 426492 12442
rect 426440 12378 426492 12384
rect 426348 5772 426400 5778
rect 426348 5714 426400 5720
rect 424968 4208 425020 4214
rect 424968 4150 425020 4156
rect 424600 4004 424652 4010
rect 424600 3946 424652 3952
rect 425152 4004 425204 4010
rect 425152 3946 425204 3952
rect 424324 3460 424376 3466
rect 424324 3402 424376 3408
rect 425164 480 425192 3946
rect 427096 3670 427124 337622
rect 427544 12436 427596 12442
rect 427544 12378 427596 12384
rect 427084 3664 427136 3670
rect 427084 3606 427136 3612
rect 426348 3120 426400 3126
rect 426348 3062 426400 3068
rect 426360 480 426388 3062
rect 427556 480 427584 12378
rect 427740 5846 427768 340054
rect 427924 337550 427952 340068
rect 428384 337618 428412 340068
rect 428858 340054 429148 340082
rect 428464 337748 428516 337754
rect 428464 337690 428516 337696
rect 428372 337612 428424 337618
rect 428372 337554 428424 337560
rect 427912 337544 427964 337550
rect 427912 337486 427964 337492
rect 427728 5840 427780 5846
rect 427728 5782 427780 5788
rect 428476 3126 428504 337690
rect 429120 5982 429148 340054
rect 429396 337754 429424 340068
rect 429752 338020 429804 338026
rect 429752 337962 429804 337968
rect 429384 337748 429436 337754
rect 429384 337690 429436 337696
rect 429764 337226 429792 337962
rect 429856 337414 429884 340068
rect 430330 340054 430436 340082
rect 429844 337408 429896 337414
rect 429844 337350 429896 337356
rect 429764 337198 429884 337226
rect 429108 5976 429160 5982
rect 429108 5918 429160 5924
rect 428464 3120 428516 3126
rect 428464 3062 428516 3068
rect 429856 2990 429884 337198
rect 430408 6118 430436 340054
rect 430488 337748 430540 337754
rect 430488 337690 430540 337696
rect 430396 6112 430448 6118
rect 430396 6054 430448 6060
rect 430500 5914 430528 337690
rect 430868 337686 430896 340068
rect 430856 337680 430908 337686
rect 430856 337622 430908 337628
rect 431328 337618 431356 340068
rect 431408 338088 431460 338094
rect 431408 338030 431460 338036
rect 431224 337612 431276 337618
rect 431224 337554 431276 337560
rect 431316 337612 431368 337618
rect 431316 337554 431368 337560
rect 430488 5908 430540 5914
rect 430488 5850 430540 5856
rect 431132 3664 431184 3670
rect 431132 3606 431184 3612
rect 429936 3188 429988 3194
rect 429936 3130 429988 3136
rect 428740 2984 428792 2990
rect 428740 2926 428792 2932
rect 429844 2984 429896 2990
rect 429844 2926 429896 2932
rect 428752 480 428780 2926
rect 429948 480 429976 3130
rect 431144 480 431172 3606
rect 431236 3194 431264 337554
rect 431420 337498 431448 338030
rect 431328 337470 431448 337498
rect 431224 3188 431276 3194
rect 431224 3130 431276 3136
rect 431328 3058 431356 337470
rect 431788 6798 431816 340068
rect 432340 337754 432368 340068
rect 432328 337748 432380 337754
rect 432328 337690 432380 337696
rect 431868 337680 431920 337686
rect 431868 337622 431920 337628
rect 431776 6792 431828 6798
rect 431776 6734 431828 6740
rect 431880 6050 431908 337622
rect 432800 337210 432828 340068
rect 433168 340054 433274 340082
rect 432788 337204 432840 337210
rect 432788 337146 432840 337152
rect 433168 6662 433196 340054
rect 433720 337754 433748 340068
rect 433248 337748 433300 337754
rect 433248 337690 433300 337696
rect 433708 337748 433760 337754
rect 433708 337690 433760 337696
rect 433260 6866 433288 337690
rect 434272 337482 434300 340068
rect 434628 337748 434680 337754
rect 434628 337690 434680 337696
rect 433984 337476 434036 337482
rect 433984 337418 434036 337424
rect 434260 337476 434312 337482
rect 434260 337418 434312 337424
rect 433524 337136 433576 337142
rect 433524 337078 433576 337084
rect 433248 6860 433300 6866
rect 433248 6802 433300 6808
rect 433156 6656 433208 6662
rect 433156 6598 433208 6604
rect 431868 6044 431920 6050
rect 431868 5986 431920 5992
rect 433536 5522 433564 337078
rect 433536 5494 433840 5522
rect 433524 5432 433576 5438
rect 433524 5374 433576 5380
rect 432328 3256 432380 3262
rect 432328 3198 432380 3204
rect 431316 3052 431368 3058
rect 431316 2994 431368 3000
rect 432340 480 432368 3198
rect 433536 480 433564 5374
rect 433812 3074 433840 5494
rect 433996 3398 434024 337418
rect 434640 6730 434668 337690
rect 434732 337686 434760 340068
rect 435192 337754 435220 340068
rect 435744 338094 435772 340068
rect 435732 338088 435784 338094
rect 435732 338030 435784 338036
rect 435180 337748 435232 337754
rect 435180 337690 435232 337696
rect 436008 337748 436060 337754
rect 436008 337690 436060 337696
rect 434720 337680 434772 337686
rect 434720 337622 434772 337628
rect 435916 337680 435968 337686
rect 435916 337622 435968 337628
rect 434628 6724 434680 6730
rect 434628 6666 434680 6672
rect 435928 6594 435956 337622
rect 435916 6588 435968 6594
rect 435916 6530 435968 6536
rect 436020 6526 436048 337690
rect 436204 337686 436232 340068
rect 436664 337754 436692 340068
rect 437216 338026 437244 340068
rect 437204 338020 437256 338026
rect 437204 337962 437256 337968
rect 437676 337754 437704 340068
rect 438124 337816 438176 337822
rect 438124 337758 438176 337764
rect 436652 337748 436704 337754
rect 436652 337690 436704 337696
rect 437388 337748 437440 337754
rect 437388 337690 437440 337696
rect 437664 337748 437716 337754
rect 437664 337690 437716 337696
rect 436192 337680 436244 337686
rect 436192 337622 436244 337628
rect 437296 337680 437348 337686
rect 437296 337622 437348 337628
rect 437202 157584 437258 157593
rect 437202 157519 437204 157528
rect 437256 157519 437258 157528
rect 437204 157490 437256 157496
rect 437202 110664 437258 110673
rect 437202 110599 437204 110608
rect 437256 110599 437258 110608
rect 437204 110570 437256 110576
rect 437204 87168 437256 87174
rect 437202 87136 437204 87145
rect 437256 87136 437258 87145
rect 437202 87071 437258 87080
rect 437202 76120 437258 76129
rect 437202 76055 437204 76064
rect 437256 76055 437258 76064
rect 437204 76026 437256 76032
rect 437202 63744 437258 63753
rect 437202 63679 437204 63688
rect 437256 63679 437258 63688
rect 437204 63650 437256 63656
rect 437204 40248 437256 40254
rect 437202 40216 437204 40225
rect 437256 40216 437258 40225
rect 437202 40151 437258 40160
rect 437202 29200 437258 29209
rect 437202 29135 437204 29144
rect 437256 29135 437258 29144
rect 437204 29106 437256 29112
rect 437202 16824 437258 16833
rect 437202 16759 437204 16768
rect 437256 16759 437258 16768
rect 437204 16730 437256 16736
rect 436008 6520 436060 6526
rect 436008 6462 436060 6468
rect 437308 6458 437336 337622
rect 437296 6452 437348 6458
rect 437296 6394 437348 6400
rect 437400 6390 437428 337690
rect 437478 157584 437534 157593
rect 437478 157519 437480 157528
rect 437532 157519 437534 157528
rect 437480 157490 437532 157496
rect 437478 110664 437534 110673
rect 437478 110599 437480 110608
rect 437532 110599 437534 110608
rect 437480 110570 437532 110576
rect 437480 87168 437532 87174
rect 437478 87136 437480 87145
rect 437532 87136 437534 87145
rect 437478 87071 437534 87080
rect 437478 76120 437534 76129
rect 437478 76055 437480 76064
rect 437532 76055 437534 76064
rect 437480 76026 437532 76032
rect 437478 63744 437534 63753
rect 437478 63679 437480 63688
rect 437532 63679 437534 63688
rect 437480 63650 437532 63656
rect 437480 40248 437532 40254
rect 437478 40216 437480 40225
rect 437532 40216 437534 40225
rect 437478 40151 437534 40160
rect 437478 29200 437534 29209
rect 437478 29135 437480 29144
rect 437532 29135 437534 29144
rect 437480 29106 437532 29112
rect 437478 16824 437534 16833
rect 437478 16759 437480 16768
rect 437532 16759 437534 16768
rect 437480 16730 437532 16736
rect 437388 6384 437440 6390
rect 437388 6326 437440 6332
rect 438136 3398 438164 337758
rect 438596 337668 438624 340190
rect 438688 337822 438716 340068
rect 438676 337816 438728 337822
rect 438676 337758 438728 337764
rect 439148 337754 439176 340068
rect 439622 340054 440096 340082
rect 438768 337748 438820 337754
rect 438768 337690 438820 337696
rect 439136 337748 439188 337754
rect 439136 337690 439188 337696
rect 438596 337640 438716 337668
rect 438688 6254 438716 337640
rect 438780 6322 438808 337690
rect 439596 337476 439648 337482
rect 439596 337418 439648 337424
rect 439504 336864 439556 336870
rect 439504 336806 439556 336812
rect 438768 6316 438820 6322
rect 438768 6258 438820 6264
rect 438676 6248 438728 6254
rect 438676 6190 438728 6196
rect 438216 4140 438268 4146
rect 438216 4082 438268 4088
rect 433984 3392 434036 3398
rect 433984 3334 434036 3340
rect 435824 3392 435876 3398
rect 435824 3334 435876 3340
rect 438124 3392 438176 3398
rect 438124 3334 438176 3340
rect 433812 3046 434668 3074
rect 434640 480 434668 3046
rect 435836 480 435864 3334
rect 437020 3256 437072 3262
rect 437020 3198 437072 3204
rect 437032 480 437060 3198
rect 438228 480 438256 4082
rect 439412 4072 439464 4078
rect 439412 4014 439464 4020
rect 439424 480 439452 4014
rect 439516 2854 439544 336806
rect 439608 4078 439636 337418
rect 440068 7342 440096 340054
rect 440160 337906 440188 340068
rect 440160 337878 440280 337906
rect 440148 337748 440200 337754
rect 440148 337690 440200 337696
rect 440056 7336 440108 7342
rect 440056 7278 440108 7284
rect 440160 6186 440188 337690
rect 440252 337550 440280 337878
rect 440620 337822 440648 340068
rect 441094 340054 441476 340082
rect 440608 337816 440660 337822
rect 440608 337758 440660 337764
rect 440240 337544 440292 337550
rect 440240 337486 440292 337492
rect 441448 7410 441476 340054
rect 441632 337822 441660 340068
rect 441528 337816 441580 337822
rect 441528 337758 441580 337764
rect 441620 337816 441672 337822
rect 441620 337758 441672 337764
rect 441436 7404 441488 7410
rect 441436 7346 441488 7352
rect 440148 6180 440200 6186
rect 440148 6122 440200 6128
rect 440608 5364 440660 5370
rect 440608 5306 440660 5312
rect 439596 4072 439648 4078
rect 439596 4014 439648 4020
rect 439504 2848 439556 2854
rect 439504 2790 439556 2796
rect 440620 480 440648 5306
rect 441540 4282 441568 337758
rect 442092 337686 442120 340068
rect 442566 340054 442856 340082
rect 442356 338020 442408 338026
rect 442356 337962 442408 337968
rect 442080 337680 442132 337686
rect 442080 337622 442132 337628
rect 442264 337612 442316 337618
rect 442264 337554 442316 337560
rect 441528 4276 441580 4282
rect 441528 4218 441580 4224
rect 442276 4146 442304 337554
rect 442264 4140 442316 4146
rect 442264 4082 442316 4088
rect 441620 3936 441672 3942
rect 441672 3884 441844 3890
rect 441620 3878 441844 3884
rect 441632 3862 441844 3878
rect 441816 480 441844 3862
rect 442368 3670 442396 337962
rect 442828 7478 442856 340054
rect 442908 337680 442960 337686
rect 442908 337622 442960 337628
rect 442816 7472 442868 7478
rect 442816 7414 442868 7420
rect 442920 4350 442948 337622
rect 443104 337482 443132 340068
rect 443564 337686 443592 340068
rect 444038 340054 444236 340082
rect 443644 337816 443696 337822
rect 443644 337758 443696 337764
rect 443552 337680 443604 337686
rect 443552 337622 443604 337628
rect 443092 337476 443144 337482
rect 443092 337418 443144 337424
rect 442908 4344 442960 4350
rect 442908 4286 442960 4292
rect 443000 3800 443052 3806
rect 443000 3742 443052 3748
rect 442356 3664 442408 3670
rect 442356 3606 442408 3612
rect 443012 480 443040 3742
rect 443656 3670 443684 337758
rect 444208 7546 444236 340054
rect 444576 337822 444604 340068
rect 444564 337816 444616 337822
rect 444564 337758 444616 337764
rect 445036 337686 445064 340068
rect 444288 337680 444340 337686
rect 444288 337622 444340 337628
rect 445024 337680 445076 337686
rect 445024 337622 445076 337628
rect 444196 7540 444248 7546
rect 444196 7482 444248 7488
rect 444196 5296 444248 5302
rect 444196 5238 444248 5244
rect 443644 3664 443696 3670
rect 443644 3606 443696 3612
rect 444208 480 444236 5238
rect 444300 4418 444328 337622
rect 445496 8294 445524 340068
rect 446048 338026 446076 340068
rect 446036 338020 446088 338026
rect 446036 337962 446088 337968
rect 445668 337816 445720 337822
rect 445668 337758 445720 337764
rect 445576 337680 445628 337686
rect 445576 337622 445628 337628
rect 445484 8288 445536 8294
rect 445484 8230 445536 8236
rect 445588 4486 445616 337622
rect 445576 4480 445628 4486
rect 445576 4422 445628 4428
rect 444288 4412 444340 4418
rect 444288 4354 444340 4360
rect 445680 4146 445708 337758
rect 446508 337686 446536 340068
rect 446496 337680 446548 337686
rect 446496 337622 446548 337628
rect 446968 8226 446996 340068
rect 447048 337680 447100 337686
rect 447048 337622 447100 337628
rect 446956 8220 447008 8226
rect 446956 8162 447008 8168
rect 447060 4554 447088 337622
rect 447520 337550 447548 340068
rect 447994 340054 448376 340082
rect 448244 337680 448296 337686
rect 448244 337622 448296 337628
rect 447508 337544 447560 337550
rect 447508 337486 447560 337492
rect 448256 8158 448284 337622
rect 448244 8152 448296 8158
rect 448244 8094 448296 8100
rect 447784 5228 447836 5234
rect 447784 5170 447836 5176
rect 447048 4548 447100 4554
rect 447048 4490 447100 4496
rect 445668 4140 445720 4146
rect 445668 4082 445720 4088
rect 445392 3868 445444 3874
rect 445392 3810 445444 3816
rect 445404 480 445432 3810
rect 446588 3664 446640 3670
rect 446232 3612 446588 3618
rect 446232 3606 446640 3612
rect 446232 3590 446628 3606
rect 446232 3262 446260 3590
rect 446588 3324 446640 3330
rect 446588 3266 446640 3272
rect 446220 3256 446272 3262
rect 446220 3198 446272 3204
rect 446600 480 446628 3266
rect 447796 480 447824 5170
rect 448348 4622 448376 340054
rect 448440 337686 448468 340068
rect 448992 337822 449020 340068
rect 449466 340054 449848 340082
rect 448980 337816 449032 337822
rect 448980 337758 449032 337764
rect 448428 337680 448480 337686
rect 448428 337622 448480 337628
rect 449164 337612 449216 337618
rect 449164 337554 449216 337560
rect 448428 337544 448480 337550
rect 448428 337486 448480 337492
rect 448336 4616 448388 4622
rect 448336 4558 448388 4564
rect 448440 4078 448468 337486
rect 448428 4072 448480 4078
rect 448428 4014 448480 4020
rect 449176 3670 449204 337554
rect 449820 4690 449848 340054
rect 449912 337686 449940 340068
rect 449900 337680 449952 337686
rect 449900 337622 449952 337628
rect 450464 337618 450492 340068
rect 450938 340054 451136 340082
rect 451004 337680 451056 337686
rect 451004 337622 451056 337628
rect 450452 337612 450504 337618
rect 450452 337554 450504 337560
rect 451016 8090 451044 337622
rect 451004 8084 451056 8090
rect 451004 8026 451056 8032
rect 451108 4758 451136 340054
rect 451384 337618 451412 340068
rect 451188 337612 451240 337618
rect 451188 337554 451240 337560
rect 451372 337612 451424 337618
rect 451372 337554 451424 337560
rect 451096 4752 451148 4758
rect 451096 4694 451148 4700
rect 449808 4684 449860 4690
rect 449808 4626 449860 4632
rect 451200 4010 451228 337554
rect 451844 336870 451872 340068
rect 452410 340054 452608 340082
rect 452476 337612 452528 337618
rect 452476 337554 452528 337560
rect 451832 336864 451884 336870
rect 451832 336806 451884 336812
rect 452488 8022 452516 337554
rect 452476 8016 452528 8022
rect 452476 7958 452528 7964
rect 452580 5506 452608 340054
rect 452856 337822 452884 340068
rect 452844 337816 452896 337822
rect 452844 337758 452896 337764
rect 453316 337618 453344 340068
rect 453764 337816 453816 337822
rect 453764 337758 453816 337764
rect 453304 337612 453356 337618
rect 453304 337554 453356 337560
rect 453776 7954 453804 337758
rect 453764 7948 453816 7954
rect 453764 7890 453816 7896
rect 452568 5500 452620 5506
rect 452568 5442 452620 5448
rect 453868 5438 453896 340068
rect 454328 337822 454356 340068
rect 454788 338026 454816 340068
rect 454776 338020 454828 338026
rect 454776 337962 454828 337968
rect 454316 337816 454368 337822
rect 454316 337758 454368 337764
rect 455236 337816 455288 337822
rect 455236 337758 455288 337764
rect 453948 337612 454000 337618
rect 453948 337554 454000 337560
rect 453856 5432 453908 5438
rect 453856 5374 453908 5380
rect 451280 5160 451332 5166
rect 451280 5102 451332 5108
rect 450176 4004 450228 4010
rect 450176 3946 450228 3952
rect 451188 4004 451240 4010
rect 451188 3946 451240 3952
rect 449164 3664 449216 3670
rect 449164 3606 449216 3612
rect 448980 2984 449032 2990
rect 448980 2926 449032 2932
rect 448992 480 449020 2926
rect 450188 480 450216 3946
rect 451292 480 451320 5102
rect 453960 3942 453988 337554
rect 455248 7886 455276 337758
rect 455236 7880 455288 7886
rect 455236 7822 455288 7828
rect 455340 5370 455368 340068
rect 455604 337952 455656 337958
rect 455604 337894 455656 337900
rect 455328 5364 455380 5370
rect 455328 5306 455380 5312
rect 454868 5092 454920 5098
rect 454868 5034 454920 5040
rect 453672 3936 453724 3942
rect 453672 3878 453724 3884
rect 453948 3936 454000 3942
rect 453948 3878 454000 3884
rect 452476 3800 452528 3806
rect 452476 3742 452528 3748
rect 452488 480 452516 3742
rect 453684 480 453712 3878
rect 454880 480 454908 5034
rect 455616 1442 455644 337894
rect 455800 337822 455828 340068
rect 456274 340054 456748 340082
rect 455788 337816 455840 337822
rect 455788 337758 455840 337764
rect 456616 337816 456668 337822
rect 456616 337758 456668 337764
rect 456522 157584 456578 157593
rect 456522 157519 456524 157528
rect 456576 157519 456578 157528
rect 456524 157490 456576 157496
rect 456524 110696 456576 110702
rect 456522 110664 456524 110673
rect 456576 110664 456578 110673
rect 456522 110599 456578 110608
rect 456524 87168 456576 87174
rect 456522 87136 456524 87145
rect 456576 87136 456578 87145
rect 456522 87071 456578 87080
rect 456522 76120 456578 76129
rect 456522 76055 456524 76064
rect 456576 76055 456578 76064
rect 456524 76026 456576 76032
rect 456522 63744 456578 63753
rect 456522 63679 456524 63688
rect 456576 63679 456578 63688
rect 456524 63650 456576 63656
rect 456522 40216 456578 40225
rect 456522 40151 456524 40160
rect 456576 40151 456578 40160
rect 456524 40122 456576 40128
rect 456524 29232 456576 29238
rect 456522 29200 456524 29209
rect 456576 29200 456578 29209
rect 456522 29135 456578 29144
rect 456524 16856 456576 16862
rect 456522 16824 456524 16833
rect 456576 16824 456578 16833
rect 456522 16759 456578 16768
rect 456628 7818 456656 337758
rect 456616 7812 456668 7818
rect 456616 7754 456668 7760
rect 456720 3806 456748 340054
rect 456812 337550 456840 340068
rect 456800 337544 456852 337550
rect 456800 337486 456852 337492
rect 457272 336802 457300 340068
rect 457732 337822 457760 340068
rect 457720 337816 457772 337822
rect 457720 337758 457772 337764
rect 458088 337544 458140 337550
rect 458088 337486 458140 337492
rect 457260 336796 457312 336802
rect 457260 336738 457312 336744
rect 457996 336796 458048 336802
rect 457996 336738 458048 336744
rect 456890 157584 456946 157593
rect 456890 157519 456892 157528
rect 456944 157519 456946 157528
rect 456892 157490 456944 157496
rect 456984 87168 457036 87174
rect 456982 87136 456984 87145
rect 457036 87136 457038 87145
rect 456982 87071 457038 87080
rect 456798 76120 456854 76129
rect 456798 76055 456800 76064
rect 456852 76055 456854 76064
rect 456800 76026 456852 76032
rect 456890 63744 456946 63753
rect 456890 63679 456892 63688
rect 456944 63679 456946 63688
rect 456892 63650 456944 63656
rect 456890 40216 456946 40225
rect 456890 40151 456892 40160
rect 456944 40151 456946 40160
rect 456892 40122 456944 40128
rect 456984 29232 457036 29238
rect 456982 29200 456984 29209
rect 457036 29200 457038 29209
rect 456982 29135 457038 29144
rect 458008 7750 458036 336738
rect 457996 7744 458048 7750
rect 457996 7686 458048 7692
rect 458100 5098 458128 337486
rect 458284 336802 458312 340068
rect 458744 337958 458772 340068
rect 458732 337952 458784 337958
rect 458732 337894 458784 337900
rect 459204 336870 459232 340068
rect 459376 337952 459428 337958
rect 459376 337894 459428 337900
rect 459192 336864 459244 336870
rect 459192 336806 459244 336812
rect 458272 336796 458324 336802
rect 458272 336738 458324 336744
rect 458824 110696 458876 110702
rect 458822 110664 458824 110673
rect 458876 110664 458878 110673
rect 458822 110599 458878 110608
rect 458824 16856 458876 16862
rect 458822 16824 458824 16833
rect 458876 16824 458878 16833
rect 458822 16759 458878 16768
rect 459388 7682 459416 337894
rect 459756 336802 459784 340068
rect 460230 340054 460428 340082
rect 460690 340054 460888 340082
rect 460296 337272 460348 337278
rect 460296 337214 460348 337220
rect 460204 336864 460256 336870
rect 460204 336806 460256 336812
rect 459468 336796 459520 336802
rect 459468 336738 459520 336744
rect 459744 336796 459796 336802
rect 459744 336738 459796 336744
rect 459376 7676 459428 7682
rect 459376 7618 459428 7624
rect 459480 5302 459508 336738
rect 459468 5296 459520 5302
rect 459468 5238 459520 5244
rect 458088 5092 458140 5098
rect 458088 5034 458140 5040
rect 458456 5024 458508 5030
rect 458456 4966 458508 4972
rect 456708 3800 456760 3806
rect 456708 3742 456760 3748
rect 457260 3596 457312 3602
rect 457260 3538 457312 3544
rect 455616 1414 456104 1442
rect 456076 480 456104 1414
rect 457272 480 457300 3538
rect 458468 480 458496 4966
rect 460112 3800 460164 3806
rect 460110 3768 460112 3777
rect 460164 3768 460166 3777
rect 460216 3738 460244 336806
rect 460308 3806 460336 337214
rect 460400 336870 460428 340054
rect 460860 338162 460888 340054
rect 460848 338156 460900 338162
rect 460848 338098 460900 338104
rect 460388 336864 460440 336870
rect 460388 336806 460440 336812
rect 460756 336864 460808 336870
rect 460756 336806 460808 336812
rect 460768 7614 460796 336806
rect 461228 336802 461256 340068
rect 461688 338026 461716 340068
rect 462162 340054 462268 340082
rect 461676 338020 461728 338026
rect 461676 337962 461728 337968
rect 460848 336796 460900 336802
rect 460848 336738 460900 336744
rect 461216 336796 461268 336802
rect 461216 336738 461268 336744
rect 462136 336796 462188 336802
rect 462136 336738 462188 336744
rect 460756 7608 460808 7614
rect 460756 7550 460808 7556
rect 460860 5234 460888 336738
rect 460848 5228 460900 5234
rect 460848 5170 460900 5176
rect 462044 5024 462096 5030
rect 462044 4966 462096 4972
rect 460296 3800 460348 3806
rect 460296 3742 460348 3748
rect 460110 3703 460166 3712
rect 460204 3732 460256 3738
rect 460204 3674 460256 3680
rect 460848 3528 460900 3534
rect 460848 3470 460900 3476
rect 459652 3052 459704 3058
rect 459652 2994 459704 3000
rect 459664 480 459692 2994
rect 460860 480 460888 3470
rect 462056 480 462084 4966
rect 462148 4826 462176 336738
rect 462136 4820 462188 4826
rect 462136 4762 462188 4768
rect 462240 3602 462268 340054
rect 462700 336802 462728 340068
rect 463174 340054 463464 340082
rect 463436 336920 463464 340054
rect 463620 337278 463648 340068
rect 463884 337340 463936 337346
rect 463884 337282 463936 337288
rect 463608 337272 463660 337278
rect 463608 337214 463660 337220
rect 463436 336892 463648 336920
rect 462688 336796 462740 336802
rect 462688 336738 462740 336744
rect 463516 336796 463568 336802
rect 463516 336738 463568 336744
rect 463528 5166 463556 336738
rect 463516 5160 463568 5166
rect 463516 5102 463568 5108
rect 463240 3800 463292 3806
rect 463240 3742 463292 3748
rect 463514 3768 463570 3777
rect 462228 3596 462280 3602
rect 462228 3538 462280 3544
rect 463252 480 463280 3742
rect 463514 3703 463570 3712
rect 463528 3602 463556 3703
rect 463620 3670 463648 336892
rect 463896 325718 463924 337282
rect 464172 336802 464200 340068
rect 464646 340054 464936 340082
rect 464908 336920 464936 340054
rect 465092 337346 465120 340068
rect 465658 340054 465948 340082
rect 466118 340054 466316 340082
rect 465080 337340 465132 337346
rect 465080 337282 465132 337288
rect 464908 336892 465120 336920
rect 465092 336802 465120 336892
rect 464160 336796 464212 336802
rect 464160 336738 464212 336744
rect 464988 336796 465040 336802
rect 464988 336738 465040 336744
rect 465080 336796 465132 336802
rect 465080 336738 465132 336744
rect 463700 325712 463752 325718
rect 463700 325654 463752 325660
rect 463884 325712 463936 325718
rect 463884 325654 463936 325660
rect 463712 316010 463740 325654
rect 463712 315982 463924 316010
rect 463896 306406 463924 315982
rect 463700 306400 463752 306406
rect 463700 306342 463752 306348
rect 463884 306400 463936 306406
rect 463884 306342 463936 306348
rect 463712 296698 463740 306342
rect 463712 296670 463924 296698
rect 463896 287094 463924 296670
rect 463700 287088 463752 287094
rect 463700 287030 463752 287036
rect 463884 287088 463936 287094
rect 463884 287030 463936 287036
rect 463712 277386 463740 287030
rect 463712 277358 463924 277386
rect 463896 267782 463924 277358
rect 463700 267776 463752 267782
rect 463884 267776 463936 267782
rect 463752 267724 463832 267730
rect 463700 267718 463832 267724
rect 463884 267718 463936 267724
rect 463712 267702 463832 267718
rect 463804 267594 463832 267702
rect 463804 267566 463924 267594
rect 463896 263514 463924 267566
rect 463804 263486 463924 263514
rect 463804 260846 463832 263486
rect 463792 260840 463844 260846
rect 463792 260782 463844 260788
rect 463700 251252 463752 251258
rect 463700 251194 463752 251200
rect 463712 244202 463740 251194
rect 463712 244174 463832 244202
rect 463804 234682 463832 244174
rect 463804 234654 464016 234682
rect 463988 231849 464016 234654
rect 463790 231840 463846 231849
rect 463790 231775 463846 231784
rect 463974 231840 464030 231849
rect 463974 231775 464030 231784
rect 463804 222222 463832 231775
rect 463792 222216 463844 222222
rect 463792 222158 463844 222164
rect 464068 222216 464120 222222
rect 464068 222158 464120 222164
rect 464080 215422 464108 222158
rect 464068 215416 464120 215422
rect 464068 215358 464120 215364
rect 463976 215280 464028 215286
rect 463976 215222 464028 215228
rect 463988 212537 464016 215222
rect 463790 212528 463846 212537
rect 463790 212463 463846 212472
rect 463974 212528 464030 212537
rect 463974 212463 464030 212472
rect 463804 202910 463832 212463
rect 463792 202904 463844 202910
rect 463792 202846 463844 202852
rect 464068 202904 464120 202910
rect 464068 202846 464120 202852
rect 464080 196110 464108 202846
rect 464068 196104 464120 196110
rect 464068 196046 464120 196052
rect 463976 195968 464028 195974
rect 463976 195910 464028 195916
rect 463988 193225 464016 195910
rect 463790 193216 463846 193225
rect 463790 193151 463846 193160
rect 463974 193216 464030 193225
rect 463974 193151 464030 193160
rect 463804 183598 463832 193151
rect 463792 183592 463844 183598
rect 463792 183534 463844 183540
rect 464068 183592 464120 183598
rect 464068 183534 464120 183540
rect 464080 176730 464108 183534
rect 463884 176724 463936 176730
rect 463884 176666 463936 176672
rect 464068 176724 464120 176730
rect 464068 176666 464120 176672
rect 463896 166954 463924 176666
rect 463804 166926 463924 166954
rect 463804 164218 463832 166926
rect 463792 164212 463844 164218
rect 463792 164154 463844 164160
rect 464068 164212 464120 164218
rect 464068 164154 464120 164160
rect 464080 154601 464108 164154
rect 463882 154592 463938 154601
rect 463882 154527 463938 154536
rect 464066 154592 464122 154601
rect 464066 154527 464122 154536
rect 463896 130422 463924 154527
rect 463884 130416 463936 130422
rect 463884 130358 463936 130364
rect 464068 130416 464120 130422
rect 464068 130358 464120 130364
rect 464080 125633 464108 130358
rect 463882 125624 463938 125633
rect 463882 125559 463938 125568
rect 464066 125624 464122 125633
rect 464066 125559 464122 125568
rect 463896 118726 463924 125559
rect 463884 118720 463936 118726
rect 463884 118662 463936 118668
rect 463976 118652 464028 118658
rect 463976 118594 464028 118600
rect 463988 109070 464016 118594
rect 463792 109064 463844 109070
rect 463792 109006 463844 109012
rect 463976 109064 464028 109070
rect 463976 109006 464028 109012
rect 463804 103578 463832 109006
rect 463804 103550 463924 103578
rect 463896 93906 463924 103550
rect 463700 93900 463752 93906
rect 463700 93842 463752 93848
rect 463884 93900 463936 93906
rect 463884 93842 463936 93848
rect 463712 93786 463740 93842
rect 463712 93758 463832 93786
rect 463804 80102 463832 93758
rect 463792 80096 463844 80102
rect 463792 80038 463844 80044
rect 463792 79960 463844 79966
rect 463792 79902 463844 79908
rect 463804 70394 463832 79902
rect 463712 70366 463832 70394
rect 463608 3664 463660 3670
rect 463608 3606 463660 3612
rect 463516 3596 463568 3602
rect 463516 3538 463568 3544
rect 463712 610 463740 70366
rect 465000 5098 465028 336738
rect 465920 331242 465948 340054
rect 465920 331214 466224 331242
rect 464988 5092 465040 5098
rect 464988 5034 465040 5040
rect 465632 5024 465684 5030
rect 465632 4966 465684 4972
rect 463700 604 463752 610
rect 463700 546 463752 552
rect 464436 604 464488 610
rect 464436 546 464488 552
rect 464448 480 464476 546
rect 465644 480 465672 4966
rect 466196 4962 466224 331214
rect 466184 4956 466236 4962
rect 466184 4898 466236 4904
rect 466288 3534 466316 340054
rect 466368 337340 466420 337346
rect 466368 337282 466420 337288
rect 466380 3602 466408 337282
rect 466564 336938 466592 340068
rect 467116 337958 467144 340068
rect 467104 337952 467156 337958
rect 467104 337894 467156 337900
rect 467576 337385 467604 340068
rect 468036 337958 468064 340068
rect 468602 340054 468984 340082
rect 467748 337952 467800 337958
rect 467748 337894 467800 337900
rect 468024 337952 468076 337958
rect 468024 337894 468076 337900
rect 467562 337376 467618 337385
rect 467562 337311 467618 337320
rect 466552 336932 466604 336938
rect 466552 336874 466604 336880
rect 467760 4865 467788 337894
rect 468760 8356 468812 8362
rect 468760 8298 468812 8304
rect 467746 4856 467802 4865
rect 467746 4791 467802 4800
rect 466368 3596 466420 3602
rect 466368 3538 466420 3544
rect 466276 3528 466328 3534
rect 466276 3470 466328 3476
rect 467932 3460 467984 3466
rect 467932 3402 467984 3408
rect 466828 2848 466880 2854
rect 466828 2790 466880 2796
rect 466840 480 466868 2790
rect 467944 480 467972 3402
rect 468772 3369 468800 8298
rect 468956 5574 468984 340054
rect 469048 8362 469076 340068
rect 469128 337952 469180 337958
rect 469128 337894 469180 337900
rect 469036 8356 469088 8362
rect 469036 8298 469088 8304
rect 469140 7970 469168 337894
rect 469508 337278 469536 340068
rect 469496 337272 469548 337278
rect 469496 337214 469548 337220
rect 469220 336864 469272 336870
rect 469220 336806 469272 336812
rect 469048 7942 469168 7970
rect 468944 5568 468996 5574
rect 468944 5510 468996 5516
rect 469048 3466 469076 7942
rect 469128 4888 469180 4894
rect 469128 4830 469180 4836
rect 469036 3460 469088 3466
rect 469036 3402 469088 3408
rect 468758 3360 468814 3369
rect 468758 3295 468814 3304
rect 469140 480 469168 4830
rect 469232 610 469260 336806
rect 469876 252550 469904 580246
rect 469968 299470 469996 580314
rect 470048 579216 470100 579222
rect 470048 579158 470100 579164
rect 470060 322930 470088 579158
rect 470152 346390 470180 581062
rect 470244 393310 470272 581130
rect 470324 579284 470376 579290
rect 470324 579226 470376 579232
rect 470336 405686 470364 579226
rect 470428 416770 470456 581198
rect 470520 440230 470548 581266
rect 471256 499526 471284 583578
rect 471348 546446 471376 583646
rect 580632 583568 580684 583574
rect 580632 583510 580684 583516
rect 580540 583500 580592 583506
rect 580540 583442 580592 583448
rect 580356 583432 580408 583438
rect 580356 583374 580408 583380
rect 580080 581052 580132 581058
rect 580080 580994 580132 581000
rect 580092 580122 580120 580994
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 580242 580212 580751
rect 580172 580236 580224 580242
rect 580172 580178 580224 580184
rect 580092 580094 580212 580122
rect 579804 579148 579856 579154
rect 579804 579090 579856 579096
rect 579712 557524 579764 557530
rect 579712 557466 579764 557472
rect 579724 557297 579752 557466
rect 579710 557288 579766 557297
rect 579710 557223 579766 557232
rect 471336 546440 471388 546446
rect 471336 546382 471388 546388
rect 579712 546440 579764 546446
rect 579712 546382 579764 546388
rect 579724 545601 579752 546382
rect 579710 545592 579766 545601
rect 579710 545527 579766 545536
rect 579712 510604 579764 510610
rect 579712 510546 579764 510552
rect 579724 510377 579752 510546
rect 579710 510368 579766 510377
rect 579710 510303 579766 510312
rect 471244 499520 471296 499526
rect 471244 499462 471296 499468
rect 579712 499520 579764 499526
rect 579712 499462 579764 499468
rect 579724 498681 579752 499462
rect 579710 498672 579766 498681
rect 579710 498607 579766 498616
rect 579712 463684 579764 463690
rect 579712 463626 579764 463632
rect 579724 463457 579752 463626
rect 579710 463448 579766 463457
rect 579710 463383 579766 463392
rect 579816 451761 579844 579090
rect 579988 579080 580040 579086
rect 579988 579022 580040 579028
rect 579896 579012 579948 579018
rect 579896 578954 579948 578960
rect 579802 451752 579858 451761
rect 579802 451687 579858 451696
rect 470508 440224 470560 440230
rect 470508 440166 470560 440172
rect 579804 440224 579856 440230
rect 579804 440166 579856 440172
rect 579816 439929 579844 440166
rect 579802 439920 579858 439929
rect 579802 439855 579858 439864
rect 470416 416764 470468 416770
rect 470416 416706 470468 416712
rect 579804 416764 579856 416770
rect 579804 416706 579856 416712
rect 579816 416537 579844 416706
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 470324 405680 470376 405686
rect 470324 405622 470376 405628
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404841 579844 405622
rect 579802 404832 579858 404841
rect 579802 404767 579858 404776
rect 470232 393304 470284 393310
rect 470232 393246 470284 393252
rect 579804 393304 579856 393310
rect 579804 393246 579856 393252
rect 579816 393009 579844 393246
rect 579802 393000 579858 393009
rect 579802 392935 579858 392944
rect 579908 369617 579936 578954
rect 579894 369608 579950 369617
rect 579894 369543 579950 369552
rect 580000 357921 580028 579022
rect 580080 578944 580132 578950
rect 580080 578886 580132 578892
rect 579986 357912 580042 357921
rect 579986 357847 580042 357856
rect 470140 346384 470192 346390
rect 470140 346326 470192 346332
rect 579988 346384 580040 346390
rect 579988 346326 580040 346332
rect 580000 346089 580028 346326
rect 579986 346080 580042 346089
rect 579986 346015 580042 346024
rect 499580 338088 499632 338094
rect 499580 338030 499632 338036
rect 470600 337340 470652 337346
rect 470600 337282 470652 337288
rect 470692 337340 470744 337346
rect 470692 337282 470744 337288
rect 470506 337240 470562 337249
rect 470506 337175 470562 337184
rect 470520 336938 470548 337175
rect 470508 336932 470560 336938
rect 470508 336874 470560 336880
rect 470612 328438 470640 337282
rect 470704 337249 470732 337282
rect 470690 337240 470746 337249
rect 470690 337175 470746 337184
rect 492680 337204 492732 337210
rect 492680 337146 492732 337152
rect 485780 337136 485832 337142
rect 485780 337078 485832 337084
rect 477592 337068 477644 337074
rect 477592 337010 477644 337016
rect 475384 337000 475436 337006
rect 475384 336942 475436 336948
rect 470600 328432 470652 328438
rect 470600 328374 470652 328380
rect 470048 322924 470100 322930
rect 470048 322866 470100 322872
rect 470600 318844 470652 318850
rect 470600 318786 470652 318792
rect 470612 309126 470640 318786
rect 470600 309120 470652 309126
rect 470600 309062 470652 309068
rect 470600 299532 470652 299538
rect 470600 299474 470652 299480
rect 469956 299464 470008 299470
rect 469956 299406 470008 299412
rect 470612 289814 470640 299474
rect 470600 289808 470652 289814
rect 470600 289750 470652 289756
rect 470600 280220 470652 280226
rect 470600 280162 470652 280168
rect 470612 270502 470640 280162
rect 470600 270496 470652 270502
rect 470600 270438 470652 270444
rect 470600 260908 470652 260914
rect 470600 260850 470652 260856
rect 469864 252544 469916 252550
rect 469864 252486 469916 252492
rect 470612 251190 470640 260850
rect 470600 251184 470652 251190
rect 470600 251126 470652 251132
rect 470600 241528 470652 241534
rect 470600 241470 470652 241476
rect 470612 231849 470640 241470
rect 470414 231840 470470 231849
rect 470414 231775 470470 231784
rect 470598 231840 470654 231849
rect 470598 231775 470654 231784
rect 470428 222222 470456 231775
rect 470416 222216 470468 222222
rect 470416 222158 470468 222164
rect 470600 222216 470652 222222
rect 470600 222158 470652 222164
rect 470612 212537 470640 222158
rect 470414 212528 470470 212537
rect 470414 212463 470470 212472
rect 470598 212528 470654 212537
rect 470598 212463 470654 212472
rect 470428 202910 470456 212463
rect 470416 202904 470468 202910
rect 470416 202846 470468 202852
rect 470600 202904 470652 202910
rect 470600 202846 470652 202852
rect 470612 193225 470640 202846
rect 470414 193216 470470 193225
rect 470414 193151 470470 193160
rect 470598 193216 470654 193225
rect 470598 193151 470654 193160
rect 470428 183598 470456 193151
rect 470416 183592 470468 183598
rect 470416 183534 470468 183540
rect 470600 183592 470652 183598
rect 470600 183534 470652 183540
rect 470612 173913 470640 183534
rect 470414 173904 470470 173913
rect 470414 173839 470470 173848
rect 470598 173904 470654 173913
rect 470598 173839 470654 173848
rect 470428 164257 470456 173839
rect 470414 164248 470470 164257
rect 470414 164183 470470 164192
rect 470598 164248 470654 164257
rect 470598 164183 470654 164192
rect 470612 154562 470640 164183
rect 470416 154556 470468 154562
rect 470416 154498 470468 154504
rect 470600 154556 470652 154562
rect 470600 154498 470652 154504
rect 470428 144945 470456 154498
rect 470414 144936 470470 144945
rect 470414 144871 470470 144880
rect 470598 144936 470654 144945
rect 470598 144871 470654 144880
rect 470612 135250 470640 144871
rect 470416 135244 470468 135250
rect 470416 135186 470468 135192
rect 470600 135244 470652 135250
rect 470600 135186 470652 135192
rect 470428 125633 470456 135186
rect 470414 125624 470470 125633
rect 470414 125559 470470 125568
rect 470598 125624 470654 125633
rect 470598 125559 470654 125568
rect 470612 57934 470640 125559
rect 470600 57928 470652 57934
rect 470600 57870 470652 57876
rect 470600 48340 470652 48346
rect 470600 48282 470652 48288
rect 470612 5642 470640 48282
rect 470600 5636 470652 5642
rect 470600 5578 470652 5584
rect 472716 4208 472768 4214
rect 472716 4150 472768 4156
rect 469220 604 469272 610
rect 469220 546 469272 552
rect 470324 604 470376 610
rect 470324 546 470376 552
rect 471520 604 471572 610
rect 471520 546 471572 552
rect 470336 480 470364 546
rect 471532 480 471560 546
rect 472728 480 472756 4150
rect 475396 3126 475424 336942
rect 476026 87272 476082 87281
rect 476026 87207 476082 87216
rect 476040 87122 476068 87207
rect 476210 87136 476266 87145
rect 476040 87094 476210 87122
rect 476210 87071 476266 87080
rect 476026 29336 476082 29345
rect 476026 29271 476082 29280
rect 476040 29186 476068 29271
rect 476210 29200 476266 29209
rect 476040 29158 476210 29186
rect 476210 29135 476266 29144
rect 476304 5772 476356 5778
rect 476304 5714 476356 5720
rect 475108 3120 475160 3126
rect 475108 3062 475160 3068
rect 475384 3120 475436 3126
rect 475384 3062 475436 3068
rect 473912 2916 473964 2922
rect 473912 2858 473964 2864
rect 473924 480 473952 2858
rect 475120 480 475148 3062
rect 476316 480 476344 5714
rect 477604 3346 477632 337010
rect 482926 111072 482982 111081
rect 482926 111007 482982 111016
rect 482940 110673 482968 111007
rect 482926 110664 482982 110673
rect 482926 110599 482982 110608
rect 482926 76528 482982 76537
rect 482926 76463 482982 76472
rect 482940 76129 482968 76463
rect 482926 76120 482982 76129
rect 482926 76055 482982 76064
rect 482926 17232 482982 17241
rect 482926 17167 482982 17176
rect 482940 16833 482968 17167
rect 482926 16824 482982 16833
rect 482926 16759 482982 16768
rect 483480 5976 483532 5982
rect 483480 5918 483532 5924
rect 479892 5840 479944 5846
rect 479892 5782 479944 5788
rect 477604 3318 478736 3346
rect 477500 3120 477552 3126
rect 477500 3062 477552 3068
rect 477512 480 477540 3062
rect 478708 480 478736 3318
rect 479904 480 479932 5782
rect 482284 3120 482336 3126
rect 482284 3062 482336 3068
rect 481088 2984 481140 2990
rect 481088 2926 481140 2932
rect 481100 480 481128 2926
rect 482296 480 482324 3062
rect 483492 480 483520 5918
rect 484584 5908 484636 5914
rect 484584 5850 484636 5856
rect 484596 480 484624 5850
rect 485792 480 485820 337078
rect 487802 110936 487858 110945
rect 487802 110871 487858 110880
rect 487816 110537 487844 110871
rect 487802 110528 487858 110537
rect 487802 110463 487858 110472
rect 491206 87408 491262 87417
rect 491206 87343 491262 87352
rect 491220 87009 491248 87343
rect 491206 87000 491262 87009
rect 491206 86935 491262 86944
rect 487802 76392 487858 76401
rect 487802 76327 487858 76336
rect 487816 75993 487844 76327
rect 487802 75984 487858 75993
rect 487802 75919 487858 75928
rect 491206 29472 491262 29481
rect 491206 29407 491262 29416
rect 491220 29073 491248 29407
rect 491206 29064 491262 29073
rect 491206 28999 491262 29008
rect 487802 17096 487858 17105
rect 487802 17031 487858 17040
rect 487816 16697 487844 17031
rect 487802 16688 487858 16697
rect 487802 16623 487858 16632
rect 491760 6860 491812 6866
rect 491760 6802 491812 6808
rect 490564 6792 490616 6798
rect 490564 6734 490616 6740
rect 486976 6112 487028 6118
rect 486976 6054 487028 6060
rect 486988 480 487016 6054
rect 488172 6044 488224 6050
rect 488172 5986 488224 5992
rect 488184 480 488212 5986
rect 489368 3052 489420 3058
rect 489368 2994 489420 3000
rect 489380 480 489408 2994
rect 490576 480 490604 6734
rect 491772 480 491800 6802
rect 492692 3482 492720 337146
rect 494612 87168 494664 87174
rect 494612 87110 494664 87116
rect 494624 87009 494652 87110
rect 494610 87000 494666 87009
rect 494610 86935 494666 86944
rect 492772 29096 492824 29102
rect 492770 29064 492772 29073
rect 492824 29064 492826 29073
rect 492770 28999 492826 29008
rect 495348 6724 495400 6730
rect 495348 6666 495400 6672
rect 494152 6656 494204 6662
rect 494152 6598 494204 6604
rect 492692 3454 492996 3482
rect 492968 480 492996 3454
rect 494164 480 494192 6598
rect 495360 480 495388 6666
rect 497740 6588 497792 6594
rect 497740 6530 497792 6536
rect 496544 3256 496596 3262
rect 496544 3198 496596 3204
rect 496556 480 496584 3198
rect 497752 480 497780 6530
rect 498936 6520 498988 6526
rect 498936 6462 498988 6468
rect 498948 480 498976 6462
rect 499592 3482 499620 338030
rect 525064 338020 525116 338026
rect 525064 337962 525116 337968
rect 523684 337884 523736 337890
rect 523684 337826 523736 337832
rect 521016 337816 521068 337822
rect 521016 337758 521068 337764
rect 506480 337748 506532 337754
rect 506480 337690 506532 337696
rect 505744 336796 505796 336802
rect 505744 336738 505796 336744
rect 502246 87272 502302 87281
rect 502246 87207 502302 87216
rect 502260 87174 502288 87207
rect 502248 87168 502300 87174
rect 502248 87110 502300 87116
rect 502246 29336 502302 29345
rect 502246 29271 502302 29280
rect 502260 29102 502288 29271
rect 502248 29096 502300 29102
rect 502248 29038 502300 29044
rect 501236 6452 501288 6458
rect 501236 6394 501288 6400
rect 499592 3454 500172 3482
rect 500144 480 500172 3454
rect 501248 480 501276 6394
rect 502432 6384 502484 6390
rect 502432 6326 502484 6332
rect 502444 480 502472 6326
rect 504824 6316 504876 6322
rect 504824 6258 504876 6264
rect 503628 3324 503680 3330
rect 503628 3266 503680 3272
rect 503640 480 503668 3266
rect 504836 480 504864 6258
rect 505756 3194 505784 336738
rect 506020 6248 506072 6254
rect 506020 6190 506072 6196
rect 505744 3188 505796 3194
rect 505744 3130 505796 3136
rect 506032 480 506060 6190
rect 506492 3482 506520 337690
rect 518164 337680 518216 337686
rect 518164 337622 518216 337628
rect 516784 337544 516836 337550
rect 516784 337486 516836 337492
rect 514024 337476 514076 337482
rect 514024 337418 514076 337424
rect 509240 337408 509292 337414
rect 509240 337350 509292 337356
rect 512642 337376 512698 337385
rect 509252 337210 509280 337350
rect 512642 337311 512698 337320
rect 509240 337204 509292 337210
rect 509240 337146 509292 337152
rect 510620 337204 510672 337210
rect 510620 337146 510672 337152
rect 509884 336864 509936 336870
rect 509884 336806 509936 336812
rect 509608 7336 509660 7342
rect 509608 7278 509660 7284
rect 508412 6180 508464 6186
rect 508412 6122 508464 6128
rect 506492 3454 507256 3482
rect 507228 480 507256 3454
rect 508424 480 508452 6122
rect 509620 480 509648 7278
rect 509896 3058 509924 336806
rect 510632 3482 510660 337146
rect 512000 4276 512052 4282
rect 512000 4218 512052 4224
rect 510632 3454 510844 3482
rect 509884 3052 509936 3058
rect 509884 2994 509936 3000
rect 510816 480 510844 3454
rect 512012 480 512040 4218
rect 512656 3262 512684 337311
rect 513196 7404 513248 7410
rect 513196 7346 513248 7352
rect 512644 3256 512696 3262
rect 512644 3198 512696 3204
rect 513208 480 513236 7346
rect 514036 3398 514064 337418
rect 516796 11778 516824 337486
rect 516704 11750 516824 11778
rect 516704 6934 516732 11750
rect 516784 7472 516836 7478
rect 516784 7414 516836 7420
rect 516692 6928 516744 6934
rect 516692 6870 516744 6876
rect 515588 4344 515640 4350
rect 515588 4286 515640 4292
rect 514024 3392 514076 3398
rect 514024 3334 514076 3340
rect 514392 3324 514444 3330
rect 514392 3266 514444 3272
rect 514404 480 514432 3266
rect 515600 480 515628 4286
rect 516796 480 516824 7414
rect 516876 6928 516928 6934
rect 516876 6870 516928 6876
rect 516888 3330 516916 6870
rect 517888 3392 517940 3398
rect 517888 3334 517940 3340
rect 516876 3324 516928 3330
rect 516876 3266 516928 3272
rect 517900 480 517928 3334
rect 518176 2854 518204 337622
rect 520924 337612 520976 337618
rect 520924 337554 520976 337560
rect 520280 7540 520332 7546
rect 520280 7482 520332 7488
rect 519084 4412 519136 4418
rect 519084 4354 519136 4360
rect 518164 2848 518216 2854
rect 518164 2790 518216 2796
rect 519096 480 519124 4354
rect 520292 480 520320 7482
rect 520936 2922 520964 337554
rect 521028 2990 521056 337758
rect 522672 4480 522724 4486
rect 522672 4422 522724 4428
rect 521476 4140 521528 4146
rect 521476 4082 521528 4088
rect 521016 2984 521068 2990
rect 521016 2926 521068 2932
rect 520924 2916 520976 2922
rect 520924 2858 520976 2864
rect 521488 480 521516 4082
rect 522684 480 522712 4422
rect 523696 3058 523724 337826
rect 523868 8288 523920 8294
rect 523868 8230 523920 8236
rect 523684 3052 523736 3058
rect 523684 2994 523736 3000
rect 523880 480 523908 8230
rect 525076 6882 525104 337962
rect 527824 337952 527876 337958
rect 527824 337894 527876 337900
rect 527456 8220 527508 8226
rect 527456 8162 527508 8168
rect 524984 6854 525104 6882
rect 524984 3126 525012 6854
rect 526260 4548 526312 4554
rect 526260 4490 526312 4496
rect 525064 3392 525116 3398
rect 525064 3334 525116 3340
rect 524972 3120 525024 3126
rect 524972 3062 525024 3068
rect 525076 480 525104 3334
rect 526272 480 526300 4490
rect 527468 480 527496 8162
rect 527836 3398 527864 337894
rect 529204 337340 529256 337346
rect 529204 337282 529256 337288
rect 529216 4146 529244 337282
rect 530584 337272 530636 337278
rect 530584 337214 530636 337220
rect 529848 4616 529900 4622
rect 529848 4558 529900 4564
rect 529204 4140 529256 4146
rect 529204 4082 529256 4088
rect 528652 4072 528704 4078
rect 528652 4014 528704 4020
rect 527824 3392 527876 3398
rect 527824 3334 527876 3340
rect 528664 480 528692 4014
rect 529860 480 529888 4558
rect 530596 4078 530624 337214
rect 579988 322924 580040 322930
rect 579988 322866 580040 322872
rect 580000 322697 580028 322866
rect 579986 322688 580042 322697
rect 579986 322623 580042 322632
rect 580092 310865 580120 578886
rect 580078 310856 580134 310865
rect 580078 310791 580134 310800
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 580184 275777 580212 580094
rect 580264 578604 580316 578610
rect 580264 578546 580316 578552
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 252544 580224 252550
rect 580172 252486 580224 252492
rect 580184 252249 580212 252486
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580276 123185 580304 578546
rect 580368 134881 580396 583374
rect 580448 578672 580500 578678
rect 580448 578614 580500 578620
rect 580460 170105 580488 578614
rect 580552 181937 580580 583442
rect 580644 205329 580672 583510
rect 580908 578876 580960 578882
rect 580908 578818 580960 578824
rect 580724 578808 580776 578814
rect 580724 578750 580776 578756
rect 580736 217025 580764 578750
rect 580816 578740 580868 578746
rect 580816 578682 580868 578688
rect 580828 228857 580856 578682
rect 580920 263945 580948 578818
rect 580906 263936 580962 263945
rect 580906 263871 580962 263880
rect 580814 228848 580870 228857
rect 580814 228783 580870 228792
rect 580722 217016 580778 217025
rect 580722 216951 580778 216960
rect 580630 205320 580686 205329
rect 580630 205255 580686 205264
rect 580538 181928 580594 181937
rect 580538 181863 580594 181872
rect 580446 170096 580502 170105
rect 580446 170031 580502 170040
rect 580354 134872 580410 134881
rect 580354 134807 580410 134816
rect 580262 123176 580318 123185
rect 580262 123111 580318 123120
rect 531044 8152 531096 8158
rect 531044 8094 531096 8100
rect 530584 4072 530636 4078
rect 530584 4014 530636 4020
rect 531056 480 531084 8094
rect 534540 8084 534592 8090
rect 534540 8026 534592 8032
rect 533436 4684 533488 4690
rect 533436 4626 533488 4632
rect 532240 2848 532292 2854
rect 532240 2790 532292 2796
rect 532252 480 532280 2790
rect 533448 480 533476 4626
rect 534552 480 534580 8026
rect 538128 8016 538180 8022
rect 538128 7958 538180 7964
rect 536932 4752 536984 4758
rect 536932 4694 536984 4700
rect 535736 4004 535788 4010
rect 535736 3946 535788 3952
rect 535748 480 535776 3946
rect 536944 480 536972 4694
rect 538140 480 538168 7958
rect 541716 7948 541768 7954
rect 541716 7890 541768 7896
rect 540520 5500 540572 5506
rect 540520 5442 540572 5448
rect 539324 2916 539376 2922
rect 539324 2858 539376 2864
rect 539336 480 539364 2858
rect 540532 480 540560 5442
rect 541728 480 541756 7890
rect 545304 7880 545356 7886
rect 545304 7822 545356 7828
rect 544108 5432 544160 5438
rect 544108 5374 544160 5380
rect 542912 3936 542964 3942
rect 542912 3878 542964 3884
rect 542924 480 542952 3878
rect 544120 480 544148 5374
rect 545316 480 545344 7822
rect 548892 7812 548944 7818
rect 548892 7754 548944 7760
rect 547696 5364 547748 5370
rect 547696 5306 547748 5312
rect 546500 2984 546552 2990
rect 546500 2926 546552 2932
rect 546512 480 546540 2926
rect 547708 480 547736 5306
rect 548904 480 548932 7754
rect 552388 7744 552440 7750
rect 552388 7686 552440 7692
rect 551192 5296 551244 5302
rect 551192 5238 551244 5244
rect 550088 3868 550140 3874
rect 550088 3810 550140 3816
rect 550100 480 550128 3810
rect 551204 480 551232 5238
rect 552400 480 552428 7686
rect 555976 7676 556028 7682
rect 555976 7618 556028 7624
rect 554780 5228 554832 5234
rect 554780 5170 554832 5176
rect 553584 3052 553636 3058
rect 553584 2994 553636 3000
rect 553596 480 553624 2994
rect 554792 480 554820 5170
rect 555988 480 556016 7618
rect 559564 7608 559616 7614
rect 559564 7550 559616 7556
rect 558368 5160 558420 5166
rect 558368 5102 558420 5108
rect 557172 3800 557224 3806
rect 557172 3742 557224 3748
rect 557184 480 557212 3742
rect 558380 480 558408 5102
rect 559576 480 559604 7550
rect 561956 5092 562008 5098
rect 561956 5034 562008 5040
rect 560760 3120 560812 3126
rect 560760 3062 560812 3068
rect 560772 480 560800 3062
rect 561968 480 561996 5034
rect 565544 5024 565596 5030
rect 565544 4966 565596 4972
rect 564348 3732 564400 3738
rect 564348 3674 564400 3680
rect 563152 3188 563204 3194
rect 563152 3130 563204 3136
rect 563164 480 563192 3130
rect 564360 480 564388 3674
rect 565556 480 565584 4966
rect 569040 4956 569092 4962
rect 569040 4898 569092 4904
rect 566740 3664 566792 3670
rect 566740 3606 566792 3612
rect 566752 480 566780 3606
rect 567844 3392 567896 3398
rect 567844 3334 567896 3340
rect 567856 480 567884 3334
rect 569052 480 569080 4898
rect 572628 4888 572680 4894
rect 572628 4830 572680 4836
rect 576214 4856 576270 4865
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 570236 3256 570288 3262
rect 570236 3198 570288 3204
rect 570248 480 570276 3198
rect 571444 480 571472 3538
rect 572640 480 572668 4830
rect 576214 4791 576270 4800
rect 579804 4820 579856 4826
rect 575020 4140 575072 4146
rect 575020 4082 575072 4088
rect 573824 3528 573876 3534
rect 573824 3470 573876 3476
rect 573836 480 573864 3470
rect 575032 480 575060 4082
rect 576228 480 576256 4791
rect 579804 4762 579856 4768
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 577412 3324 577464 3330
rect 577412 3266 577464 3272
rect 577424 480 577452 3266
rect 578620 480 578648 3402
rect 579816 480 579844 4762
rect 582196 4072 582248 4078
rect 582196 4014 582248 4020
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 4014
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 4802 583480 4858 583536
rect 3054 567332 3056 567352
rect 3056 567332 3108 567352
rect 3108 567332 3110 567352
rect 3054 567296 3110 567332
rect 2778 553052 2780 553072
rect 2780 553052 2832 553072
rect 2832 553052 2834 553072
rect 2778 553016 2834 553052
rect 3054 538636 3056 538656
rect 3056 538636 3108 538656
rect 3108 538636 3110 538656
rect 3054 538600 3110 538636
rect 3054 509904 3110 509960
rect 2778 495488 2834 495544
rect 2962 481108 2964 481128
rect 2964 481108 3016 481128
rect 3016 481108 3018 481128
rect 2962 481072 3018 481108
rect 3146 452376 3202 452432
rect 3146 437960 3202 438016
rect 3146 423680 3202 423736
rect 3238 394984 3294 395040
rect 3238 380568 3294 380624
rect 3330 366152 3386 366208
rect 3330 323040 3386 323096
rect 2778 308796 2780 308816
rect 2780 308796 2832 308816
rect 2832 308796 2834 308816
rect 2778 308760 2834 308796
rect 2962 295160 3018 295216
rect 2962 294344 3018 294400
rect 2778 251232 2834 251288
rect 3054 236952 3110 237008
rect 2778 165008 2834 165064
rect 3330 150728 3386 150784
rect 2778 136312 2834 136368
rect 2778 122032 2834 122088
rect 4066 280064 4122 280120
rect 3974 265648 4030 265704
rect 3882 222536 3938 222592
rect 3790 208120 3846 208176
rect 3698 193840 3754 193896
rect 3606 179424 3662 179480
rect 3514 107616 3570 107672
rect 3422 93200 3478 93256
rect 2778 78920 2834 78976
rect 3330 64504 3386 64560
rect 5078 582528 5134 582584
rect 2778 50088 2834 50144
rect 10322 337320 10378 337376
rect 3146 35844 3148 35864
rect 3148 35844 3200 35864
rect 3200 35844 3202 35864
rect 3146 35808 3202 35844
rect 3146 11600 3202 11656
rect 3146 7112 3202 7168
rect 6458 3304 6514 3360
rect 17222 582800 17278 582856
rect 24122 582664 24178 582720
rect 293958 583208 294014 583264
rect 300306 583344 300362 583400
rect 378138 700304 378194 700360
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 460294 583480 460350 583536
rect 420274 583072 420330 583128
rect 426622 582936 426678 582992
rect 449806 582800 449862 582856
rect 447690 582528 447746 582584
rect 462410 582664 462466 582720
rect 468482 579672 468538 579728
rect 231122 579264 231178 579320
rect 232962 579264 233018 579320
rect 235262 579264 235318 579320
rect 237194 579264 237250 579320
rect 239402 579264 239458 579320
rect 241426 579264 241482 579320
rect 243634 579264 243690 579320
rect 249522 579264 249578 579320
rect 466458 579264 466514 579320
rect 51630 6160 51686 6216
rect 57978 337748 58034 337784
rect 57978 337728 57980 337748
rect 57980 337728 58032 337748
rect 58032 337728 58034 337748
rect 67546 337748 67602 337784
rect 67546 337728 67548 337748
rect 67548 337728 67600 337748
rect 67600 337728 67602 337748
rect 77298 337748 77354 337784
rect 77298 337728 77300 337748
rect 77300 337728 77352 337748
rect 77352 337728 77354 337748
rect 86866 337748 86922 337784
rect 86866 337728 86868 337748
rect 86868 337728 86920 337748
rect 86920 337728 86922 337748
rect 95238 337748 95294 337784
rect 95238 337728 95240 337748
rect 95240 337728 95292 337748
rect 95292 337728 95294 337748
rect 104806 337748 104862 337784
rect 104806 337728 104808 337748
rect 104808 337728 104860 337748
rect 104860 337728 104862 337748
rect 114558 337748 114614 337784
rect 114558 337728 114560 337748
rect 114560 337728 114612 337748
rect 114612 337728 114614 337748
rect 124126 337748 124182 337784
rect 124126 337728 124128 337748
rect 124128 337728 124180 337748
rect 124180 337728 124182 337748
rect 133878 337748 133934 337784
rect 133878 337728 133880 337748
rect 133880 337728 133932 337748
rect 133932 337728 133934 337748
rect 143446 337748 143502 337784
rect 143446 337728 143448 337748
rect 143448 337728 143500 337748
rect 143500 337728 143502 337748
rect 153198 337748 153254 337784
rect 153198 337728 153200 337748
rect 153200 337728 153252 337748
rect 153252 337728 153254 337748
rect 162766 337748 162822 337784
rect 162766 337728 162768 337748
rect 162768 337728 162820 337748
rect 162820 337728 162822 337748
rect 172518 337748 172574 337784
rect 172518 337728 172520 337748
rect 172520 337728 172572 337748
rect 172572 337728 172574 337748
rect 182086 337748 182142 337784
rect 182086 337728 182088 337748
rect 182088 337728 182140 337748
rect 182140 337728 182142 337748
rect 191838 337748 191894 337784
rect 191838 337728 191840 337748
rect 191840 337728 191892 337748
rect 191892 337728 191894 337748
rect 201406 337748 201462 337784
rect 201406 337728 201408 337748
rect 201408 337728 201460 337748
rect 201460 337728 201462 337748
rect 211158 337748 211214 337784
rect 211158 337728 211160 337748
rect 211160 337728 211212 337748
rect 211212 337728 211214 337748
rect 220726 337748 220782 337784
rect 220726 337728 220728 337748
rect 220728 337728 220780 337748
rect 220780 337728 220782 337748
rect 132498 337220 132500 337240
rect 132500 337220 132552 337240
rect 132552 337220 132554 337240
rect 132498 337184 132554 337220
rect 142066 337220 142068 337240
rect 142068 337220 142120 337240
rect 142120 337220 142122 337240
rect 142066 337184 142122 337220
rect 151818 337220 151820 337240
rect 151820 337220 151872 337240
rect 151872 337220 151874 337240
rect 151818 337184 151874 337220
rect 161386 337220 161388 337240
rect 161388 337220 161440 337240
rect 161440 337220 161442 337240
rect 161386 337184 161442 337220
rect 171138 337220 171140 337240
rect 171140 337220 171192 337240
rect 171192 337220 171194 337240
rect 171138 337184 171194 337220
rect 180706 337220 180708 337240
rect 180708 337220 180760 337240
rect 180760 337220 180762 337240
rect 180706 337184 180762 337220
rect 190458 337220 190460 337240
rect 190460 337220 190512 337240
rect 190512 337220 190514 337240
rect 190458 337184 190514 337220
rect 200026 337220 200028 337240
rect 200028 337220 200080 337240
rect 200080 337220 200082 337240
rect 200026 337184 200082 337220
rect 209778 337220 209780 337240
rect 209780 337220 209832 337240
rect 209832 337220 209834 337240
rect 209778 337184 209834 337220
rect 219346 337220 219348 337240
rect 219348 337220 219400 337240
rect 219400 337220 219402 337240
rect 219346 337184 219402 337220
rect 221002 337220 221004 337240
rect 221004 337220 221056 337240
rect 221056 337220 221058 337240
rect 221002 337184 221058 337220
rect 132590 8880 132646 8936
rect 129002 7520 129058 7576
rect 208674 4800 208730 4856
rect 231950 337320 232006 337376
rect 232226 318824 232282 318880
rect 232410 318824 232466 318880
rect 232226 249736 232282 249792
rect 232502 249736 232558 249792
rect 232226 230424 232282 230480
rect 232502 230424 232558 230480
rect 232042 3304 232098 3360
rect 234618 337220 234620 337240
rect 234620 337220 234672 337240
rect 234672 337220 234674 337240
rect 234618 337184 234674 337220
rect 236274 172488 236330 172544
rect 236458 172488 236514 172544
rect 236274 135224 236330 135280
rect 236458 135224 236514 135280
rect 236274 115912 236330 115968
rect 236458 115912 236514 115968
rect 236274 96600 236330 96656
rect 236642 96600 236698 96656
rect 238758 29164 238814 29200
rect 238758 29144 238760 29164
rect 238760 29144 238812 29164
rect 238812 29144 238814 29164
rect 239310 240080 239366 240136
rect 239494 240080 239550 240136
rect 239126 212472 239182 212528
rect 239310 212472 239366 212528
rect 239034 201456 239090 201512
rect 239218 201456 239274 201512
rect 239126 138080 239182 138136
rect 239126 135244 239182 135280
rect 239126 135224 239128 135244
rect 239128 135224 239180 135244
rect 239180 135224 239182 135244
rect 239126 115912 239182 115968
rect 239310 115912 239366 115968
rect 239126 96600 239182 96656
rect 239310 96600 239366 96656
rect 244462 267688 244518 267744
rect 244646 267688 244702 267744
rect 244278 219408 244334 219464
rect 244554 219428 244610 219464
rect 244554 219408 244556 219428
rect 244556 219408 244608 219428
rect 244608 219408 244610 219428
rect 244462 145016 244518 145072
rect 244462 144880 244518 144936
rect 245566 48320 245622 48376
rect 245566 48184 245622 48240
rect 245934 325624 245990 325680
rect 246118 325624 246174 325680
rect 245842 316004 245844 316024
rect 245844 316004 245896 316024
rect 245896 316004 245898 316024
rect 245842 315968 245898 316004
rect 245934 315832 245990 315888
rect 245934 267688 245990 267744
rect 246118 267688 246174 267744
rect 245842 258032 245898 258088
rect 246118 258032 246174 258088
rect 245842 240116 245844 240136
rect 245844 240116 245896 240136
rect 245896 240116 245898 240136
rect 245842 240080 245898 240116
rect 246118 240080 246174 240136
rect 245934 164192 245990 164248
rect 245842 164056 245898 164112
rect 245842 133864 245898 133920
rect 246118 133864 246174 133920
rect 245934 125568 245990 125624
rect 246118 125568 246174 125624
rect 249246 336640 249302 336696
rect 249246 316240 249302 316296
rect 249246 306312 249302 306368
rect 249246 296928 249302 296984
rect 249430 275032 249486 275088
rect 249430 267824 249486 267880
rect 249246 257896 249302 257952
rect 249246 248376 249302 248432
rect 249614 209616 249670 209672
rect 249614 200096 249670 200152
rect 249338 193160 249394 193216
rect 249338 182144 249394 182200
rect 250074 278704 250130 278760
rect 250258 278704 250314 278760
rect 250074 193196 250076 193216
rect 250076 193196 250128 193216
rect 250128 193196 250130 193216
rect 250074 193160 250130 193196
rect 250258 193196 250260 193216
rect 250260 193196 250312 193216
rect 250312 193196 250314 193216
rect 250258 193160 250314 193196
rect 249982 6160 250038 6216
rect 251178 280064 251234 280120
rect 251178 260752 251234 260808
rect 251086 240080 251142 240136
rect 251178 162832 251234 162888
rect 251086 87488 251142 87544
rect 251086 87216 251142 87272
rect 251178 87100 251234 87136
rect 251178 87080 251180 87100
rect 251180 87080 251232 87100
rect 251232 87080 251234 87100
rect 251086 76064 251142 76120
rect 251086 75656 251142 75712
rect 251546 307672 251602 307728
rect 251546 298152 251602 298208
rect 251362 280064 251418 280120
rect 251362 260752 251418 260808
rect 251362 240116 251364 240136
rect 251364 240116 251416 240136
rect 251416 240116 251418 240136
rect 251362 240080 251418 240116
rect 251362 230460 251364 230480
rect 251364 230460 251416 230480
rect 251416 230460 251418 230480
rect 251362 230424 251418 230460
rect 251546 230424 251602 230480
rect 251362 162832 251418 162888
rect 251454 143520 251510 143576
rect 251638 143520 251694 143576
rect 251454 48456 251510 48512
rect 251362 48320 251418 48376
rect 251362 26288 251418 26344
rect 251638 26152 251694 26208
rect 256606 29008 256662 29064
rect 257986 29280 258042 29336
rect 257986 29008 258042 29064
rect 259366 63960 259422 64016
rect 259366 63552 259422 63608
rect 259734 306312 259790 306368
rect 259918 306312 259974 306368
rect 259642 295296 259698 295352
rect 259918 295296 259974 295352
rect 259734 258032 259790 258088
rect 259918 258032 259974 258088
rect 259642 240080 259698 240136
rect 259826 240080 259882 240136
rect 259642 222128 259698 222184
rect 259734 221856 259790 221912
rect 259642 202816 259698 202872
rect 259918 202816 259974 202872
rect 259550 96600 259606 96656
rect 259734 96600 259790 96656
rect 260654 87100 260710 87136
rect 260654 87080 260656 87100
rect 260656 87080 260708 87100
rect 260708 87080 260710 87100
rect 263414 29280 263470 29336
rect 263598 29280 263654 29336
rect 264978 314608 265034 314664
rect 264978 304952 265034 305008
rect 264978 258032 265034 258088
rect 265162 314608 265218 314664
rect 265254 304952 265310 305008
rect 265162 258032 265218 258088
rect 267830 315968 267886 316024
rect 268014 315968 268070 316024
rect 267738 277344 267794 277400
rect 268014 277344 268070 277400
rect 267922 240080 267978 240136
rect 268106 240080 268162 240136
rect 267738 183540 267740 183560
rect 267740 183540 267792 183560
rect 267792 183540 267794 183560
rect 267738 183504 267794 183540
rect 267922 183504 267978 183560
rect 266634 135224 266690 135280
rect 266818 135224 266874 135280
rect 266634 115912 266690 115968
rect 266818 115912 266874 115968
rect 266726 96736 266782 96792
rect 266634 96600 266690 96656
rect 267738 29180 267740 29200
rect 267740 29180 267792 29200
rect 267792 29180 267794 29200
rect 267738 29144 267794 29180
rect 265254 9560 265310 9616
rect 265438 9560 265494 9616
rect 270498 183504 270554 183560
rect 270498 164192 270554 164248
rect 270682 202816 270738 202872
rect 270682 202680 270738 202736
rect 270682 183540 270684 183560
rect 270684 183540 270736 183560
rect 270736 183540 270738 183560
rect 270682 183504 270738 183540
rect 270682 164192 270738 164248
rect 270682 125588 270738 125624
rect 270682 125568 270684 125588
rect 270684 125568 270736 125588
rect 270736 125568 270738 125588
rect 270958 125588 271014 125624
rect 270958 125568 270960 125588
rect 270960 125568 271012 125588
rect 271012 125568 271014 125588
rect 272154 278704 272210 278760
rect 272338 278704 272394 278760
rect 272154 241440 272210 241496
rect 272338 241304 272394 241360
rect 272154 222128 272210 222184
rect 272246 221992 272302 222048
rect 272154 202816 272210 202872
rect 272246 202680 272302 202736
rect 272062 164192 272118 164248
rect 272246 164192 272302 164248
rect 272154 133864 272210 133920
rect 272338 133864 272394 133920
rect 273074 315968 273130 316024
rect 273258 315968 273314 316024
rect 275558 63824 275614 63880
rect 275558 63552 275614 63608
rect 277306 29280 277362 29336
rect 278778 110744 278834 110800
rect 278778 110608 278834 110664
rect 279974 40296 280030 40352
rect 280158 40296 280214 40352
rect 283102 7520 283158 7576
rect 283470 87080 283526 87136
rect 283654 87080 283710 87136
rect 284574 278704 284630 278760
rect 284758 278704 284814 278760
rect 284666 220768 284722 220824
rect 284850 220768 284906 220824
rect 284482 8880 284538 8936
rect 285770 202816 285826 202872
rect 286046 261024 286102 261080
rect 285954 260888 286010 260944
rect 286046 249772 286048 249792
rect 286048 249772 286100 249792
rect 286100 249772 286102 249792
rect 286046 249736 286102 249772
rect 285954 249600 286010 249656
rect 285954 222128 286010 222184
rect 286138 222128 286194 222184
rect 285954 220768 286010 220824
rect 286138 220768 286194 220824
rect 285954 202852 285956 202872
rect 285956 202852 286008 202872
rect 286008 202852 286010 202872
rect 285954 202816 286010 202852
rect 285954 124072 286010 124128
rect 286230 123936 286286 123992
rect 288346 16768 288402 16824
rect 288346 16224 288402 16280
rect 288806 248376 288862 248432
rect 288990 248376 289046 248432
rect 288806 180784 288862 180840
rect 288990 180784 289046 180840
rect 288898 44104 288954 44160
rect 289082 44104 289138 44160
rect 289266 16788 289322 16824
rect 289266 16768 289268 16788
rect 289268 16768 289320 16788
rect 289320 16768 289322 16788
rect 290002 284280 290058 284336
rect 290278 284280 290334 284336
rect 290002 172624 290058 172680
rect 290002 172488 290058 172544
rect 290094 102040 290150 102096
rect 289910 101904 289966 101960
rect 289910 16496 289966 16552
rect 291474 172624 291530 172680
rect 291474 172488 291530 172544
rect 295246 296656 295302 296712
rect 294142 267688 294198 267744
rect 294418 267688 294474 267744
rect 294234 258052 294290 258088
rect 294234 258032 294236 258052
rect 294236 258032 294288 258052
rect 294288 258032 294290 258052
rect 294418 258032 294474 258088
rect 295246 157936 295302 157992
rect 295246 157528 295302 157584
rect 294142 27648 294198 27704
rect 294142 27512 294198 27568
rect 295522 296656 295578 296712
rect 296534 76200 296590 76256
rect 296534 75792 296590 75848
rect 296902 248376 296958 248432
rect 297178 248376 297234 248432
rect 296810 93744 296866 93800
rect 297178 93608 297234 93664
rect 297546 87100 297602 87136
rect 297546 87080 297548 87100
rect 297548 87080 297600 87100
rect 297600 87080 297602 87100
rect 298006 157548 298062 157584
rect 298006 157528 298008 157548
rect 298008 157528 298060 157548
rect 298060 157528 298062 157548
rect 298006 29416 298062 29472
rect 298006 29144 298062 29200
rect 298098 16532 298100 16552
rect 298100 16532 298152 16552
rect 298152 16532 298154 16552
rect 298098 16496 298154 16532
rect 298466 17040 298522 17096
rect 299662 277344 299718 277400
rect 299938 277344 299994 277400
rect 301134 325624 301190 325680
rect 301318 325624 301374 325680
rect 301226 306312 301282 306368
rect 301410 306312 301466 306368
rect 301042 296692 301044 296712
rect 301044 296692 301096 296712
rect 301096 296692 301098 296712
rect 301042 296656 301098 296692
rect 301134 296520 301190 296576
rect 301042 241440 301098 241496
rect 301134 241304 301190 241360
rect 301042 222128 301098 222184
rect 301134 221992 301190 222048
rect 301042 202816 301098 202872
rect 301134 202680 301190 202736
rect 301042 164192 301098 164248
rect 301226 164192 301282 164248
rect 301042 144880 301098 144936
rect 301226 144880 301282 144936
rect 301042 125568 301098 125624
rect 301226 125568 301282 125624
rect 302422 249736 302478 249792
rect 302606 249736 302662 249792
rect 302606 162852 302662 162888
rect 302606 162832 302608 162852
rect 302608 162832 302660 162852
rect 302660 162832 302662 162852
rect 302790 162832 302846 162888
rect 302606 143540 302662 143576
rect 302606 143520 302608 143540
rect 302608 143520 302660 143540
rect 302660 143520 302662 143540
rect 302790 143520 302846 143576
rect 302790 29008 302846 29064
rect 302790 28736 302846 28792
rect 306286 157392 306342 157448
rect 306286 86944 306342 87000
rect 306378 75948 306434 75984
rect 306378 75928 306380 75948
rect 306380 75928 306432 75948
rect 306432 75928 306434 75948
rect 306378 40180 306434 40216
rect 306378 40160 306380 40180
rect 306380 40160 306432 40180
rect 306432 40160 306434 40180
rect 306378 28772 306380 28792
rect 306380 28772 306432 28792
rect 306432 28772 306434 28792
rect 306378 28736 306434 28772
rect 306378 17060 306434 17096
rect 306378 17040 306380 17060
rect 306380 17040 306432 17060
rect 306432 17040 306434 17060
rect 307758 337592 307814 337648
rect 306746 287000 306802 287056
rect 307022 287000 307078 287056
rect 306930 249772 306932 249792
rect 306932 249772 306984 249792
rect 306984 249772 306986 249792
rect 306930 249736 306986 249772
rect 307114 249736 307170 249792
rect 306838 162852 306894 162888
rect 306838 162832 306840 162852
rect 306840 162832 306892 162852
rect 306892 162832 306894 162852
rect 307022 162832 307078 162888
rect 307574 157428 307576 157448
rect 307576 157428 307628 157448
rect 307628 157428 307630 157448
rect 307574 157392 307630 157428
rect 307574 16496 307630 16552
rect 307390 3304 307446 3360
rect 310794 193160 310850 193216
rect 311070 193160 311126 193216
rect 310886 153312 310942 153368
rect 310794 153196 310850 153232
rect 310794 153176 310796 153196
rect 310796 153176 310848 153196
rect 310848 153176 310850 153196
rect 311254 75948 311310 75984
rect 311254 75928 311256 75948
rect 311256 75928 311308 75948
rect 311308 75928 311310 75948
rect 310794 16496 310850 16552
rect 315946 157428 315948 157448
rect 315948 157428 316000 157448
rect 316000 157428 316002 157448
rect 315946 157392 316002 157428
rect 315946 40024 316002 40080
rect 315946 28872 316002 28928
rect 315946 16632 316002 16688
rect 314658 4800 314714 4856
rect 317326 337592 317382 337648
rect 317326 157664 317382 157720
rect 317326 157392 317382 157448
rect 317326 29280 317382 29336
rect 317326 28872 317382 28928
rect 323306 211112 323362 211168
rect 323490 211112 323546 211168
rect 323306 193196 323308 193216
rect 323308 193196 323360 193216
rect 323360 193196 323362 193216
rect 323306 193160 323362 193196
rect 323490 193196 323492 193216
rect 323492 193196 323544 193216
rect 323544 193196 323546 193216
rect 323490 193160 323546 193196
rect 324594 182144 324650 182200
rect 324870 182144 324926 182200
rect 325882 249772 325884 249792
rect 325884 249772 325936 249792
rect 325936 249772 325938 249792
rect 325882 249736 325938 249772
rect 326158 249736 326214 249792
rect 325882 202852 325884 202872
rect 325884 202852 325936 202872
rect 325936 202852 325938 202872
rect 325882 202816 325938 202852
rect 325974 202680 326030 202736
rect 325882 144900 325938 144936
rect 325882 144880 325884 144900
rect 325884 144880 325936 144900
rect 325936 144880 325938 144900
rect 326066 144900 326122 144936
rect 326066 144880 326068 144900
rect 326068 144880 326120 144900
rect 326120 144880 326122 144900
rect 327170 288396 327172 288416
rect 327172 288396 327224 288416
rect 327224 288396 327226 288416
rect 327170 288360 327226 288396
rect 327538 288360 327594 288416
rect 327170 230424 327226 230480
rect 327538 230424 327594 230480
rect 327262 212472 327318 212528
rect 327354 212336 327410 212392
rect 327170 183504 327226 183560
rect 327354 183504 327410 183560
rect 327262 172488 327318 172544
rect 327538 172488 327594 172544
rect 327262 153176 327318 153232
rect 327446 153176 327502 153232
rect 327170 144900 327226 144936
rect 327170 144880 327172 144900
rect 327172 144880 327224 144900
rect 327224 144880 327226 144900
rect 327354 144880 327410 144936
rect 327170 125588 327226 125624
rect 327170 125568 327172 125588
rect 327172 125568 327224 125588
rect 327224 125568 327226 125588
rect 327354 125568 327410 125624
rect 328274 110744 328330 110800
rect 328458 110744 328514 110800
rect 329930 219408 329986 219464
rect 329930 172488 329986 172544
rect 330206 315968 330262 316024
rect 330390 315968 330446 316024
rect 330206 298016 330262 298072
rect 330390 298016 330446 298072
rect 330206 248376 330262 248432
rect 330390 248376 330446 248432
rect 330206 229064 330262 229120
rect 330390 229064 330446 229120
rect 330114 219428 330170 219464
rect 330114 219408 330116 219428
rect 330116 219408 330168 219428
rect 330168 219408 330170 219428
rect 330114 183504 330170 183560
rect 330114 183368 330170 183424
rect 330206 172488 330262 172544
rect 330482 157936 330538 157992
rect 330482 157664 330538 157720
rect 330482 29280 330538 29336
rect 330482 29008 330538 29064
rect 330114 28872 330170 28928
rect 330206 28736 330262 28792
rect 336738 249872 336794 249928
rect 336738 183504 336794 183560
rect 336646 17040 336702 17096
rect 336646 16632 336702 16688
rect 337106 249872 337162 249928
rect 337106 249736 337162 249792
rect 337290 249736 337346 249792
rect 337198 230424 337254 230480
rect 337382 230424 337438 230480
rect 337106 202816 337162 202872
rect 337382 202816 337438 202872
rect 336922 183504 336978 183560
rect 337198 66136 337254 66192
rect 337290 56616 337346 56672
rect 339498 172488 339554 172544
rect 339866 172488 339922 172544
rect 339682 144880 339738 144936
rect 339866 144880 339922 144936
rect 340878 125568 340934 125624
rect 341246 299376 341302 299432
rect 341246 289856 341302 289912
rect 341246 280064 341302 280120
rect 341246 270544 341302 270600
rect 341246 260752 341302 260808
rect 341246 251232 341302 251288
rect 341154 240080 341210 240136
rect 341430 240080 341486 240136
rect 341154 202852 341156 202872
rect 341156 202852 341208 202872
rect 341208 202852 341210 202872
rect 341154 202816 341210 202852
rect 341430 202816 341486 202872
rect 341062 144880 341118 144936
rect 341246 144880 341302 144936
rect 341246 135244 341302 135280
rect 341246 135224 341248 135244
rect 341248 135224 341300 135244
rect 341300 135224 341302 135244
rect 341430 135224 341486 135280
rect 341062 125588 341118 125624
rect 341062 125568 341064 125588
rect 341064 125568 341116 125588
rect 341116 125568 341118 125588
rect 341246 106256 341302 106312
rect 341430 106256 341486 106312
rect 341246 48456 341302 48512
rect 341430 48320 341486 48376
rect 342718 337492 342720 337512
rect 342720 337492 342772 337512
rect 342772 337492 342774 337512
rect 342718 337456 342774 337492
rect 345754 337456 345810 337512
rect 346306 87080 346362 87136
rect 346306 86944 346362 87000
rect 347778 110508 347780 110528
rect 347780 110508 347832 110528
rect 347832 110508 347834 110528
rect 347778 110472 347834 110508
rect 347778 86980 347780 87000
rect 347780 86980 347832 87000
rect 347832 86980 347834 87000
rect 347778 86944 347834 86980
rect 347778 29044 347780 29064
rect 347780 29044 347832 29064
rect 347832 29044 347834 29064
rect 347778 29008 347834 29044
rect 347778 16924 347834 16960
rect 347778 16904 347780 16924
rect 347780 16904 347832 16924
rect 347832 16904 347834 16924
rect 352654 16632 352710 16688
rect 356242 3304 356298 3360
rect 357438 325624 357494 325680
rect 357622 325624 357678 325680
rect 357438 287000 357494 287056
rect 357806 287000 357862 287056
rect 357530 182144 357586 182200
rect 357714 182144 357770 182200
rect 357346 110744 357402 110800
rect 357346 87216 357402 87272
rect 357346 29280 357402 29336
rect 358542 316104 358598 316160
rect 358542 315968 358598 316024
rect 358726 261160 358782 261216
rect 358726 260888 358782 260944
rect 358542 259392 358598 259448
rect 358726 259392 358782 259448
rect 358542 240080 358598 240136
rect 358726 240080 358782 240136
rect 358542 220768 358598 220824
rect 358726 220768 358782 220824
rect 358542 172488 358598 172544
rect 358726 172488 358782 172544
rect 358634 85584 358690 85640
rect 359002 182144 359058 182200
rect 359186 182144 359242 182200
rect 359002 85312 359058 85368
rect 360474 182416 360530 182472
rect 360290 182144 360346 182200
rect 360474 95240 360530 95296
rect 360382 95104 360438 95160
rect 362038 306312 362094 306368
rect 362406 306312 362462 306368
rect 362314 133864 362370 133920
rect 362498 133864 362554 133920
rect 366822 241440 366878 241496
rect 366822 202816 366878 202872
rect 366822 106256 366878 106312
rect 367006 241476 367008 241496
rect 367008 241476 367060 241496
rect 367060 241476 367062 241496
rect 367006 241440 367062 241476
rect 367006 202816 367062 202872
rect 367006 106256 367062 106312
rect 367006 96872 367062 96928
rect 367006 96620 367062 96656
rect 367006 96600 367008 96620
rect 367008 96600 367060 96620
rect 367060 96600 367062 96620
rect 367098 76064 367154 76120
rect 367098 29144 367154 29200
rect 367098 29008 367154 29064
rect 368202 110472 368258 110528
rect 372526 241440 372582 241496
rect 372710 241440 372766 241496
rect 372526 222128 372582 222184
rect 372710 222128 372766 222184
rect 372526 202816 372582 202872
rect 372710 202816 372766 202872
rect 372802 173848 372858 173904
rect 372986 173848 373042 173904
rect 372802 164212 372858 164248
rect 372802 164192 372804 164212
rect 372804 164192 372856 164212
rect 372856 164192 372858 164212
rect 372986 164192 373042 164248
rect 376942 241440 376998 241496
rect 377126 241440 377182 241496
rect 376942 222128 376998 222184
rect 377126 222128 377182 222184
rect 376942 202816 376998 202872
rect 377126 202816 377182 202872
rect 376942 183504 376998 183560
rect 377126 183504 377182 183560
rect 376942 154536 376998 154592
rect 377126 154536 377182 154592
rect 376942 135224 376998 135280
rect 377126 135224 377182 135280
rect 376666 110744 376722 110800
rect 376758 87100 376814 87136
rect 376758 87080 376760 87100
rect 376760 87080 376812 87100
rect 376812 87080 376814 87100
rect 376666 76220 376722 76256
rect 376666 76200 376668 76220
rect 376668 76200 376720 76220
rect 376720 76200 376722 76220
rect 377126 29008 377182 29064
rect 377310 29008 377366 29064
rect 385130 16804 385132 16824
rect 385132 16804 385184 16824
rect 385184 16804 385186 16824
rect 385130 16768 385186 16804
rect 386234 86944 386290 87000
rect 386418 86944 386474 87000
rect 386418 76472 386474 76528
rect 386418 76200 386474 76256
rect 388994 251096 389050 251152
rect 388994 48184 389050 48240
rect 389178 251096 389234 251152
rect 389270 231784 389326 231840
rect 389454 231784 389510 231840
rect 389270 212472 389326 212528
rect 389454 212472 389510 212528
rect 389270 193160 389326 193216
rect 389454 193160 389510 193216
rect 389362 144880 389418 144936
rect 389638 144880 389694 144936
rect 389270 118768 389326 118824
rect 389454 108840 389510 108896
rect 389178 48184 389234 48240
rect 395986 87080 396042 87136
rect 396078 76084 396134 76120
rect 396078 76064 396080 76084
rect 396080 76064 396132 76084
rect 396132 76064 396134 76084
rect 396078 40196 396080 40216
rect 396080 40196 396132 40216
rect 396132 40196 396134 40216
rect 396078 40160 396134 40196
rect 395894 17040 395950 17096
rect 399390 76084 399446 76120
rect 399390 76064 399392 76084
rect 399392 76064 399444 76084
rect 399444 76064 399446 76084
rect 399022 40196 399024 40216
rect 399024 40196 399076 40216
rect 399076 40196 399078 40216
rect 399022 40160 399078 40196
rect 398746 16632 398802 16688
rect 398930 16632 398986 16688
rect 414018 110628 414074 110664
rect 414018 110608 414020 110628
rect 414020 110608 414072 110628
rect 414072 110608 414074 110628
rect 414018 63724 414020 63744
rect 414020 63724 414072 63744
rect 414072 63724 414074 63744
rect 414018 63688 414074 63724
rect 417882 157564 417884 157584
rect 417884 157564 417936 157584
rect 417936 157564 417938 157584
rect 417882 157528 417938 157564
rect 417882 40180 417938 40216
rect 417882 40160 417884 40180
rect 417884 40160 417936 40180
rect 417936 40160 417938 40180
rect 417882 16804 417884 16824
rect 417884 16804 417936 16824
rect 417936 16804 417938 16824
rect 417882 16768 417938 16804
rect 418250 157564 418252 157584
rect 418252 157564 418304 157584
rect 418304 157564 418306 157584
rect 418250 157528 418306 157564
rect 418894 63724 418896 63744
rect 418896 63724 418948 63744
rect 418948 63724 418950 63744
rect 418894 63688 418950 63724
rect 418250 40180 418306 40216
rect 418250 40160 418252 40180
rect 418252 40160 418304 40180
rect 418304 40160 418306 40180
rect 418250 16804 418252 16824
rect 418252 16804 418304 16824
rect 418304 16804 418306 16824
rect 418250 16768 418306 16804
rect 421194 278704 421250 278760
rect 421378 278704 421434 278760
rect 421194 259392 421250 259448
rect 421378 259392 421434 259448
rect 421194 241712 421250 241768
rect 421194 241576 421250 241632
rect 421194 240080 421250 240136
rect 421378 240080 421434 240136
rect 421194 220768 421250 220824
rect 421378 220768 421434 220824
rect 421102 196560 421158 196616
rect 421194 183640 421250 183696
rect 421194 172488 421250 172544
rect 421378 172488 421434 172544
rect 421010 67632 421066 67688
rect 421194 67632 421250 67688
rect 423494 110472 423550 110528
rect 421378 3440 421434 3496
rect 421562 3440 421618 3496
rect 424598 212472 424654 212528
rect 424782 212472 424838 212528
rect 437202 157548 437258 157584
rect 437202 157528 437204 157548
rect 437204 157528 437256 157548
rect 437256 157528 437258 157548
rect 437202 110628 437258 110664
rect 437202 110608 437204 110628
rect 437204 110608 437256 110628
rect 437256 110608 437258 110628
rect 437202 87116 437204 87136
rect 437204 87116 437256 87136
rect 437256 87116 437258 87136
rect 437202 87080 437258 87116
rect 437202 76084 437258 76120
rect 437202 76064 437204 76084
rect 437204 76064 437256 76084
rect 437256 76064 437258 76084
rect 437202 63708 437258 63744
rect 437202 63688 437204 63708
rect 437204 63688 437256 63708
rect 437256 63688 437258 63708
rect 437202 40196 437204 40216
rect 437204 40196 437256 40216
rect 437256 40196 437258 40216
rect 437202 40160 437258 40196
rect 437202 29164 437258 29200
rect 437202 29144 437204 29164
rect 437204 29144 437256 29164
rect 437256 29144 437258 29164
rect 437202 16788 437258 16824
rect 437202 16768 437204 16788
rect 437204 16768 437256 16788
rect 437256 16768 437258 16788
rect 437478 157548 437534 157584
rect 437478 157528 437480 157548
rect 437480 157528 437532 157548
rect 437532 157528 437534 157548
rect 437478 110628 437534 110664
rect 437478 110608 437480 110628
rect 437480 110608 437532 110628
rect 437532 110608 437534 110628
rect 437478 87116 437480 87136
rect 437480 87116 437532 87136
rect 437532 87116 437534 87136
rect 437478 87080 437534 87116
rect 437478 76084 437534 76120
rect 437478 76064 437480 76084
rect 437480 76064 437532 76084
rect 437532 76064 437534 76084
rect 437478 63708 437534 63744
rect 437478 63688 437480 63708
rect 437480 63688 437532 63708
rect 437532 63688 437534 63708
rect 437478 40196 437480 40216
rect 437480 40196 437532 40216
rect 437532 40196 437534 40216
rect 437478 40160 437534 40196
rect 437478 29164 437534 29200
rect 437478 29144 437480 29164
rect 437480 29144 437532 29164
rect 437532 29144 437534 29164
rect 437478 16788 437534 16824
rect 437478 16768 437480 16788
rect 437480 16768 437532 16788
rect 437532 16768 437534 16788
rect 456522 157548 456578 157584
rect 456522 157528 456524 157548
rect 456524 157528 456576 157548
rect 456576 157528 456578 157548
rect 456522 110644 456524 110664
rect 456524 110644 456576 110664
rect 456576 110644 456578 110664
rect 456522 110608 456578 110644
rect 456522 87116 456524 87136
rect 456524 87116 456576 87136
rect 456576 87116 456578 87136
rect 456522 87080 456578 87116
rect 456522 76084 456578 76120
rect 456522 76064 456524 76084
rect 456524 76064 456576 76084
rect 456576 76064 456578 76084
rect 456522 63708 456578 63744
rect 456522 63688 456524 63708
rect 456524 63688 456576 63708
rect 456576 63688 456578 63708
rect 456522 40180 456578 40216
rect 456522 40160 456524 40180
rect 456524 40160 456576 40180
rect 456576 40160 456578 40180
rect 456522 29180 456524 29200
rect 456524 29180 456576 29200
rect 456576 29180 456578 29200
rect 456522 29144 456578 29180
rect 456522 16804 456524 16824
rect 456524 16804 456576 16824
rect 456576 16804 456578 16824
rect 456522 16768 456578 16804
rect 456890 157548 456946 157584
rect 456890 157528 456892 157548
rect 456892 157528 456944 157548
rect 456944 157528 456946 157548
rect 456982 87116 456984 87136
rect 456984 87116 457036 87136
rect 457036 87116 457038 87136
rect 456982 87080 457038 87116
rect 456798 76084 456854 76120
rect 456798 76064 456800 76084
rect 456800 76064 456852 76084
rect 456852 76064 456854 76084
rect 456890 63708 456946 63744
rect 456890 63688 456892 63708
rect 456892 63688 456944 63708
rect 456944 63688 456946 63708
rect 456890 40180 456946 40216
rect 456890 40160 456892 40180
rect 456892 40160 456944 40180
rect 456944 40160 456946 40180
rect 456982 29180 456984 29200
rect 456984 29180 457036 29200
rect 457036 29180 457038 29200
rect 456982 29144 457038 29180
rect 458822 110644 458824 110664
rect 458824 110644 458876 110664
rect 458876 110644 458878 110664
rect 458822 110608 458878 110644
rect 458822 16804 458824 16824
rect 458824 16804 458876 16824
rect 458876 16804 458878 16824
rect 458822 16768 458878 16804
rect 460110 3748 460112 3768
rect 460112 3748 460164 3768
rect 460164 3748 460166 3768
rect 460110 3712 460166 3748
rect 463514 3712 463570 3768
rect 463790 231784 463846 231840
rect 463974 231784 464030 231840
rect 463790 212472 463846 212528
rect 463974 212472 464030 212528
rect 463790 193160 463846 193216
rect 463974 193160 464030 193216
rect 463882 154536 463938 154592
rect 464066 154536 464122 154592
rect 463882 125568 463938 125624
rect 464066 125568 464122 125624
rect 467562 337320 467618 337376
rect 467746 4800 467802 4856
rect 468758 3304 468814 3360
rect 580170 580760 580226 580816
rect 579710 557232 579766 557288
rect 579710 545536 579766 545592
rect 579710 510312 579766 510368
rect 579710 498616 579766 498672
rect 579710 463392 579766 463448
rect 579802 451696 579858 451752
rect 579802 439864 579858 439920
rect 579802 416472 579858 416528
rect 579802 404776 579858 404832
rect 579802 392944 579858 393000
rect 579894 369552 579950 369608
rect 579986 357856 580042 357912
rect 579986 346024 580042 346080
rect 470506 337184 470562 337240
rect 470690 337184 470746 337240
rect 470414 231784 470470 231840
rect 470598 231784 470654 231840
rect 470414 212472 470470 212528
rect 470598 212472 470654 212528
rect 470414 193160 470470 193216
rect 470598 193160 470654 193216
rect 470414 173848 470470 173904
rect 470598 173848 470654 173904
rect 470414 164192 470470 164248
rect 470598 164192 470654 164248
rect 470414 144880 470470 144936
rect 470598 144880 470654 144936
rect 470414 125568 470470 125624
rect 470598 125568 470654 125624
rect 476026 87216 476082 87272
rect 476210 87080 476266 87136
rect 476026 29280 476082 29336
rect 476210 29144 476266 29200
rect 482926 111016 482982 111072
rect 482926 110608 482982 110664
rect 482926 76472 482982 76528
rect 482926 76064 482982 76120
rect 482926 17176 482982 17232
rect 482926 16768 482982 16824
rect 487802 110880 487858 110936
rect 487802 110472 487858 110528
rect 491206 87352 491262 87408
rect 491206 86944 491262 87000
rect 487802 76336 487858 76392
rect 487802 75928 487858 75984
rect 491206 29416 491262 29472
rect 491206 29008 491262 29064
rect 487802 17040 487858 17096
rect 487802 16632 487858 16688
rect 494610 86944 494666 87000
rect 492770 29044 492772 29064
rect 492772 29044 492824 29064
rect 492824 29044 492826 29064
rect 492770 29008 492826 29044
rect 502246 87216 502302 87272
rect 502246 29280 502302 29336
rect 512642 337320 512698 337376
rect 579986 322632 580042 322688
rect 580078 310800 580134 310856
rect 579802 299104 579858 299160
rect 580170 275712 580226 275768
rect 580170 252184 580226 252240
rect 580906 263880 580962 263936
rect 580814 228792 580870 228848
rect 580722 216960 580778 217016
rect 580630 205264 580686 205320
rect 580538 181872 580594 181928
rect 580446 170040 580502 170096
rect 580354 134816 580410 134872
rect 580262 123120 580318 123176
rect 576214 4800 576270 4856
rect 580998 3304 581054 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 378133 700362 378199 700365
rect 8109 700360 378199 700362
rect 8109 700304 8114 700360
rect 8170 700304 378138 700360
rect 378194 700304 378199 700360
rect 8109 700302 378199 700304
rect 8109 700299 8175 700302
rect 378133 700299 378199 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect 4797 583538 4863 583541
rect 460289 583538 460355 583541
rect 4797 583536 460355 583538
rect 4797 583480 4802 583536
rect 4858 583480 460294 583536
rect 460350 583480 460355 583536
rect 4797 583478 460355 583480
rect 4797 583475 4863 583478
rect 460289 583475 460355 583478
rect 300301 583402 300367 583405
rect 465942 583402 465948 583404
rect 300301 583400 465948 583402
rect 300301 583344 300306 583400
rect 300362 583344 465948 583400
rect 300301 583342 465948 583344
rect 300301 583339 300367 583342
rect 465942 583340 465948 583342
rect 466012 583340 466018 583404
rect 293953 583266 294019 583269
rect 465758 583266 465764 583268
rect 293953 583264 465764 583266
rect 293953 583208 293958 583264
rect 294014 583208 465764 583264
rect 293953 583206 465764 583208
rect 293953 583203 294019 583206
rect 465758 583204 465764 583206
rect 465828 583204 465834 583268
rect 242750 583068 242756 583132
rect 242820 583130 242826 583132
rect 420269 583130 420335 583133
rect 242820 583128 420335 583130
rect 242820 583072 420274 583128
rect 420330 583072 420335 583128
rect 242820 583070 420335 583072
rect 242820 583068 242826 583070
rect 420269 583067 420335 583070
rect 239254 582932 239260 582996
rect 239324 582994 239330 582996
rect 426617 582994 426683 582997
rect 239324 582992 426683 582994
rect 239324 582936 426622 582992
rect 426678 582936 426683 582992
rect 239324 582934 426683 582936
rect 239324 582932 239330 582934
rect 426617 582931 426683 582934
rect 17217 582858 17283 582861
rect 449801 582858 449867 582861
rect 17217 582856 449867 582858
rect 17217 582800 17222 582856
rect 17278 582800 449806 582856
rect 449862 582800 449867 582856
rect 17217 582798 449867 582800
rect 17217 582795 17283 582798
rect 449801 582795 449867 582798
rect 24117 582722 24183 582725
rect 462405 582722 462471 582725
rect 24117 582720 462471 582722
rect 24117 582664 24122 582720
rect 24178 582664 462410 582720
rect 462466 582664 462471 582720
rect 24117 582662 462471 582664
rect 24117 582659 24183 582662
rect 462405 582659 462471 582662
rect 5073 582586 5139 582589
rect 447685 582586 447751 582589
rect 5073 582584 447751 582586
rect 5073 582528 5078 582584
rect 5134 582528 447690 582584
rect 447746 582528 447751 582584
rect 5073 582526 447751 582528
rect 5073 582523 5139 582526
rect 447685 582523 447751 582526
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 465574 579668 465580 579732
rect 465644 579730 465650 579732
rect 468477 579730 468543 579733
rect 465644 579728 468543 579730
rect 465644 579672 468482 579728
rect 468538 579672 468543 579728
rect 465644 579670 468543 579672
rect 465644 579668 465650 579670
rect 468477 579667 468543 579670
rect 231117 579322 231183 579325
rect 232957 579324 233023 579325
rect 231710 579322 231716 579324
rect 231117 579320 231716 579322
rect 231117 579264 231122 579320
rect 231178 579264 231716 579320
rect 231117 579262 231716 579264
rect 231117 579259 231183 579262
rect 231710 579260 231716 579262
rect 231780 579260 231786 579324
rect 232957 579320 233004 579324
rect 233068 579322 233074 579324
rect 235257 579322 235323 579325
rect 237189 579324 237255 579325
rect 235758 579322 235764 579324
rect 232957 579264 232962 579320
rect 232957 579260 233004 579264
rect 233068 579262 233114 579322
rect 235257 579320 235764 579322
rect 235257 579264 235262 579320
rect 235318 579264 235764 579320
rect 235257 579262 235764 579264
rect 233068 579260 233074 579262
rect 232957 579259 233023 579260
rect 235257 579259 235323 579262
rect 235758 579260 235764 579262
rect 235828 579260 235834 579324
rect 237189 579320 237236 579324
rect 237300 579322 237306 579324
rect 239397 579322 239463 579325
rect 239990 579322 239996 579324
rect 237189 579264 237194 579320
rect 237189 579260 237236 579264
rect 237300 579262 237346 579322
rect 239397 579320 239996 579322
rect 239397 579264 239402 579320
rect 239458 579264 239996 579320
rect 239397 579262 239996 579264
rect 237300 579260 237306 579262
rect 237189 579259 237255 579260
rect 239397 579259 239463 579262
rect 239990 579260 239996 579262
rect 240060 579260 240066 579324
rect 241278 579260 241284 579324
rect 241348 579322 241354 579324
rect 241421 579322 241487 579325
rect 241348 579320 241487 579322
rect 241348 579264 241426 579320
rect 241482 579264 241487 579320
rect 241348 579262 241487 579264
rect 241348 579260 241354 579262
rect 241421 579259 241487 579262
rect 243629 579322 243695 579325
rect 249517 579324 249583 579325
rect 466453 579324 466519 579325
rect 244038 579322 244044 579324
rect 243629 579320 244044 579322
rect 243629 579264 243634 579320
rect 243690 579264 244044 579320
rect 243629 579262 244044 579264
rect 243629 579259 243695 579262
rect 244038 579260 244044 579262
rect 244108 579260 244114 579324
rect 249517 579320 249564 579324
rect 249628 579322 249634 579324
rect 249517 579264 249522 579320
rect 249517 579260 249564 579264
rect 249628 579262 249674 579322
rect 466453 579320 466500 579324
rect 466564 579322 466570 579324
rect 466453 579264 466458 579320
rect 249628 579260 249634 579262
rect 466453 579260 466500 579264
rect 466564 579262 466610 579322
rect 466564 579260 466570 579262
rect 249517 579259 249583 579260
rect 466453 579259 466519 579260
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3049 567354 3115 567357
rect -960 567352 3115 567354
rect -960 567296 3054 567352
rect 3110 567296 3115 567352
rect -960 567294 3115 567296
rect -960 567204 480 567294
rect 3049 567291 3115 567294
rect 579705 557290 579771 557293
rect 583520 557290 584960 557380
rect 579705 557288 584960 557290
rect 579705 557232 579710 557288
rect 579766 557232 584960 557288
rect 579705 557230 584960 557232
rect 579705 557227 579771 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 2773 553074 2839 553077
rect -960 553072 2839 553074
rect -960 553016 2778 553072
rect 2834 553016 2839 553072
rect -960 553014 2839 553016
rect -960 552924 480 553014
rect 2773 553011 2839 553014
rect 579705 545594 579771 545597
rect 583520 545594 584960 545684
rect 579705 545592 584960 545594
rect 579705 545536 579710 545592
rect 579766 545536 584960 545592
rect 579705 545534 584960 545536
rect 579705 545531 579771 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3049 538658 3115 538661
rect -960 538656 3115 538658
rect -960 538600 3054 538656
rect 3110 538600 3115 538656
rect -960 538598 3115 538600
rect -960 538508 480 538598
rect 3049 538595 3115 538598
rect 583520 533898 584960 533988
rect 583342 533838 584960 533898
rect 465942 533020 465948 533084
rect 466012 533082 466018 533084
rect 466012 533022 470610 533082
rect 466012 533020 466018 533022
rect 470550 532946 470610 533022
rect 480302 533022 489930 533082
rect 470550 532886 480178 532946
rect 480118 532810 480178 532886
rect 480302 532810 480362 533022
rect 489870 532946 489930 533022
rect 499622 533022 509250 533082
rect 489870 532886 499498 532946
rect 480118 532750 480362 532810
rect 499438 532810 499498 532886
rect 499622 532810 499682 533022
rect 509190 532946 509250 533022
rect 518942 533022 528570 533082
rect 509190 532886 518818 532946
rect 499438 532750 499682 532810
rect 518758 532810 518818 532886
rect 518942 532810 519002 533022
rect 528510 532946 528570 533022
rect 538262 533022 547890 533082
rect 528510 532886 538138 532946
rect 518758 532750 519002 532810
rect 538078 532810 538138 532886
rect 538262 532810 538322 533022
rect 547830 532946 547890 533022
rect 557582 533022 567210 533082
rect 547830 532886 557458 532946
rect 538078 532750 538322 532810
rect 557398 532810 557458 532886
rect 557582 532810 557642 533022
rect 567150 532946 567210 533022
rect 583342 532946 583402 533838
rect 583520 533748 584960 533838
rect 567150 532886 576778 532946
rect 557398 532750 557642 532810
rect 576718 532810 576778 532886
rect 576902 532886 583402 532946
rect 576902 532810 576962 532886
rect 576718 532750 576962 532810
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579705 510370 579771 510373
rect 583520 510370 584960 510460
rect 579705 510368 584960 510370
rect 579705 510312 579710 510368
rect 579766 510312 584960 510368
rect 579705 510310 584960 510312
rect 579705 510307 579771 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3049 509962 3115 509965
rect -960 509960 3115 509962
rect -960 509904 3054 509960
rect 3110 509904 3115 509960
rect -960 509902 3115 509904
rect -960 509812 480 509902
rect 3049 509899 3115 509902
rect 579705 498674 579771 498677
rect 583520 498674 584960 498764
rect 579705 498672 584960 498674
rect 579705 498616 579710 498672
rect 579766 498616 584960 498672
rect 579705 498614 584960 498616
rect 579705 498611 579771 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 583520 486842 584960 486932
rect 583342 486782 584960 486842
rect 465758 486100 465764 486164
rect 465828 486162 465834 486164
rect 465828 486102 470610 486162
rect 465828 486100 465834 486102
rect 470550 486026 470610 486102
rect 480302 486102 489930 486162
rect 470550 485966 480178 486026
rect 480118 485890 480178 485966
rect 480302 485890 480362 486102
rect 489870 486026 489930 486102
rect 499622 486102 509250 486162
rect 489870 485966 499498 486026
rect 480118 485830 480362 485890
rect 499438 485890 499498 485966
rect 499622 485890 499682 486102
rect 509190 486026 509250 486102
rect 518942 486102 528570 486162
rect 509190 485966 518818 486026
rect 499438 485830 499682 485890
rect 518758 485890 518818 485966
rect 518942 485890 519002 486102
rect 528510 486026 528570 486102
rect 538262 486102 547890 486162
rect 528510 485966 538138 486026
rect 518758 485830 519002 485890
rect 538078 485890 538138 485966
rect 538262 485890 538322 486102
rect 547830 486026 547890 486102
rect 557582 486102 567210 486162
rect 547830 485966 557458 486026
rect 538078 485830 538322 485890
rect 557398 485890 557458 485966
rect 557582 485890 557642 486102
rect 567150 486026 567210 486102
rect 583342 486026 583402 486782
rect 583520 486692 584960 486782
rect 567150 485966 576778 486026
rect 557398 485830 557642 485890
rect 576718 485890 576778 485966
rect 576902 485966 583402 486026
rect 576902 485890 576962 485966
rect 576718 485830 576962 485890
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579705 463450 579771 463453
rect 583520 463450 584960 463540
rect 579705 463448 584960 463450
rect 579705 463392 579710 463448
rect 579766 463392 584960 463448
rect 579705 463390 584960 463392
rect 579705 463387 579771 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3141 452434 3207 452437
rect -960 452432 3207 452434
rect -960 452376 3146 452432
rect 3202 452376 3207 452432
rect -960 452374 3207 452376
rect -960 452284 480 452374
rect 3141 452371 3207 452374
rect 579797 451754 579863 451757
rect 583520 451754 584960 451844
rect 579797 451752 584960 451754
rect 579797 451696 579802 451752
rect 579858 451696 584960 451752
rect 579797 451694 584960 451696
rect 579797 451691 579863 451694
rect 583520 451604 584960 451694
rect 579797 439922 579863 439925
rect 583520 439922 584960 440012
rect 579797 439920 584960 439922
rect 579797 439864 579802 439920
rect 579858 439864 584960 439920
rect 579797 439862 584960 439864
rect 579797 439859 579863 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3141 423738 3207 423741
rect -960 423736 3207 423738
rect -960 423680 3146 423736
rect 3202 423680 3207 423736
rect -960 423678 3207 423680
rect -960 423588 480 423678
rect 3141 423675 3207 423678
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579797 404834 579863 404837
rect 583520 404834 584960 404924
rect 579797 404832 584960 404834
rect 579797 404776 579802 404832
rect 579858 404776 584960 404832
rect 579797 404774 584960 404776
rect 579797 404771 579863 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3233 395042 3299 395045
rect -960 395040 3299 395042
rect -960 394984 3238 395040
rect 3294 394984 3299 395040
rect -960 394982 3299 394984
rect -960 394892 480 394982
rect 3233 394979 3299 394982
rect 579797 393002 579863 393005
rect 583520 393002 584960 393092
rect 579797 393000 584960 393002
rect 579797 392944 579802 393000
rect 579858 392944 584960 393000
rect 579797 392942 584960 392944
rect 579797 392939 579863 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 579889 369610 579955 369613
rect 583520 369610 584960 369700
rect 579889 369608 584960 369610
rect 579889 369552 579894 369608
rect 579950 369552 584960 369608
rect 579889 369550 584960 369552
rect 579889 369547 579955 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3325 366210 3391 366213
rect -960 366208 3391 366210
rect -960 366152 3330 366208
rect 3386 366152 3391 366208
rect -960 366150 3391 366152
rect -960 366060 480 366150
rect 3325 366147 3391 366150
rect 579981 357914 580047 357917
rect 583520 357914 584960 358004
rect 579981 357912 584960 357914
rect 579981 357856 579986 357912
rect 580042 357856 584960 357912
rect 579981 357854 584960 357856
rect 579981 357851 580047 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579981 346082 580047 346085
rect 583520 346082 584960 346172
rect 579981 346080 584960 346082
rect 579981 346024 579986 346080
rect 580042 346024 584960 346080
rect 579981 346022 584960 346024
rect 579981 346019 580047 346022
rect 583520 345932 584960 346022
rect 243670 340580 243676 340644
rect 243740 340642 243746 340644
rect 249558 340642 249564 340644
rect 243740 340582 249564 340642
rect 243740 340580 243746 340582
rect 249558 340580 249564 340582
rect 249628 340580 249634 340644
rect 242750 338058 242756 338060
rect 614 337998 242756 338058
rect -960 337514 480 337604
rect 614 337514 674 337998
rect 242750 337996 242756 337998
rect 242820 337996 242826 338060
rect 57973 337786 58039 337789
rect 67541 337786 67607 337789
rect 57973 337784 67607 337786
rect 57973 337728 57978 337784
rect 58034 337728 67546 337784
rect 67602 337728 67607 337784
rect 57973 337726 67607 337728
rect 57973 337723 58039 337726
rect 67541 337723 67607 337726
rect 77293 337786 77359 337789
rect 86861 337786 86927 337789
rect 77293 337784 86927 337786
rect 77293 337728 77298 337784
rect 77354 337728 86866 337784
rect 86922 337728 86927 337784
rect 77293 337726 86927 337728
rect 77293 337723 77359 337726
rect 86861 337723 86927 337726
rect 95233 337786 95299 337789
rect 104801 337786 104867 337789
rect 95233 337784 104867 337786
rect 95233 337728 95238 337784
rect 95294 337728 104806 337784
rect 104862 337728 104867 337784
rect 95233 337726 104867 337728
rect 95233 337723 95299 337726
rect 104801 337723 104867 337726
rect 114553 337786 114619 337789
rect 124121 337786 124187 337789
rect 114553 337784 124187 337786
rect 114553 337728 114558 337784
rect 114614 337728 124126 337784
rect 124182 337728 124187 337784
rect 114553 337726 124187 337728
rect 114553 337723 114619 337726
rect 124121 337723 124187 337726
rect 133873 337786 133939 337789
rect 143441 337786 143507 337789
rect 133873 337784 143507 337786
rect 133873 337728 133878 337784
rect 133934 337728 143446 337784
rect 143502 337728 143507 337784
rect 133873 337726 143507 337728
rect 133873 337723 133939 337726
rect 143441 337723 143507 337726
rect 153193 337786 153259 337789
rect 162761 337786 162827 337789
rect 153193 337784 162827 337786
rect 153193 337728 153198 337784
rect 153254 337728 162766 337784
rect 162822 337728 162827 337784
rect 153193 337726 162827 337728
rect 153193 337723 153259 337726
rect 162761 337723 162827 337726
rect 172513 337786 172579 337789
rect 182081 337786 182147 337789
rect 172513 337784 182147 337786
rect 172513 337728 172518 337784
rect 172574 337728 182086 337784
rect 182142 337728 182147 337784
rect 172513 337726 182147 337728
rect 172513 337723 172579 337726
rect 182081 337723 182147 337726
rect 191833 337786 191899 337789
rect 201401 337786 201467 337789
rect 191833 337784 201467 337786
rect 191833 337728 191838 337784
rect 191894 337728 201406 337784
rect 201462 337728 201467 337784
rect 191833 337726 201467 337728
rect 191833 337723 191899 337726
rect 201401 337723 201467 337726
rect 211153 337786 211219 337789
rect 220721 337786 220787 337789
rect 211153 337784 220787 337786
rect 211153 337728 211158 337784
rect 211214 337728 220726 337784
rect 220782 337728 220787 337784
rect 211153 337726 220787 337728
rect 211153 337723 211219 337726
rect 220721 337723 220787 337726
rect 307753 337650 307819 337653
rect 317321 337650 317387 337653
rect 307753 337648 317387 337650
rect 307753 337592 307758 337648
rect 307814 337592 317326 337648
rect 317382 337592 317387 337648
rect 307753 337590 317387 337592
rect 307753 337587 307819 337590
rect 317321 337587 317387 337590
rect -960 337454 674 337514
rect 342713 337514 342779 337517
rect 345749 337514 345815 337517
rect 342713 337512 345815 337514
rect 342713 337456 342718 337512
rect 342774 337456 345754 337512
rect 345810 337456 345815 337512
rect 342713 337454 345815 337456
rect -960 337364 480 337454
rect 342713 337451 342779 337454
rect 345749 337451 345815 337454
rect 10317 337378 10383 337381
rect 231945 337378 232011 337381
rect 10317 337376 232011 337378
rect 10317 337320 10322 337376
rect 10378 337320 231950 337376
rect 232006 337320 232011 337376
rect 10317 337318 232011 337320
rect 10317 337315 10383 337318
rect 231945 337315 232011 337318
rect 467557 337378 467623 337381
rect 512637 337378 512703 337381
rect 467557 337376 512703 337378
rect 467557 337320 467562 337376
rect 467618 337320 512642 337376
rect 512698 337320 512703 337376
rect 467557 337318 512703 337320
rect 467557 337315 467623 337318
rect 512637 337315 512703 337318
rect 132493 337242 132559 337245
rect 142061 337242 142127 337245
rect 132493 337240 142127 337242
rect 132493 337184 132498 337240
rect 132554 337184 142066 337240
rect 142122 337184 142127 337240
rect 132493 337182 142127 337184
rect 132493 337179 132559 337182
rect 142061 337179 142127 337182
rect 151813 337242 151879 337245
rect 161381 337242 161447 337245
rect 151813 337240 161447 337242
rect 151813 337184 151818 337240
rect 151874 337184 161386 337240
rect 161442 337184 161447 337240
rect 151813 337182 161447 337184
rect 151813 337179 151879 337182
rect 161381 337179 161447 337182
rect 171133 337242 171199 337245
rect 180701 337242 180767 337245
rect 171133 337240 180767 337242
rect 171133 337184 171138 337240
rect 171194 337184 180706 337240
rect 180762 337184 180767 337240
rect 171133 337182 180767 337184
rect 171133 337179 171199 337182
rect 180701 337179 180767 337182
rect 190453 337242 190519 337245
rect 200021 337242 200087 337245
rect 190453 337240 200087 337242
rect 190453 337184 190458 337240
rect 190514 337184 200026 337240
rect 200082 337184 200087 337240
rect 190453 337182 200087 337184
rect 190453 337179 190519 337182
rect 200021 337179 200087 337182
rect 209773 337242 209839 337245
rect 219341 337242 219407 337245
rect 209773 337240 219407 337242
rect 209773 337184 209778 337240
rect 209834 337184 219346 337240
rect 219402 337184 219407 337240
rect 209773 337182 219407 337184
rect 209773 337179 209839 337182
rect 219341 337179 219407 337182
rect 220997 337242 221063 337245
rect 234613 337242 234679 337245
rect 220997 337240 234679 337242
rect 220997 337184 221002 337240
rect 221058 337184 234618 337240
rect 234674 337184 234679 337240
rect 220997 337182 234679 337184
rect 220997 337179 221063 337182
rect 234613 337179 234679 337182
rect 470501 337242 470567 337245
rect 470685 337242 470751 337245
rect 470501 337240 470751 337242
rect 470501 337184 470506 337240
rect 470562 337184 470690 337240
rect 470746 337184 470751 337240
rect 470501 337182 470751 337184
rect 470501 337179 470567 337182
rect 470685 337179 470751 337182
rect 249241 336698 249307 336701
rect 249558 336698 249564 336700
rect 249241 336696 249564 336698
rect 249241 336640 249246 336696
rect 249302 336640 249564 336696
rect 249241 336638 249564 336640
rect 249241 336635 249307 336638
rect 249558 336636 249564 336638
rect 249628 336636 249634 336700
rect 583520 334236 584960 334476
rect 245929 325682 245995 325685
rect 246113 325682 246179 325685
rect 245929 325680 246179 325682
rect 245929 325624 245934 325680
rect 245990 325624 246118 325680
rect 246174 325624 246179 325680
rect 245929 325622 246179 325624
rect 245929 325619 245995 325622
rect 246113 325619 246179 325622
rect 301129 325682 301195 325685
rect 301313 325682 301379 325685
rect 301129 325680 301379 325682
rect 301129 325624 301134 325680
rect 301190 325624 301318 325680
rect 301374 325624 301379 325680
rect 301129 325622 301379 325624
rect 301129 325619 301195 325622
rect 301313 325619 301379 325622
rect 357433 325682 357499 325685
rect 357617 325682 357683 325685
rect 357433 325680 357683 325682
rect 357433 325624 357438 325680
rect 357494 325624 357622 325680
rect 357678 325624 357683 325680
rect 357433 325622 357683 325624
rect 357433 325619 357499 325622
rect 357617 325619 357683 325622
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 579981 322690 580047 322693
rect 583520 322690 584960 322780
rect 579981 322688 584960 322690
rect 579981 322632 579986 322688
rect 580042 322632 584960 322688
rect 579981 322630 584960 322632
rect 579981 322627 580047 322630
rect 583520 322540 584960 322630
rect 232221 318882 232287 318885
rect 232405 318882 232471 318885
rect 232221 318880 232471 318882
rect 232221 318824 232226 318880
rect 232282 318824 232410 318880
rect 232466 318824 232471 318880
rect 232221 318822 232471 318824
rect 232221 318819 232287 318822
rect 232405 318819 232471 318822
rect 249241 316298 249307 316301
rect 249198 316296 249307 316298
rect 249198 316240 249246 316296
rect 249302 316240 249307 316296
rect 249198 316235 249307 316240
rect 249198 316164 249258 316235
rect 249190 316100 249196 316164
rect 249260 316100 249266 316164
rect 358537 316162 358603 316165
rect 358537 316160 358738 316162
rect 358537 316104 358542 316160
rect 358598 316104 358738 316160
rect 358537 316102 358738 316104
rect 358537 316099 358603 316102
rect 245837 316026 245903 316029
rect 245702 316024 245903 316026
rect 245702 315968 245842 316024
rect 245898 315968 245903 316024
rect 245702 315966 245903 315968
rect 245702 315890 245762 315966
rect 245837 315963 245903 315966
rect 267825 316026 267891 316029
rect 268009 316026 268075 316029
rect 267825 316024 268075 316026
rect 267825 315968 267830 316024
rect 267886 315968 268014 316024
rect 268070 315968 268075 316024
rect 267825 315966 268075 315968
rect 267825 315963 267891 315966
rect 268009 315963 268075 315966
rect 273069 316026 273135 316029
rect 273253 316026 273319 316029
rect 273069 316024 273319 316026
rect 273069 315968 273074 316024
rect 273130 315968 273258 316024
rect 273314 315968 273319 316024
rect 273069 315966 273319 315968
rect 273069 315963 273135 315966
rect 273253 315963 273319 315966
rect 330201 316026 330267 316029
rect 330385 316026 330451 316029
rect 330201 316024 330451 316026
rect 330201 315968 330206 316024
rect 330262 315968 330390 316024
rect 330446 315968 330451 316024
rect 330201 315966 330451 315968
rect 330201 315963 330267 315966
rect 330385 315963 330451 315966
rect 358537 316026 358603 316029
rect 358678 316026 358738 316102
rect 358537 316024 358738 316026
rect 358537 315968 358542 316024
rect 358598 315968 358738 316024
rect 358537 315966 358738 315968
rect 358537 315963 358603 315966
rect 245929 315890 245995 315893
rect 245702 315888 245995 315890
rect 245702 315832 245934 315888
rect 245990 315832 245995 315888
rect 245702 315830 245995 315832
rect 245929 315827 245995 315830
rect 264973 314666 265039 314669
rect 265157 314666 265223 314669
rect 264973 314664 265223 314666
rect 264973 314608 264978 314664
rect 265034 314608 265162 314664
rect 265218 314608 265223 314664
rect 264973 314606 265223 314608
rect 264973 314603 265039 314606
rect 265157 314603 265223 314606
rect 249190 312020 249196 312084
rect 249260 312020 249266 312084
rect 249198 311810 249258 312020
rect 249374 311810 249380 311812
rect 249198 311750 249380 311810
rect 249374 311748 249380 311750
rect 249444 311748 249450 311812
rect 580073 310858 580139 310861
rect 583520 310858 584960 310948
rect 580073 310856 584960 310858
rect 580073 310800 580078 310856
rect 580134 310800 584960 310856
rect 580073 310798 584960 310800
rect 580073 310795 580139 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 2773 308818 2839 308821
rect -960 308816 2839 308818
rect -960 308760 2778 308816
rect 2834 308760 2839 308816
rect -960 308758 2839 308760
rect -960 308668 480 308758
rect 2773 308755 2839 308758
rect 251398 307668 251404 307732
rect 251468 307730 251474 307732
rect 251541 307730 251607 307733
rect 251468 307728 251607 307730
rect 251468 307672 251546 307728
rect 251602 307672 251607 307728
rect 251468 307670 251607 307672
rect 251468 307668 251474 307670
rect 251541 307667 251607 307670
rect 249241 306370 249307 306373
rect 249374 306370 249380 306372
rect 249241 306368 249380 306370
rect 249241 306312 249246 306368
rect 249302 306312 249380 306368
rect 249241 306310 249380 306312
rect 249241 306307 249307 306310
rect 249374 306308 249380 306310
rect 249444 306308 249450 306372
rect 259729 306370 259795 306373
rect 259913 306370 259979 306373
rect 259729 306368 259979 306370
rect 259729 306312 259734 306368
rect 259790 306312 259918 306368
rect 259974 306312 259979 306368
rect 259729 306310 259979 306312
rect 259729 306307 259795 306310
rect 259913 306307 259979 306310
rect 301221 306370 301287 306373
rect 301405 306370 301471 306373
rect 301221 306368 301471 306370
rect 301221 306312 301226 306368
rect 301282 306312 301410 306368
rect 301466 306312 301471 306368
rect 301221 306310 301471 306312
rect 301221 306307 301287 306310
rect 301405 306307 301471 306310
rect 362033 306370 362099 306373
rect 362401 306370 362467 306373
rect 362033 306368 362467 306370
rect 362033 306312 362038 306368
rect 362094 306312 362406 306368
rect 362462 306312 362467 306368
rect 362033 306310 362467 306312
rect 362033 306307 362099 306310
rect 362401 306307 362467 306310
rect 264973 305010 265039 305013
rect 265249 305010 265315 305013
rect 264973 305008 265315 305010
rect 264973 304952 264978 305008
rect 265034 304952 265254 305008
rect 265310 304952 265315 305008
rect 264973 304950 265315 304952
rect 264973 304947 265039 304950
rect 265249 304947 265315 304950
rect 341241 299434 341307 299437
rect 341374 299434 341380 299436
rect 341241 299432 341380 299434
rect 341241 299376 341246 299432
rect 341302 299376 341380 299432
rect 341241 299374 341380 299376
rect 341241 299371 341307 299374
rect 341374 299372 341380 299374
rect 341444 299372 341450 299436
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 251398 298148 251404 298212
rect 251468 298210 251474 298212
rect 251541 298210 251607 298213
rect 251468 298208 251607 298210
rect 251468 298152 251546 298208
rect 251602 298152 251607 298208
rect 251468 298150 251607 298152
rect 251468 298148 251474 298150
rect 251541 298147 251607 298150
rect 330201 298074 330267 298077
rect 330385 298074 330451 298077
rect 330201 298072 330451 298074
rect 330201 298016 330206 298072
rect 330262 298016 330390 298072
rect 330446 298016 330451 298072
rect 330201 298014 330451 298016
rect 330201 298011 330267 298014
rect 330385 298011 330451 298014
rect 249241 296986 249307 296989
rect 249198 296984 249307 296986
rect 249198 296928 249246 296984
rect 249302 296928 249307 296984
rect 249198 296923 249307 296928
rect 249198 296852 249258 296923
rect 249190 296788 249196 296852
rect 249260 296788 249266 296852
rect 295241 296714 295307 296717
rect 295517 296714 295583 296717
rect 301037 296714 301103 296717
rect 295241 296712 295583 296714
rect 295241 296656 295246 296712
rect 295302 296656 295522 296712
rect 295578 296656 295583 296712
rect 295241 296654 295583 296656
rect 295241 296651 295307 296654
rect 295517 296651 295583 296654
rect 300902 296712 301103 296714
rect 300902 296656 301042 296712
rect 301098 296656 301103 296712
rect 300902 296654 301103 296656
rect 300902 296578 300962 296654
rect 301037 296651 301103 296654
rect 301129 296578 301195 296581
rect 300902 296576 301195 296578
rect 300902 296520 301134 296576
rect 301190 296520 301195 296576
rect 300902 296518 301195 296520
rect 301129 296515 301195 296518
rect 259637 295354 259703 295357
rect 259913 295354 259979 295357
rect 259637 295352 259979 295354
rect 259637 295296 259642 295352
rect 259698 295296 259918 295352
rect 259974 295296 259979 295352
rect 259637 295294 259979 295296
rect 259637 295291 259703 295294
rect 259913 295291 259979 295294
rect 2957 295218 3023 295221
rect 239254 295218 239260 295220
rect 2957 295216 239260 295218
rect 2957 295160 2962 295216
rect 3018 295160 239260 295216
rect 2957 295158 239260 295160
rect 2957 295155 3023 295158
rect 239254 295156 239260 295158
rect 239324 295156 239330 295220
rect -960 294402 480 294492
rect 2957 294402 3023 294405
rect -960 294400 3023 294402
rect -960 294344 2962 294400
rect 3018 294344 3023 294400
rect -960 294342 3023 294344
rect -960 294252 480 294342
rect 2957 294339 3023 294342
rect 341241 289914 341307 289917
rect 341374 289914 341380 289916
rect 341241 289912 341380 289914
rect 341241 289856 341246 289912
rect 341302 289856 341380 289912
rect 341241 289854 341380 289856
rect 341241 289851 341307 289854
rect 341374 289852 341380 289854
rect 341444 289852 341450 289916
rect 327165 288418 327231 288421
rect 327533 288418 327599 288421
rect 327165 288416 327599 288418
rect 327165 288360 327170 288416
rect 327226 288360 327538 288416
rect 327594 288360 327599 288416
rect 327165 288358 327599 288360
rect 327165 288355 327231 288358
rect 327533 288355 327599 288358
rect 583520 287316 584960 287556
rect 306741 287058 306807 287061
rect 307017 287058 307083 287061
rect 306741 287056 307083 287058
rect 306741 287000 306746 287056
rect 306802 287000 307022 287056
rect 307078 287000 307083 287056
rect 306741 286998 307083 287000
rect 306741 286995 306807 286998
rect 307017 286995 307083 286998
rect 357433 287058 357499 287061
rect 357801 287058 357867 287061
rect 357433 287056 357867 287058
rect 357433 287000 357438 287056
rect 357494 287000 357806 287056
rect 357862 287000 357867 287056
rect 357433 286998 357867 287000
rect 357433 286995 357499 286998
rect 357801 286995 357867 286998
rect 289997 284338 290063 284341
rect 290273 284338 290339 284341
rect 289997 284336 290339 284338
rect 289997 284280 290002 284336
rect 290058 284280 290278 284336
rect 290334 284280 290339 284336
rect 289997 284278 290339 284280
rect 289997 284275 290063 284278
rect 290273 284275 290339 284278
rect -960 280122 480 280212
rect 4061 280122 4127 280125
rect -960 280120 4127 280122
rect -960 280064 4066 280120
rect 4122 280064 4127 280120
rect -960 280062 4127 280064
rect -960 279972 480 280062
rect 4061 280059 4127 280062
rect 251173 280122 251239 280125
rect 251357 280122 251423 280125
rect 251173 280120 251423 280122
rect 251173 280064 251178 280120
rect 251234 280064 251362 280120
rect 251418 280064 251423 280120
rect 251173 280062 251423 280064
rect 251173 280059 251239 280062
rect 251357 280059 251423 280062
rect 341241 280122 341307 280125
rect 341374 280122 341380 280124
rect 341241 280120 341380 280122
rect 341241 280064 341246 280120
rect 341302 280064 341380 280120
rect 341241 280062 341380 280064
rect 341241 280059 341307 280062
rect 341374 280060 341380 280062
rect 341444 280060 341450 280124
rect 250069 278762 250135 278765
rect 250253 278762 250319 278765
rect 250069 278760 250319 278762
rect 250069 278704 250074 278760
rect 250130 278704 250258 278760
rect 250314 278704 250319 278760
rect 250069 278702 250319 278704
rect 250069 278699 250135 278702
rect 250253 278699 250319 278702
rect 272149 278762 272215 278765
rect 272333 278762 272399 278765
rect 272149 278760 272399 278762
rect 272149 278704 272154 278760
rect 272210 278704 272338 278760
rect 272394 278704 272399 278760
rect 272149 278702 272399 278704
rect 272149 278699 272215 278702
rect 272333 278699 272399 278702
rect 284569 278762 284635 278765
rect 284753 278762 284819 278765
rect 284569 278760 284819 278762
rect 284569 278704 284574 278760
rect 284630 278704 284758 278760
rect 284814 278704 284819 278760
rect 284569 278702 284819 278704
rect 284569 278699 284635 278702
rect 284753 278699 284819 278702
rect 421189 278762 421255 278765
rect 421373 278762 421439 278765
rect 421189 278760 421439 278762
rect 421189 278704 421194 278760
rect 421250 278704 421378 278760
rect 421434 278704 421439 278760
rect 421189 278702 421439 278704
rect 421189 278699 421255 278702
rect 421373 278699 421439 278702
rect 267733 277402 267799 277405
rect 268009 277402 268075 277405
rect 267733 277400 268075 277402
rect 267733 277344 267738 277400
rect 267794 277344 268014 277400
rect 268070 277344 268075 277400
rect 267733 277342 268075 277344
rect 267733 277339 267799 277342
rect 268009 277339 268075 277342
rect 299657 277402 299723 277405
rect 299933 277402 299999 277405
rect 299657 277400 299999 277402
rect 299657 277344 299662 277400
rect 299718 277344 299938 277400
rect 299994 277344 299999 277400
rect 299657 277342 299999 277344
rect 299657 277339 299723 277342
rect 299933 277339 299999 277342
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 249190 275028 249196 275092
rect 249260 275090 249266 275092
rect 249425 275090 249491 275093
rect 249260 275088 249491 275090
rect 249260 275032 249430 275088
rect 249486 275032 249491 275088
rect 249260 275030 249491 275032
rect 249260 275028 249266 275030
rect 249425 275027 249491 275030
rect 341241 270602 341307 270605
rect 341374 270602 341380 270604
rect 341241 270600 341380 270602
rect 341241 270544 341246 270600
rect 341302 270544 341380 270600
rect 341241 270542 341380 270544
rect 341241 270539 341307 270542
rect 341374 270540 341380 270542
rect 341444 270540 341450 270604
rect 249425 267884 249491 267885
rect 249374 267820 249380 267884
rect 249444 267882 249491 267884
rect 249444 267880 249536 267882
rect 249486 267824 249536 267880
rect 249444 267822 249536 267824
rect 249444 267820 249491 267822
rect 249425 267819 249491 267820
rect 244457 267746 244523 267749
rect 244641 267746 244707 267749
rect 244457 267744 244707 267746
rect 244457 267688 244462 267744
rect 244518 267688 244646 267744
rect 244702 267688 244707 267744
rect 244457 267686 244707 267688
rect 244457 267683 244523 267686
rect 244641 267683 244707 267686
rect 245929 267746 245995 267749
rect 246113 267746 246179 267749
rect 245929 267744 246179 267746
rect 245929 267688 245934 267744
rect 245990 267688 246118 267744
rect 246174 267688 246179 267744
rect 245929 267686 246179 267688
rect 245929 267683 245995 267686
rect 246113 267683 246179 267686
rect 294137 267746 294203 267749
rect 294413 267746 294479 267749
rect 294137 267744 294479 267746
rect 294137 267688 294142 267744
rect 294198 267688 294418 267744
rect 294474 267688 294479 267744
rect 294137 267686 294479 267688
rect 294137 267683 294203 267686
rect 294413 267683 294479 267686
rect -960 265706 480 265796
rect 3969 265706 4035 265709
rect -960 265704 4035 265706
rect -960 265648 3974 265704
rect 4030 265648 4035 265704
rect -960 265646 4035 265648
rect -960 265556 480 265646
rect 3969 265643 4035 265646
rect 580901 263938 580967 263941
rect 583520 263938 584960 264028
rect 580901 263936 584960 263938
rect 580901 263880 580906 263936
rect 580962 263880 584960 263936
rect 580901 263878 584960 263880
rect 580901 263875 580967 263878
rect 583520 263788 584960 263878
rect 358721 261218 358787 261221
rect 358721 261216 358922 261218
rect 358721 261160 358726 261216
rect 358782 261160 358922 261216
rect 358721 261158 358922 261160
rect 358721 261155 358787 261158
rect 286041 261082 286107 261085
rect 285814 261080 286107 261082
rect 285814 261024 286046 261080
rect 286102 261024 286107 261080
rect 285814 261022 286107 261024
rect 285814 260946 285874 261022
rect 286041 261019 286107 261022
rect 285949 260946 286015 260949
rect 285814 260944 286015 260946
rect 285814 260888 285954 260944
rect 286010 260888 286015 260944
rect 285814 260886 286015 260888
rect 285949 260883 286015 260886
rect 358721 260946 358787 260949
rect 358862 260946 358922 261158
rect 358721 260944 358922 260946
rect 358721 260888 358726 260944
rect 358782 260888 358922 260944
rect 358721 260886 358922 260888
rect 358721 260883 358787 260886
rect 251173 260810 251239 260813
rect 251357 260810 251423 260813
rect 251173 260808 251423 260810
rect 251173 260752 251178 260808
rect 251234 260752 251362 260808
rect 251418 260752 251423 260808
rect 251173 260750 251423 260752
rect 251173 260747 251239 260750
rect 251357 260747 251423 260750
rect 341241 260810 341307 260813
rect 341374 260810 341380 260812
rect 341241 260808 341380 260810
rect 341241 260752 341246 260808
rect 341302 260752 341380 260808
rect 341241 260750 341380 260752
rect 341241 260747 341307 260750
rect 341374 260748 341380 260750
rect 341444 260748 341450 260812
rect 358537 259450 358603 259453
rect 358721 259450 358787 259453
rect 358537 259448 358787 259450
rect 358537 259392 358542 259448
rect 358598 259392 358726 259448
rect 358782 259392 358787 259448
rect 358537 259390 358787 259392
rect 358537 259387 358603 259390
rect 358721 259387 358787 259390
rect 421189 259450 421255 259453
rect 421373 259450 421439 259453
rect 421189 259448 421439 259450
rect 421189 259392 421194 259448
rect 421250 259392 421378 259448
rect 421434 259392 421439 259448
rect 421189 259390 421439 259392
rect 421189 259387 421255 259390
rect 421373 259387 421439 259390
rect 245837 258090 245903 258093
rect 246113 258090 246179 258093
rect 245837 258088 246179 258090
rect 245837 258032 245842 258088
rect 245898 258032 246118 258088
rect 246174 258032 246179 258088
rect 245837 258030 246179 258032
rect 245837 258027 245903 258030
rect 246113 258027 246179 258030
rect 259729 258090 259795 258093
rect 259913 258090 259979 258093
rect 259729 258088 259979 258090
rect 259729 258032 259734 258088
rect 259790 258032 259918 258088
rect 259974 258032 259979 258088
rect 259729 258030 259979 258032
rect 259729 258027 259795 258030
rect 259913 258027 259979 258030
rect 264973 258090 265039 258093
rect 265157 258090 265223 258093
rect 264973 258088 265223 258090
rect 264973 258032 264978 258088
rect 265034 258032 265162 258088
rect 265218 258032 265223 258088
rect 264973 258030 265223 258032
rect 264973 258027 265039 258030
rect 265157 258027 265223 258030
rect 294229 258090 294295 258093
rect 294413 258090 294479 258093
rect 294229 258088 294479 258090
rect 294229 258032 294234 258088
rect 294290 258032 294418 258088
rect 294474 258032 294479 258088
rect 294229 258030 294479 258032
rect 294229 258027 294295 258030
rect 294413 258027 294479 258030
rect 249241 257956 249307 257957
rect 249190 257892 249196 257956
rect 249260 257954 249307 257956
rect 249260 257952 249352 257954
rect 249302 257896 249352 257952
rect 249260 257894 249352 257896
rect 249260 257892 249307 257894
rect 249241 257891 249307 257892
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 2773 251290 2839 251293
rect -960 251288 2839 251290
rect -960 251232 2778 251288
rect 2834 251232 2839 251288
rect -960 251230 2839 251232
rect -960 251140 480 251230
rect 2773 251227 2839 251230
rect 341241 251290 341307 251293
rect 341374 251290 341380 251292
rect 341241 251288 341380 251290
rect 341241 251232 341246 251288
rect 341302 251232 341380 251288
rect 341241 251230 341380 251232
rect 341241 251227 341307 251230
rect 341374 251228 341380 251230
rect 341444 251228 341450 251292
rect 388989 251154 389055 251157
rect 389173 251154 389239 251157
rect 388989 251152 389239 251154
rect 388989 251096 388994 251152
rect 389050 251096 389178 251152
rect 389234 251096 389239 251152
rect 388989 251094 389239 251096
rect 388989 251091 389055 251094
rect 389173 251091 389239 251094
rect 336733 249930 336799 249933
rect 337101 249930 337167 249933
rect 336733 249928 337167 249930
rect 336733 249872 336738 249928
rect 336794 249872 337106 249928
rect 337162 249872 337167 249928
rect 336733 249870 337167 249872
rect 336733 249867 336799 249870
rect 337101 249867 337167 249870
rect 232221 249794 232287 249797
rect 232497 249794 232563 249797
rect 286041 249794 286107 249797
rect 232221 249792 232563 249794
rect 232221 249736 232226 249792
rect 232282 249736 232502 249792
rect 232558 249736 232563 249792
rect 232221 249734 232563 249736
rect 232221 249731 232287 249734
rect 232497 249731 232563 249734
rect 285998 249792 286107 249794
rect 285998 249736 286046 249792
rect 286102 249736 286107 249792
rect 285998 249731 286107 249736
rect 302417 249794 302483 249797
rect 302601 249794 302667 249797
rect 302417 249792 302667 249794
rect 302417 249736 302422 249792
rect 302478 249736 302606 249792
rect 302662 249736 302667 249792
rect 302417 249734 302667 249736
rect 302417 249731 302483 249734
rect 302601 249731 302667 249734
rect 306925 249794 306991 249797
rect 307109 249794 307175 249797
rect 306925 249792 307175 249794
rect 306925 249736 306930 249792
rect 306986 249736 307114 249792
rect 307170 249736 307175 249792
rect 306925 249734 307175 249736
rect 306925 249731 306991 249734
rect 307109 249731 307175 249734
rect 325877 249794 325943 249797
rect 326153 249794 326219 249797
rect 325877 249792 326219 249794
rect 325877 249736 325882 249792
rect 325938 249736 326158 249792
rect 326214 249736 326219 249792
rect 325877 249734 326219 249736
rect 325877 249731 325943 249734
rect 326153 249731 326219 249734
rect 337101 249794 337167 249797
rect 337285 249794 337351 249797
rect 337101 249792 337351 249794
rect 337101 249736 337106 249792
rect 337162 249736 337290 249792
rect 337346 249736 337351 249792
rect 337101 249734 337351 249736
rect 337101 249731 337167 249734
rect 337285 249731 337351 249734
rect 285998 249661 286058 249731
rect 285949 249656 286058 249661
rect 285949 249600 285954 249656
rect 286010 249600 286058 249656
rect 285949 249598 286058 249600
rect 285949 249595 286015 249598
rect 249006 248372 249012 248436
rect 249076 248434 249082 248436
rect 249241 248434 249307 248437
rect 249076 248432 249307 248434
rect 249076 248376 249246 248432
rect 249302 248376 249307 248432
rect 249076 248374 249307 248376
rect 249076 248372 249082 248374
rect 249241 248371 249307 248374
rect 288801 248434 288867 248437
rect 288985 248434 289051 248437
rect 288801 248432 289051 248434
rect 288801 248376 288806 248432
rect 288862 248376 288990 248432
rect 289046 248376 289051 248432
rect 288801 248374 289051 248376
rect 288801 248371 288867 248374
rect 288985 248371 289051 248374
rect 296897 248434 296963 248437
rect 297173 248434 297239 248437
rect 296897 248432 297239 248434
rect 296897 248376 296902 248432
rect 296958 248376 297178 248432
rect 297234 248376 297239 248432
rect 296897 248374 297239 248376
rect 296897 248371 296963 248374
rect 297173 248371 297239 248374
rect 330201 248434 330267 248437
rect 330385 248434 330451 248437
rect 330201 248432 330451 248434
rect 330201 248376 330206 248432
rect 330262 248376 330390 248432
rect 330446 248376 330451 248432
rect 330201 248374 330451 248376
rect 330201 248371 330267 248374
rect 330385 248371 330451 248374
rect 421189 241770 421255 241773
rect 421054 241768 421255 241770
rect 421054 241712 421194 241768
rect 421250 241712 421255 241768
rect 421054 241710 421255 241712
rect 421054 241634 421114 241710
rect 421189 241707 421255 241710
rect 421189 241634 421255 241637
rect 421054 241632 421255 241634
rect 421054 241576 421194 241632
rect 421250 241576 421255 241632
rect 421054 241574 421255 241576
rect 421189 241571 421255 241574
rect 272149 241498 272215 241501
rect 301037 241498 301103 241501
rect 366817 241498 366883 241501
rect 367001 241498 367067 241501
rect 272149 241496 272258 241498
rect 272149 241440 272154 241496
rect 272210 241440 272258 241496
rect 272149 241435 272258 241440
rect 301037 241496 301146 241498
rect 301037 241440 301042 241496
rect 301098 241440 301146 241496
rect 301037 241435 301146 241440
rect 366817 241496 367067 241498
rect 366817 241440 366822 241496
rect 366878 241440 367006 241496
rect 367062 241440 367067 241496
rect 366817 241438 367067 241440
rect 366817 241435 366883 241438
rect 367001 241435 367067 241438
rect 372521 241498 372587 241501
rect 372705 241498 372771 241501
rect 372521 241496 372771 241498
rect 372521 241440 372526 241496
rect 372582 241440 372710 241496
rect 372766 241440 372771 241496
rect 372521 241438 372771 241440
rect 372521 241435 372587 241438
rect 372705 241435 372771 241438
rect 376937 241498 377003 241501
rect 377121 241498 377187 241501
rect 376937 241496 377187 241498
rect 376937 241440 376942 241496
rect 376998 241440 377126 241496
rect 377182 241440 377187 241496
rect 376937 241438 377187 241440
rect 376937 241435 377003 241438
rect 377121 241435 377187 241438
rect 272198 241362 272258 241435
rect 301086 241365 301146 241435
rect 272333 241362 272399 241365
rect 272198 241360 272399 241362
rect 272198 241304 272338 241360
rect 272394 241304 272399 241360
rect 272198 241302 272399 241304
rect 301086 241360 301195 241365
rect 301086 241304 301134 241360
rect 301190 241304 301195 241360
rect 301086 241302 301195 241304
rect 272333 241299 272399 241302
rect 301129 241299 301195 241302
rect 583520 240396 584960 240636
rect 239305 240138 239371 240141
rect 239489 240138 239555 240141
rect 239305 240136 239555 240138
rect 239305 240080 239310 240136
rect 239366 240080 239494 240136
rect 239550 240080 239555 240136
rect 239305 240078 239555 240080
rect 239305 240075 239371 240078
rect 239489 240075 239555 240078
rect 245837 240138 245903 240141
rect 246113 240138 246179 240141
rect 245837 240136 246179 240138
rect 245837 240080 245842 240136
rect 245898 240080 246118 240136
rect 246174 240080 246179 240136
rect 245837 240078 246179 240080
rect 245837 240075 245903 240078
rect 246113 240075 246179 240078
rect 251081 240138 251147 240141
rect 251357 240138 251423 240141
rect 251081 240136 251423 240138
rect 251081 240080 251086 240136
rect 251142 240080 251362 240136
rect 251418 240080 251423 240136
rect 251081 240078 251423 240080
rect 251081 240075 251147 240078
rect 251357 240075 251423 240078
rect 259637 240138 259703 240141
rect 259821 240138 259887 240141
rect 259637 240136 259887 240138
rect 259637 240080 259642 240136
rect 259698 240080 259826 240136
rect 259882 240080 259887 240136
rect 259637 240078 259887 240080
rect 259637 240075 259703 240078
rect 259821 240075 259887 240078
rect 267917 240138 267983 240141
rect 268101 240138 268167 240141
rect 267917 240136 268167 240138
rect 267917 240080 267922 240136
rect 267978 240080 268106 240136
rect 268162 240080 268167 240136
rect 267917 240078 268167 240080
rect 267917 240075 267983 240078
rect 268101 240075 268167 240078
rect 341149 240138 341215 240141
rect 341425 240138 341491 240141
rect 341149 240136 341491 240138
rect 341149 240080 341154 240136
rect 341210 240080 341430 240136
rect 341486 240080 341491 240136
rect 341149 240078 341491 240080
rect 341149 240075 341215 240078
rect 341425 240075 341491 240078
rect 358537 240138 358603 240141
rect 358721 240138 358787 240141
rect 358537 240136 358787 240138
rect 358537 240080 358542 240136
rect 358598 240080 358726 240136
rect 358782 240080 358787 240136
rect 358537 240078 358787 240080
rect 358537 240075 358603 240078
rect 358721 240075 358787 240078
rect 421189 240138 421255 240141
rect 421373 240138 421439 240141
rect 421189 240136 421439 240138
rect 421189 240080 421194 240136
rect 421250 240080 421378 240136
rect 421434 240080 421439 240136
rect 421189 240078 421439 240080
rect 421189 240075 421255 240078
rect 421373 240075 421439 240078
rect -960 237010 480 237100
rect 3049 237010 3115 237013
rect -960 237008 3115 237010
rect -960 236952 3054 237008
rect 3110 236952 3115 237008
rect -960 236950 3115 236952
rect -960 236860 480 236950
rect 3049 236947 3115 236950
rect 389265 231842 389331 231845
rect 389449 231842 389515 231845
rect 389265 231840 389515 231842
rect 389265 231784 389270 231840
rect 389326 231784 389454 231840
rect 389510 231784 389515 231840
rect 389265 231782 389515 231784
rect 389265 231779 389331 231782
rect 389449 231779 389515 231782
rect 463785 231842 463851 231845
rect 463969 231842 464035 231845
rect 463785 231840 464035 231842
rect 463785 231784 463790 231840
rect 463846 231784 463974 231840
rect 464030 231784 464035 231840
rect 463785 231782 464035 231784
rect 463785 231779 463851 231782
rect 463969 231779 464035 231782
rect 470409 231842 470475 231845
rect 470593 231842 470659 231845
rect 470409 231840 470659 231842
rect 470409 231784 470414 231840
rect 470470 231784 470598 231840
rect 470654 231784 470659 231840
rect 470409 231782 470659 231784
rect 470409 231779 470475 231782
rect 470593 231779 470659 231782
rect 249006 230556 249012 230620
rect 249076 230618 249082 230620
rect 249076 230558 249442 230618
rect 249076 230556 249082 230558
rect 232221 230482 232287 230485
rect 232497 230482 232563 230485
rect 249382 230484 249442 230558
rect 232221 230480 232563 230482
rect 232221 230424 232226 230480
rect 232282 230424 232502 230480
rect 232558 230424 232563 230480
rect 232221 230422 232563 230424
rect 232221 230419 232287 230422
rect 232497 230419 232563 230422
rect 249374 230420 249380 230484
rect 249444 230420 249450 230484
rect 251357 230482 251423 230485
rect 251541 230482 251607 230485
rect 251357 230480 251607 230482
rect 251357 230424 251362 230480
rect 251418 230424 251546 230480
rect 251602 230424 251607 230480
rect 251357 230422 251607 230424
rect 251357 230419 251423 230422
rect 251541 230419 251607 230422
rect 327165 230482 327231 230485
rect 327533 230482 327599 230485
rect 327165 230480 327599 230482
rect 327165 230424 327170 230480
rect 327226 230424 327538 230480
rect 327594 230424 327599 230480
rect 327165 230422 327599 230424
rect 327165 230419 327231 230422
rect 327533 230419 327599 230422
rect 337193 230482 337259 230485
rect 337377 230482 337443 230485
rect 337193 230480 337443 230482
rect 337193 230424 337198 230480
rect 337254 230424 337382 230480
rect 337438 230424 337443 230480
rect 337193 230422 337443 230424
rect 337193 230419 337259 230422
rect 337377 230419 337443 230422
rect 330201 229122 330267 229125
rect 330385 229122 330451 229125
rect 330201 229120 330451 229122
rect 330201 229064 330206 229120
rect 330262 229064 330390 229120
rect 330446 229064 330451 229120
rect 330201 229062 330451 229064
rect 330201 229059 330267 229062
rect 330385 229059 330451 229062
rect 580809 228850 580875 228853
rect 583520 228850 584960 228940
rect 580809 228848 584960 228850
rect 580809 228792 580814 228848
rect 580870 228792 584960 228848
rect 580809 228790 584960 228792
rect 580809 228787 580875 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3877 222594 3943 222597
rect -960 222592 3943 222594
rect -960 222536 3882 222592
rect 3938 222536 3943 222592
rect -960 222534 3943 222536
rect -960 222444 480 222534
rect 3877 222531 3943 222534
rect 259637 222186 259703 222189
rect 259502 222184 259703 222186
rect 259502 222128 259642 222184
rect 259698 222128 259703 222184
rect 259502 222126 259703 222128
rect 259502 221914 259562 222126
rect 259637 222123 259703 222126
rect 272149 222186 272215 222189
rect 285949 222186 286015 222189
rect 286133 222186 286199 222189
rect 272149 222184 272258 222186
rect 272149 222128 272154 222184
rect 272210 222128 272258 222184
rect 272149 222123 272258 222128
rect 285949 222184 286199 222186
rect 285949 222128 285954 222184
rect 286010 222128 286138 222184
rect 286194 222128 286199 222184
rect 285949 222126 286199 222128
rect 285949 222123 286015 222126
rect 286133 222123 286199 222126
rect 301037 222186 301103 222189
rect 372521 222186 372587 222189
rect 372705 222186 372771 222189
rect 301037 222184 301146 222186
rect 301037 222128 301042 222184
rect 301098 222128 301146 222184
rect 301037 222123 301146 222128
rect 372521 222184 372771 222186
rect 372521 222128 372526 222184
rect 372582 222128 372710 222184
rect 372766 222128 372771 222184
rect 372521 222126 372771 222128
rect 372521 222123 372587 222126
rect 372705 222123 372771 222126
rect 376937 222186 377003 222189
rect 377121 222186 377187 222189
rect 376937 222184 377187 222186
rect 376937 222128 376942 222184
rect 376998 222128 377126 222184
rect 377182 222128 377187 222184
rect 376937 222126 377187 222128
rect 376937 222123 377003 222126
rect 377121 222123 377187 222126
rect 272198 222053 272258 222123
rect 301086 222053 301146 222123
rect 272198 222048 272307 222053
rect 272198 221992 272246 222048
rect 272302 221992 272307 222048
rect 272198 221990 272307 221992
rect 301086 222048 301195 222053
rect 301086 221992 301134 222048
rect 301190 221992 301195 222048
rect 301086 221990 301195 221992
rect 272241 221987 272307 221990
rect 301129 221987 301195 221990
rect 259729 221914 259795 221917
rect 259502 221912 259795 221914
rect 259502 221856 259734 221912
rect 259790 221856 259795 221912
rect 259502 221854 259795 221856
rect 259729 221851 259795 221854
rect 284661 220826 284727 220829
rect 284845 220826 284911 220829
rect 284661 220824 284911 220826
rect 284661 220768 284666 220824
rect 284722 220768 284850 220824
rect 284906 220768 284911 220824
rect 284661 220766 284911 220768
rect 284661 220763 284727 220766
rect 284845 220763 284911 220766
rect 285949 220826 286015 220829
rect 286133 220826 286199 220829
rect 285949 220824 286199 220826
rect 285949 220768 285954 220824
rect 286010 220768 286138 220824
rect 286194 220768 286199 220824
rect 285949 220766 286199 220768
rect 285949 220763 286015 220766
rect 286133 220763 286199 220766
rect 358537 220826 358603 220829
rect 358721 220826 358787 220829
rect 358537 220824 358787 220826
rect 358537 220768 358542 220824
rect 358598 220768 358726 220824
rect 358782 220768 358787 220824
rect 358537 220766 358787 220768
rect 358537 220763 358603 220766
rect 358721 220763 358787 220766
rect 421189 220826 421255 220829
rect 421373 220826 421439 220829
rect 421189 220824 421439 220826
rect 421189 220768 421194 220824
rect 421250 220768 421378 220824
rect 421434 220768 421439 220824
rect 421189 220766 421439 220768
rect 421189 220763 421255 220766
rect 421373 220763 421439 220766
rect 244273 219466 244339 219469
rect 244549 219466 244615 219469
rect 244273 219464 244615 219466
rect 244273 219408 244278 219464
rect 244334 219408 244554 219464
rect 244610 219408 244615 219464
rect 244273 219406 244615 219408
rect 244273 219403 244339 219406
rect 244549 219403 244615 219406
rect 329925 219466 329991 219469
rect 330109 219466 330175 219469
rect 329925 219464 330175 219466
rect 329925 219408 329930 219464
rect 329986 219408 330114 219464
rect 330170 219408 330175 219464
rect 329925 219406 330175 219408
rect 329925 219403 329991 219406
rect 330109 219403 330175 219406
rect 249374 219268 249380 219332
rect 249444 219268 249450 219332
rect 249382 219194 249442 219268
rect 249742 219194 249748 219196
rect 249382 219134 249748 219194
rect 249742 219132 249748 219134
rect 249812 219132 249818 219196
rect 580717 217018 580783 217021
rect 583520 217018 584960 217108
rect 580717 217016 584960 217018
rect 580717 216960 580722 217016
rect 580778 216960 584960 217016
rect 580717 216958 584960 216960
rect 580717 216955 580783 216958
rect 583520 216868 584960 216958
rect 239121 212530 239187 212533
rect 239305 212530 239371 212533
rect 327257 212530 327323 212533
rect 239121 212528 239371 212530
rect 239121 212472 239126 212528
rect 239182 212472 239310 212528
rect 239366 212472 239371 212528
rect 239121 212470 239371 212472
rect 239121 212467 239187 212470
rect 239305 212467 239371 212470
rect 327214 212528 327323 212530
rect 327214 212472 327262 212528
rect 327318 212472 327323 212528
rect 327214 212467 327323 212472
rect 389265 212530 389331 212533
rect 389449 212530 389515 212533
rect 389265 212528 389515 212530
rect 389265 212472 389270 212528
rect 389326 212472 389454 212528
rect 389510 212472 389515 212528
rect 389265 212470 389515 212472
rect 389265 212467 389331 212470
rect 389449 212467 389515 212470
rect 424593 212530 424659 212533
rect 424777 212530 424843 212533
rect 424593 212528 424843 212530
rect 424593 212472 424598 212528
rect 424654 212472 424782 212528
rect 424838 212472 424843 212528
rect 424593 212470 424843 212472
rect 424593 212467 424659 212470
rect 424777 212467 424843 212470
rect 463785 212530 463851 212533
rect 463969 212530 464035 212533
rect 463785 212528 464035 212530
rect 463785 212472 463790 212528
rect 463846 212472 463974 212528
rect 464030 212472 464035 212528
rect 463785 212470 464035 212472
rect 463785 212467 463851 212470
rect 463969 212467 464035 212470
rect 470409 212530 470475 212533
rect 470593 212530 470659 212533
rect 470409 212528 470659 212530
rect 470409 212472 470414 212528
rect 470470 212472 470598 212528
rect 470654 212472 470659 212528
rect 470409 212470 470659 212472
rect 470409 212467 470475 212470
rect 470593 212467 470659 212470
rect 327214 212394 327274 212467
rect 327349 212394 327415 212397
rect 327214 212392 327415 212394
rect 327214 212336 327354 212392
rect 327410 212336 327415 212392
rect 327214 212334 327415 212336
rect 327349 212331 327415 212334
rect 323301 211170 323367 211173
rect 323485 211170 323551 211173
rect 323301 211168 323551 211170
rect 323301 211112 323306 211168
rect 323362 211112 323490 211168
rect 323546 211112 323551 211168
rect 323301 211110 323551 211112
rect 323301 211107 323367 211110
rect 323485 211107 323551 211110
rect 249609 209674 249675 209677
rect 249742 209674 249748 209676
rect 249609 209672 249748 209674
rect 249609 209616 249614 209672
rect 249670 209616 249748 209672
rect 249609 209614 249748 209616
rect 249609 209611 249675 209614
rect 249742 209612 249748 209614
rect 249812 209612 249818 209676
rect -960 208178 480 208268
rect 3785 208178 3851 208181
rect -960 208176 3851 208178
rect -960 208120 3790 208176
rect 3846 208120 3851 208176
rect -960 208118 3851 208120
rect -960 208028 480 208118
rect 3785 208115 3851 208118
rect 580625 205322 580691 205325
rect 583520 205322 584960 205412
rect 580625 205320 584960 205322
rect 580625 205264 580630 205320
rect 580686 205264 584960 205320
rect 580625 205262 584960 205264
rect 580625 205259 580691 205262
rect 583520 205172 584960 205262
rect 259637 202874 259703 202877
rect 259913 202874 259979 202877
rect 270677 202874 270743 202877
rect 272149 202874 272215 202877
rect 259637 202872 259979 202874
rect 259637 202816 259642 202872
rect 259698 202816 259918 202872
rect 259974 202816 259979 202872
rect 259637 202814 259979 202816
rect 259637 202811 259703 202814
rect 259913 202811 259979 202814
rect 270542 202872 270743 202874
rect 270542 202816 270682 202872
rect 270738 202816 270743 202872
rect 270542 202814 270743 202816
rect 270542 202738 270602 202814
rect 270677 202811 270743 202814
rect 272014 202872 272215 202874
rect 272014 202816 272154 202872
rect 272210 202816 272215 202872
rect 272014 202814 272215 202816
rect 270677 202738 270743 202741
rect 270542 202736 270743 202738
rect 270542 202680 270682 202736
rect 270738 202680 270743 202736
rect 270542 202678 270743 202680
rect 272014 202738 272074 202814
rect 272149 202811 272215 202814
rect 285765 202874 285831 202877
rect 285949 202874 286015 202877
rect 285765 202872 286015 202874
rect 285765 202816 285770 202872
rect 285826 202816 285954 202872
rect 286010 202816 286015 202872
rect 285765 202814 286015 202816
rect 285765 202811 285831 202814
rect 285949 202811 286015 202814
rect 301037 202874 301103 202877
rect 325877 202874 325943 202877
rect 337101 202874 337167 202877
rect 337377 202874 337443 202877
rect 301037 202872 301146 202874
rect 301037 202816 301042 202872
rect 301098 202816 301146 202872
rect 301037 202811 301146 202816
rect 325877 202872 325986 202874
rect 325877 202816 325882 202872
rect 325938 202816 325986 202872
rect 325877 202811 325986 202816
rect 337101 202872 337443 202874
rect 337101 202816 337106 202872
rect 337162 202816 337382 202872
rect 337438 202816 337443 202872
rect 337101 202814 337443 202816
rect 337101 202811 337167 202814
rect 337377 202811 337443 202814
rect 341149 202874 341215 202877
rect 341425 202874 341491 202877
rect 341149 202872 341491 202874
rect 341149 202816 341154 202872
rect 341210 202816 341430 202872
rect 341486 202816 341491 202872
rect 341149 202814 341491 202816
rect 341149 202811 341215 202814
rect 341425 202811 341491 202814
rect 366817 202874 366883 202877
rect 367001 202874 367067 202877
rect 366817 202872 367067 202874
rect 366817 202816 366822 202872
rect 366878 202816 367006 202872
rect 367062 202816 367067 202872
rect 366817 202814 367067 202816
rect 366817 202811 366883 202814
rect 367001 202811 367067 202814
rect 372521 202874 372587 202877
rect 372705 202874 372771 202877
rect 372521 202872 372771 202874
rect 372521 202816 372526 202872
rect 372582 202816 372710 202872
rect 372766 202816 372771 202872
rect 372521 202814 372771 202816
rect 372521 202811 372587 202814
rect 372705 202811 372771 202814
rect 376937 202874 377003 202877
rect 377121 202874 377187 202877
rect 376937 202872 377187 202874
rect 376937 202816 376942 202872
rect 376998 202816 377126 202872
rect 377182 202816 377187 202872
rect 376937 202814 377187 202816
rect 376937 202811 377003 202814
rect 377121 202811 377187 202814
rect 301086 202741 301146 202811
rect 325926 202741 325986 202811
rect 272241 202738 272307 202741
rect 272014 202736 272307 202738
rect 272014 202680 272246 202736
rect 272302 202680 272307 202736
rect 272014 202678 272307 202680
rect 301086 202736 301195 202741
rect 301086 202680 301134 202736
rect 301190 202680 301195 202736
rect 301086 202678 301195 202680
rect 325926 202736 326035 202741
rect 325926 202680 325974 202736
rect 326030 202680 326035 202736
rect 325926 202678 326035 202680
rect 270677 202675 270743 202678
rect 272241 202675 272307 202678
rect 301129 202675 301195 202678
rect 325969 202675 326035 202678
rect 239029 201514 239095 201517
rect 239213 201514 239279 201517
rect 239029 201512 239279 201514
rect 239029 201456 239034 201512
rect 239090 201456 239218 201512
rect 239274 201456 239279 201512
rect 239029 201454 239279 201456
rect 239029 201451 239095 201454
rect 239213 201451 239279 201454
rect 249609 200156 249675 200157
rect 249558 200154 249564 200156
rect 249518 200094 249564 200154
rect 249628 200152 249675 200156
rect 249670 200096 249675 200152
rect 249558 200092 249564 200094
rect 249628 200092 249675 200096
rect 249609 200091 249675 200092
rect 421097 196618 421163 196621
rect 421230 196618 421236 196620
rect 421097 196616 421236 196618
rect 421097 196560 421102 196616
rect 421158 196560 421236 196616
rect 421097 196558 421236 196560
rect 421097 196555 421163 196558
rect 421230 196556 421236 196558
rect 421300 196556 421306 196620
rect -960 193898 480 193988
rect 3693 193898 3759 193901
rect -960 193896 3759 193898
rect -960 193840 3698 193896
rect 3754 193840 3759 193896
rect -960 193838 3759 193840
rect -960 193748 480 193838
rect 3693 193835 3759 193838
rect 583520 193476 584960 193716
rect 249333 193218 249399 193221
rect 249558 193218 249564 193220
rect 249333 193216 249564 193218
rect 249333 193160 249338 193216
rect 249394 193160 249564 193216
rect 249333 193158 249564 193160
rect 249333 193155 249399 193158
rect 249558 193156 249564 193158
rect 249628 193156 249634 193220
rect 250069 193218 250135 193221
rect 250253 193218 250319 193221
rect 250069 193216 250319 193218
rect 250069 193160 250074 193216
rect 250130 193160 250258 193216
rect 250314 193160 250319 193216
rect 250069 193158 250319 193160
rect 250069 193155 250135 193158
rect 250253 193155 250319 193158
rect 310789 193218 310855 193221
rect 311065 193218 311131 193221
rect 310789 193216 311131 193218
rect 310789 193160 310794 193216
rect 310850 193160 311070 193216
rect 311126 193160 311131 193216
rect 310789 193158 311131 193160
rect 310789 193155 310855 193158
rect 311065 193155 311131 193158
rect 323301 193218 323367 193221
rect 323485 193218 323551 193221
rect 323301 193216 323551 193218
rect 323301 193160 323306 193216
rect 323362 193160 323490 193216
rect 323546 193160 323551 193216
rect 323301 193158 323551 193160
rect 323301 193155 323367 193158
rect 323485 193155 323551 193158
rect 389265 193218 389331 193221
rect 389449 193218 389515 193221
rect 389265 193216 389515 193218
rect 389265 193160 389270 193216
rect 389326 193160 389454 193216
rect 389510 193160 389515 193216
rect 389265 193158 389515 193160
rect 389265 193155 389331 193158
rect 389449 193155 389515 193158
rect 463785 193218 463851 193221
rect 463969 193218 464035 193221
rect 463785 193216 464035 193218
rect 463785 193160 463790 193216
rect 463846 193160 463974 193216
rect 464030 193160 464035 193216
rect 463785 193158 464035 193160
rect 463785 193155 463851 193158
rect 463969 193155 464035 193158
rect 470409 193218 470475 193221
rect 470593 193218 470659 193221
rect 470409 193216 470659 193218
rect 470409 193160 470414 193216
rect 470470 193160 470598 193216
rect 470654 193160 470659 193216
rect 470409 193158 470659 193160
rect 470409 193155 470475 193158
rect 470593 193155 470659 193158
rect 421189 183700 421255 183701
rect 421189 183698 421236 183700
rect 421144 183696 421236 183698
rect 421144 183640 421194 183696
rect 421144 183638 421236 183640
rect 421189 183636 421236 183638
rect 421300 183636 421306 183700
rect 421189 183635 421255 183636
rect 267733 183562 267799 183565
rect 267917 183562 267983 183565
rect 267733 183560 267983 183562
rect 267733 183504 267738 183560
rect 267794 183504 267922 183560
rect 267978 183504 267983 183560
rect 267733 183502 267983 183504
rect 267733 183499 267799 183502
rect 267917 183499 267983 183502
rect 270493 183562 270559 183565
rect 270677 183562 270743 183565
rect 270493 183560 270743 183562
rect 270493 183504 270498 183560
rect 270554 183504 270682 183560
rect 270738 183504 270743 183560
rect 270493 183502 270743 183504
rect 270493 183499 270559 183502
rect 270677 183499 270743 183502
rect 327165 183562 327231 183565
rect 327349 183562 327415 183565
rect 327165 183560 327415 183562
rect 327165 183504 327170 183560
rect 327226 183504 327354 183560
rect 327410 183504 327415 183560
rect 327165 183502 327415 183504
rect 327165 183499 327231 183502
rect 327349 183499 327415 183502
rect 330109 183562 330175 183565
rect 336733 183562 336799 183565
rect 336917 183562 336983 183565
rect 330109 183560 330218 183562
rect 330109 183504 330114 183560
rect 330170 183504 330218 183560
rect 330109 183499 330218 183504
rect 336733 183560 336983 183562
rect 336733 183504 336738 183560
rect 336794 183504 336922 183560
rect 336978 183504 336983 183560
rect 336733 183502 336983 183504
rect 336733 183499 336799 183502
rect 336917 183499 336983 183502
rect 376937 183562 377003 183565
rect 377121 183562 377187 183565
rect 376937 183560 377187 183562
rect 376937 183504 376942 183560
rect 376998 183504 377126 183560
rect 377182 183504 377187 183560
rect 376937 183502 377187 183504
rect 376937 183499 377003 183502
rect 377121 183499 377187 183502
rect 330158 183429 330218 183499
rect 330109 183424 330218 183429
rect 330109 183368 330114 183424
rect 330170 183368 330218 183424
rect 330109 183366 330218 183368
rect 330109 183363 330175 183366
rect 360469 182474 360535 182477
rect 360150 182472 360535 182474
rect 360150 182416 360474 182472
rect 360530 182416 360535 182472
rect 360150 182414 360535 182416
rect 249006 182140 249012 182204
rect 249076 182202 249082 182204
rect 249333 182202 249399 182205
rect 249076 182200 249399 182202
rect 249076 182144 249338 182200
rect 249394 182144 249399 182200
rect 249076 182142 249399 182144
rect 249076 182140 249082 182142
rect 249333 182139 249399 182142
rect 324589 182202 324655 182205
rect 324865 182202 324931 182205
rect 324589 182200 324931 182202
rect 324589 182144 324594 182200
rect 324650 182144 324870 182200
rect 324926 182144 324931 182200
rect 324589 182142 324931 182144
rect 324589 182139 324655 182142
rect 324865 182139 324931 182142
rect 357525 182202 357591 182205
rect 357709 182202 357775 182205
rect 357525 182200 357775 182202
rect 357525 182144 357530 182200
rect 357586 182144 357714 182200
rect 357770 182144 357775 182200
rect 357525 182142 357775 182144
rect 357525 182139 357591 182142
rect 357709 182139 357775 182142
rect 358997 182202 359063 182205
rect 359181 182202 359247 182205
rect 358997 182200 359247 182202
rect 358997 182144 359002 182200
rect 359058 182144 359186 182200
rect 359242 182144 359247 182200
rect 358997 182142 359247 182144
rect 360150 182202 360210 182414
rect 360469 182411 360535 182414
rect 360285 182202 360351 182205
rect 360150 182200 360351 182202
rect 360150 182144 360290 182200
rect 360346 182144 360351 182200
rect 360150 182142 360351 182144
rect 358997 182139 359063 182142
rect 359181 182139 359247 182142
rect 360285 182139 360351 182142
rect 580533 181930 580599 181933
rect 583520 181930 584960 182020
rect 580533 181928 584960 181930
rect 580533 181872 580538 181928
rect 580594 181872 584960 181928
rect 580533 181870 584960 181872
rect 580533 181867 580599 181870
rect 583520 181780 584960 181870
rect 288801 180842 288867 180845
rect 288985 180842 289051 180845
rect 288801 180840 289051 180842
rect 288801 180784 288806 180840
rect 288862 180784 288990 180840
rect 289046 180784 289051 180840
rect 288801 180782 289051 180784
rect 288801 180779 288867 180782
rect 288985 180779 289051 180782
rect -960 179482 480 179572
rect 3601 179482 3667 179485
rect -960 179480 3667 179482
rect -960 179424 3606 179480
rect 3662 179424 3667 179480
rect -960 179422 3667 179424
rect -960 179332 480 179422
rect 3601 179419 3667 179422
rect 372797 173906 372863 173909
rect 372981 173906 373047 173909
rect 372797 173904 373047 173906
rect 372797 173848 372802 173904
rect 372858 173848 372986 173904
rect 373042 173848 373047 173904
rect 372797 173846 373047 173848
rect 372797 173843 372863 173846
rect 372981 173843 373047 173846
rect 470409 173906 470475 173909
rect 470593 173906 470659 173909
rect 470409 173904 470659 173906
rect 470409 173848 470414 173904
rect 470470 173848 470598 173904
rect 470654 173848 470659 173904
rect 470409 173846 470659 173848
rect 470409 173843 470475 173846
rect 470593 173843 470659 173846
rect 289997 172682 290063 172685
rect 291469 172682 291535 172685
rect 289997 172680 290106 172682
rect 289997 172624 290002 172680
rect 290058 172624 290106 172680
rect 289997 172619 290106 172624
rect 291469 172680 291578 172682
rect 291469 172624 291474 172680
rect 291530 172624 291578 172680
rect 291469 172619 291578 172624
rect 290046 172549 290106 172619
rect 291518 172549 291578 172619
rect 236269 172546 236335 172549
rect 236453 172546 236519 172549
rect 236269 172544 236519 172546
rect 236269 172488 236274 172544
rect 236330 172488 236458 172544
rect 236514 172488 236519 172544
rect 236269 172486 236519 172488
rect 236269 172483 236335 172486
rect 236453 172483 236519 172486
rect 289997 172544 290106 172549
rect 289997 172488 290002 172544
rect 290058 172488 290106 172544
rect 289997 172486 290106 172488
rect 291469 172544 291578 172549
rect 291469 172488 291474 172544
rect 291530 172488 291578 172544
rect 291469 172486 291578 172488
rect 327257 172546 327323 172549
rect 327533 172546 327599 172549
rect 327257 172544 327599 172546
rect 327257 172488 327262 172544
rect 327318 172488 327538 172544
rect 327594 172488 327599 172544
rect 327257 172486 327599 172488
rect 289997 172483 290063 172486
rect 291469 172483 291535 172486
rect 327257 172483 327323 172486
rect 327533 172483 327599 172486
rect 329925 172546 329991 172549
rect 330201 172546 330267 172549
rect 329925 172544 330267 172546
rect 329925 172488 329930 172544
rect 329986 172488 330206 172544
rect 330262 172488 330267 172544
rect 329925 172486 330267 172488
rect 329925 172483 329991 172486
rect 330201 172483 330267 172486
rect 339493 172546 339559 172549
rect 339861 172546 339927 172549
rect 339493 172544 339927 172546
rect 339493 172488 339498 172544
rect 339554 172488 339866 172544
rect 339922 172488 339927 172544
rect 339493 172486 339927 172488
rect 339493 172483 339559 172486
rect 339861 172483 339927 172486
rect 358537 172546 358603 172549
rect 358721 172546 358787 172549
rect 358537 172544 358787 172546
rect 358537 172488 358542 172544
rect 358598 172488 358726 172544
rect 358782 172488 358787 172544
rect 358537 172486 358787 172488
rect 358537 172483 358603 172486
rect 358721 172483 358787 172486
rect 421189 172546 421255 172549
rect 421373 172546 421439 172549
rect 421189 172544 421439 172546
rect 421189 172488 421194 172544
rect 421250 172488 421378 172544
rect 421434 172488 421439 172544
rect 421189 172486 421439 172488
rect 421189 172483 421255 172486
rect 421373 172483 421439 172486
rect 580441 170098 580507 170101
rect 583520 170098 584960 170188
rect 580441 170096 584960 170098
rect 580441 170040 580446 170096
rect 580502 170040 584960 170096
rect 580441 170038 584960 170040
rect 580441 170035 580507 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 245929 164250 245995 164253
rect 245702 164248 245995 164250
rect 245702 164192 245934 164248
rect 245990 164192 245995 164248
rect 245702 164190 245995 164192
rect 245702 164114 245762 164190
rect 245929 164187 245995 164190
rect 270493 164250 270559 164253
rect 270677 164250 270743 164253
rect 270493 164248 270743 164250
rect 270493 164192 270498 164248
rect 270554 164192 270682 164248
rect 270738 164192 270743 164248
rect 270493 164190 270743 164192
rect 270493 164187 270559 164190
rect 270677 164187 270743 164190
rect 272057 164250 272123 164253
rect 272241 164250 272307 164253
rect 272057 164248 272307 164250
rect 272057 164192 272062 164248
rect 272118 164192 272246 164248
rect 272302 164192 272307 164248
rect 272057 164190 272307 164192
rect 272057 164187 272123 164190
rect 272241 164187 272307 164190
rect 301037 164250 301103 164253
rect 301221 164250 301287 164253
rect 301037 164248 301287 164250
rect 301037 164192 301042 164248
rect 301098 164192 301226 164248
rect 301282 164192 301287 164248
rect 301037 164190 301287 164192
rect 301037 164187 301103 164190
rect 301221 164187 301287 164190
rect 372797 164250 372863 164253
rect 372981 164250 373047 164253
rect 372797 164248 373047 164250
rect 372797 164192 372802 164248
rect 372858 164192 372986 164248
rect 373042 164192 373047 164248
rect 372797 164190 373047 164192
rect 372797 164187 372863 164190
rect 372981 164187 373047 164190
rect 470409 164250 470475 164253
rect 470593 164250 470659 164253
rect 470409 164248 470659 164250
rect 470409 164192 470414 164248
rect 470470 164192 470598 164248
rect 470654 164192 470659 164248
rect 470409 164190 470659 164192
rect 470409 164187 470475 164190
rect 470593 164187 470659 164190
rect 245837 164114 245903 164117
rect 245702 164112 245903 164114
rect 245702 164056 245842 164112
rect 245898 164056 245903 164112
rect 245702 164054 245903 164056
rect 245837 164051 245903 164054
rect 251173 162890 251239 162893
rect 251357 162890 251423 162893
rect 251173 162888 251423 162890
rect 251173 162832 251178 162888
rect 251234 162832 251362 162888
rect 251418 162832 251423 162888
rect 251173 162830 251423 162832
rect 251173 162827 251239 162830
rect 251357 162827 251423 162830
rect 302601 162890 302667 162893
rect 302785 162890 302851 162893
rect 302601 162888 302851 162890
rect 302601 162832 302606 162888
rect 302662 162832 302790 162888
rect 302846 162832 302851 162888
rect 302601 162830 302851 162832
rect 302601 162827 302667 162830
rect 302785 162827 302851 162830
rect 306833 162890 306899 162893
rect 307017 162890 307083 162893
rect 306833 162888 307083 162890
rect 306833 162832 306838 162888
rect 306894 162832 307022 162888
rect 307078 162832 307083 162888
rect 306833 162830 307083 162832
rect 306833 162827 306899 162830
rect 307017 162827 307083 162830
rect 583520 158402 584960 158492
rect 583342 158342 584960 158402
rect 285622 157932 285628 157996
rect 285692 157994 285698 157996
rect 295241 157994 295307 157997
rect 330477 157994 330543 157997
rect 285692 157992 295307 157994
rect 285692 157936 295246 157992
rect 295302 157936 295307 157992
rect 285692 157934 295307 157936
rect 285692 157932 285698 157934
rect 295241 157931 295307 157934
rect 325742 157992 330543 157994
rect 325742 157936 330482 157992
rect 330538 157936 330543 157992
rect 325742 157934 330543 157936
rect 277342 157660 277348 157724
rect 277412 157722 277418 157724
rect 285622 157722 285628 157724
rect 277412 157662 285628 157722
rect 277412 157660 277418 157662
rect 285622 157660 285628 157662
rect 285692 157660 285698 157724
rect 317321 157722 317387 157725
rect 325742 157722 325802 157934
rect 330477 157931 330543 157934
rect 405406 157858 405412 157860
rect 398606 157798 405412 157858
rect 317321 157720 325802 157722
rect 317321 157664 317326 157720
rect 317382 157664 325802 157720
rect 317321 157662 325802 157664
rect 330477 157722 330543 157725
rect 330477 157720 340890 157722
rect 330477 157664 330482 157720
rect 330538 157664 340890 157720
rect 330477 157662 340890 157664
rect 317321 157659 317387 157662
rect 330477 157659 330543 157662
rect 249558 157524 249564 157588
rect 249628 157586 249634 157588
rect 295241 157586 295307 157589
rect 298001 157586 298067 157589
rect 249628 157526 254042 157586
rect 249628 157524 249634 157526
rect 253982 157450 254042 157526
rect 295241 157584 298067 157586
rect 295241 157528 295246 157584
rect 295302 157528 298006 157584
rect 298062 157528 298067 157584
rect 295241 157526 298067 157528
rect 295241 157523 295307 157526
rect 298001 157523 298067 157526
rect 277342 157450 277348 157452
rect 253982 157390 277348 157450
rect 277342 157388 277348 157390
rect 277412 157388 277418 157452
rect 306281 157450 306347 157453
rect 307569 157450 307635 157453
rect 306281 157448 307635 157450
rect 306281 157392 306286 157448
rect 306342 157392 307574 157448
rect 307630 157392 307635 157448
rect 306281 157390 307635 157392
rect 306281 157387 306347 157390
rect 307569 157387 307635 157390
rect 315941 157450 316007 157453
rect 317321 157450 317387 157453
rect 315941 157448 317387 157450
rect 315941 157392 315946 157448
rect 316002 157392 317326 157448
rect 317382 157392 317387 157448
rect 315941 157390 317387 157392
rect 340830 157450 340890 157662
rect 398606 157586 398666 157798
rect 405406 157796 405412 157798
rect 405476 157796 405482 157860
rect 470550 157662 480178 157722
rect 417877 157586 417943 157589
rect 389222 157526 398666 157586
rect 408542 157584 417943 157586
rect 408542 157528 417882 157584
rect 417938 157528 417943 157584
rect 408542 157526 417943 157528
rect 389222 157450 389282 157526
rect 340830 157390 389282 157450
rect 315941 157387 316007 157390
rect 317321 157387 317387 157390
rect 405590 157388 405596 157452
rect 405660 157450 405666 157452
rect 408542 157450 408602 157526
rect 417877 157523 417943 157526
rect 418245 157586 418311 157589
rect 437197 157586 437263 157589
rect 418245 157584 427738 157586
rect 418245 157528 418250 157584
rect 418306 157528 427738 157584
rect 418245 157526 427738 157528
rect 418245 157523 418311 157526
rect 405660 157390 408602 157450
rect 427678 157450 427738 157526
rect 427862 157584 437263 157586
rect 427862 157528 437202 157584
rect 437258 157528 437263 157584
rect 427862 157526 437263 157528
rect 427862 157450 427922 157526
rect 437197 157523 437263 157526
rect 437473 157586 437539 157589
rect 456517 157586 456583 157589
rect 437473 157584 444298 157586
rect 437473 157528 437478 157584
rect 437534 157528 444298 157584
rect 437473 157526 444298 157528
rect 437473 157523 437539 157526
rect 427678 157390 427922 157450
rect 444238 157450 444298 157526
rect 447182 157584 456583 157586
rect 447182 157528 456522 157584
rect 456578 157528 456583 157584
rect 447182 157526 456583 157528
rect 447182 157450 447242 157526
rect 456517 157523 456583 157526
rect 456885 157586 456951 157589
rect 456885 157584 466378 157586
rect 456885 157528 456890 157584
rect 456946 157528 466378 157584
rect 456885 157526 466378 157528
rect 456885 157523 456951 157526
rect 444238 157390 447242 157450
rect 466318 157450 466378 157526
rect 470550 157450 470610 157662
rect 466318 157390 470610 157450
rect 480118 157450 480178 157662
rect 480302 157662 489930 157722
rect 480302 157450 480362 157662
rect 489870 157586 489930 157662
rect 499622 157662 509250 157722
rect 489870 157526 499498 157586
rect 480118 157390 480362 157450
rect 499438 157450 499498 157526
rect 499622 157450 499682 157662
rect 509190 157586 509250 157662
rect 518942 157662 528570 157722
rect 509190 157526 518818 157586
rect 499438 157390 499682 157450
rect 518758 157450 518818 157526
rect 518942 157450 519002 157662
rect 528510 157586 528570 157662
rect 538262 157662 547890 157722
rect 528510 157526 538138 157586
rect 518758 157390 519002 157450
rect 538078 157450 538138 157526
rect 538262 157450 538322 157662
rect 547830 157586 547890 157662
rect 557582 157662 567210 157722
rect 547830 157526 557458 157586
rect 538078 157390 538322 157450
rect 557398 157450 557458 157526
rect 557582 157450 557642 157662
rect 567150 157586 567210 157662
rect 583342 157586 583402 158342
rect 583520 158252 584960 158342
rect 567150 157526 576778 157586
rect 557398 157390 557642 157450
rect 576718 157450 576778 157526
rect 576902 157526 583402 157586
rect 576902 157450 576962 157526
rect 576718 157390 576962 157450
rect 405660 157388 405666 157390
rect 376937 154594 377003 154597
rect 377121 154594 377187 154597
rect 376937 154592 377187 154594
rect 376937 154536 376942 154592
rect 376998 154536 377126 154592
rect 377182 154536 377187 154592
rect 376937 154534 377187 154536
rect 376937 154531 377003 154534
rect 377121 154531 377187 154534
rect 463877 154594 463943 154597
rect 464061 154594 464127 154597
rect 463877 154592 464127 154594
rect 463877 154536 463882 154592
rect 463938 154536 464066 154592
rect 464122 154536 464127 154592
rect 463877 154534 464127 154536
rect 463877 154531 463943 154534
rect 464061 154531 464127 154534
rect 310881 153370 310947 153373
rect 310838 153368 310947 153370
rect 310838 153312 310886 153368
rect 310942 153312 310947 153368
rect 310838 153307 310947 153312
rect 310838 153237 310898 153307
rect 310789 153232 310898 153237
rect 310789 153176 310794 153232
rect 310850 153176 310898 153232
rect 310789 153174 310898 153176
rect 327257 153234 327323 153237
rect 327441 153234 327507 153237
rect 327257 153232 327507 153234
rect 327257 153176 327262 153232
rect 327318 153176 327446 153232
rect 327502 153176 327507 153232
rect 327257 153174 327507 153176
rect 310789 153171 310855 153174
rect 327257 153171 327323 153174
rect 327441 153171 327507 153174
rect -960 150786 480 150876
rect 3325 150786 3391 150789
rect -960 150784 3391 150786
rect -960 150728 3330 150784
rect 3386 150728 3391 150784
rect -960 150726 3391 150728
rect -960 150636 480 150726
rect 3325 150723 3391 150726
rect 583520 146556 584960 146796
rect 244457 145074 244523 145077
rect 244457 145072 244658 145074
rect 244457 145016 244462 145072
rect 244518 145016 244658 145072
rect 244457 145014 244658 145016
rect 244457 145011 244523 145014
rect 244457 144938 244523 144941
rect 244598 144938 244658 145014
rect 244457 144936 244658 144938
rect 244457 144880 244462 144936
rect 244518 144880 244658 144936
rect 244457 144878 244658 144880
rect 301037 144938 301103 144941
rect 301221 144938 301287 144941
rect 301037 144936 301287 144938
rect 301037 144880 301042 144936
rect 301098 144880 301226 144936
rect 301282 144880 301287 144936
rect 301037 144878 301287 144880
rect 244457 144875 244523 144878
rect 301037 144875 301103 144878
rect 301221 144875 301287 144878
rect 325877 144938 325943 144941
rect 326061 144938 326127 144941
rect 325877 144936 326127 144938
rect 325877 144880 325882 144936
rect 325938 144880 326066 144936
rect 326122 144880 326127 144936
rect 325877 144878 326127 144880
rect 325877 144875 325943 144878
rect 326061 144875 326127 144878
rect 327165 144938 327231 144941
rect 327349 144938 327415 144941
rect 327165 144936 327415 144938
rect 327165 144880 327170 144936
rect 327226 144880 327354 144936
rect 327410 144880 327415 144936
rect 327165 144878 327415 144880
rect 327165 144875 327231 144878
rect 327349 144875 327415 144878
rect 339677 144938 339743 144941
rect 339861 144938 339927 144941
rect 339677 144936 339927 144938
rect 339677 144880 339682 144936
rect 339738 144880 339866 144936
rect 339922 144880 339927 144936
rect 339677 144878 339927 144880
rect 339677 144875 339743 144878
rect 339861 144875 339927 144878
rect 341057 144938 341123 144941
rect 341241 144938 341307 144941
rect 341057 144936 341307 144938
rect 341057 144880 341062 144936
rect 341118 144880 341246 144936
rect 341302 144880 341307 144936
rect 341057 144878 341307 144880
rect 341057 144875 341123 144878
rect 341241 144875 341307 144878
rect 389357 144938 389423 144941
rect 389633 144938 389699 144941
rect 389357 144936 389699 144938
rect 389357 144880 389362 144936
rect 389418 144880 389638 144936
rect 389694 144880 389699 144936
rect 389357 144878 389699 144880
rect 389357 144875 389423 144878
rect 389633 144875 389699 144878
rect 470409 144938 470475 144941
rect 470593 144938 470659 144941
rect 470409 144936 470659 144938
rect 470409 144880 470414 144936
rect 470470 144880 470598 144936
rect 470654 144880 470659 144936
rect 470409 144878 470659 144880
rect 470409 144875 470475 144878
rect 470593 144875 470659 144878
rect 251449 143578 251515 143581
rect 251633 143578 251699 143581
rect 251449 143576 251699 143578
rect 251449 143520 251454 143576
rect 251510 143520 251638 143576
rect 251694 143520 251699 143576
rect 251449 143518 251699 143520
rect 251449 143515 251515 143518
rect 251633 143515 251699 143518
rect 302601 143578 302667 143581
rect 302785 143578 302851 143581
rect 302601 143576 302851 143578
rect 302601 143520 302606 143576
rect 302662 143520 302790 143576
rect 302846 143520 302851 143576
rect 302601 143518 302851 143520
rect 302601 143515 302667 143518
rect 302785 143515 302851 143518
rect 239121 138140 239187 138141
rect 239070 138138 239076 138140
rect 239030 138078 239076 138138
rect 239140 138136 239187 138140
rect 239182 138080 239187 138136
rect 239070 138076 239076 138078
rect 239140 138076 239187 138080
rect 239121 138075 239187 138076
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 236269 135282 236335 135285
rect 236453 135282 236519 135285
rect 239121 135284 239187 135285
rect 236269 135280 236519 135282
rect 236269 135224 236274 135280
rect 236330 135224 236458 135280
rect 236514 135224 236519 135280
rect 236269 135222 236519 135224
rect 236269 135219 236335 135222
rect 236453 135219 236519 135222
rect 239070 135220 239076 135284
rect 239140 135282 239187 135284
rect 266629 135282 266695 135285
rect 266813 135282 266879 135285
rect 239140 135280 239232 135282
rect 239182 135224 239232 135280
rect 239140 135222 239232 135224
rect 266629 135280 266879 135282
rect 266629 135224 266634 135280
rect 266690 135224 266818 135280
rect 266874 135224 266879 135280
rect 266629 135222 266879 135224
rect 239140 135220 239187 135222
rect 239121 135219 239187 135220
rect 266629 135219 266695 135222
rect 266813 135219 266879 135222
rect 341241 135282 341307 135285
rect 341425 135282 341491 135285
rect 341241 135280 341491 135282
rect 341241 135224 341246 135280
rect 341302 135224 341430 135280
rect 341486 135224 341491 135280
rect 341241 135222 341491 135224
rect 341241 135219 341307 135222
rect 341425 135219 341491 135222
rect 376937 135282 377003 135285
rect 377121 135282 377187 135285
rect 376937 135280 377187 135282
rect 376937 135224 376942 135280
rect 376998 135224 377126 135280
rect 377182 135224 377187 135280
rect 376937 135222 377187 135224
rect 376937 135219 377003 135222
rect 377121 135219 377187 135222
rect 580349 134874 580415 134877
rect 583520 134874 584960 134964
rect 580349 134872 584960 134874
rect 580349 134816 580354 134872
rect 580410 134816 584960 134872
rect 580349 134814 584960 134816
rect 580349 134811 580415 134814
rect 583520 134724 584960 134814
rect 245837 133922 245903 133925
rect 246113 133922 246179 133925
rect 245837 133920 246179 133922
rect 245837 133864 245842 133920
rect 245898 133864 246118 133920
rect 246174 133864 246179 133920
rect 245837 133862 246179 133864
rect 245837 133859 245903 133862
rect 246113 133859 246179 133862
rect 272149 133922 272215 133925
rect 272333 133922 272399 133925
rect 272149 133920 272399 133922
rect 272149 133864 272154 133920
rect 272210 133864 272338 133920
rect 272394 133864 272399 133920
rect 272149 133862 272399 133864
rect 272149 133859 272215 133862
rect 272333 133859 272399 133862
rect 362309 133922 362375 133925
rect 362493 133922 362559 133925
rect 362309 133920 362559 133922
rect 362309 133864 362314 133920
rect 362370 133864 362498 133920
rect 362554 133864 362559 133920
rect 362309 133862 362559 133864
rect 362309 133859 362375 133862
rect 362493 133859 362559 133862
rect 245929 125626 245995 125629
rect 246113 125626 246179 125629
rect 245929 125624 246179 125626
rect 245929 125568 245934 125624
rect 245990 125568 246118 125624
rect 246174 125568 246179 125624
rect 245929 125566 246179 125568
rect 245929 125563 245995 125566
rect 246113 125563 246179 125566
rect 270677 125626 270743 125629
rect 270953 125626 271019 125629
rect 270677 125624 271019 125626
rect 270677 125568 270682 125624
rect 270738 125568 270958 125624
rect 271014 125568 271019 125624
rect 270677 125566 271019 125568
rect 270677 125563 270743 125566
rect 270953 125563 271019 125566
rect 301037 125626 301103 125629
rect 301221 125626 301287 125629
rect 301037 125624 301287 125626
rect 301037 125568 301042 125624
rect 301098 125568 301226 125624
rect 301282 125568 301287 125624
rect 301037 125566 301287 125568
rect 301037 125563 301103 125566
rect 301221 125563 301287 125566
rect 327165 125626 327231 125629
rect 327349 125626 327415 125629
rect 327165 125624 327415 125626
rect 327165 125568 327170 125624
rect 327226 125568 327354 125624
rect 327410 125568 327415 125624
rect 327165 125566 327415 125568
rect 327165 125563 327231 125566
rect 327349 125563 327415 125566
rect 340873 125626 340939 125629
rect 341057 125626 341123 125629
rect 340873 125624 341123 125626
rect 340873 125568 340878 125624
rect 340934 125568 341062 125624
rect 341118 125568 341123 125624
rect 340873 125566 341123 125568
rect 340873 125563 340939 125566
rect 341057 125563 341123 125566
rect 463877 125626 463943 125629
rect 464061 125626 464127 125629
rect 463877 125624 464127 125626
rect 463877 125568 463882 125624
rect 463938 125568 464066 125624
rect 464122 125568 464127 125624
rect 463877 125566 464127 125568
rect 463877 125563 463943 125566
rect 464061 125563 464127 125566
rect 470409 125626 470475 125629
rect 470593 125626 470659 125629
rect 470409 125624 470659 125626
rect 470409 125568 470414 125624
rect 470470 125568 470598 125624
rect 470654 125568 470659 125624
rect 470409 125566 470659 125568
rect 470409 125563 470475 125566
rect 470593 125563 470659 125566
rect 285949 124130 286015 124133
rect 285814 124128 286015 124130
rect 285814 124072 285954 124128
rect 286010 124072 286015 124128
rect 285814 124070 286015 124072
rect 285814 123994 285874 124070
rect 285949 124067 286015 124070
rect 286225 123994 286291 123997
rect 285814 123992 286291 123994
rect 285814 123936 286230 123992
rect 286286 123936 286291 123992
rect 285814 123934 286291 123936
rect 286225 123931 286291 123934
rect 580257 123178 580323 123181
rect 583520 123178 584960 123268
rect 580257 123176 584960 123178
rect 580257 123120 580262 123176
rect 580318 123120 584960 123176
rect 580257 123118 584960 123120
rect 580257 123115 580323 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 389265 118826 389331 118829
rect 389398 118826 389404 118828
rect 389265 118824 389404 118826
rect 389265 118768 389270 118824
rect 389326 118768 389404 118824
rect 389265 118766 389404 118768
rect 389265 118763 389331 118766
rect 389398 118764 389404 118766
rect 389468 118764 389474 118828
rect 236269 115970 236335 115973
rect 236453 115970 236519 115973
rect 236269 115968 236519 115970
rect 236269 115912 236274 115968
rect 236330 115912 236458 115968
rect 236514 115912 236519 115968
rect 236269 115910 236519 115912
rect 236269 115907 236335 115910
rect 236453 115907 236519 115910
rect 239121 115970 239187 115973
rect 239305 115970 239371 115973
rect 239121 115968 239371 115970
rect 239121 115912 239126 115968
rect 239182 115912 239310 115968
rect 239366 115912 239371 115968
rect 239121 115910 239371 115912
rect 239121 115907 239187 115910
rect 239305 115907 239371 115910
rect 266629 115970 266695 115973
rect 266813 115970 266879 115973
rect 266629 115968 266879 115970
rect 266629 115912 266634 115968
rect 266690 115912 266818 115968
rect 266874 115912 266879 115968
rect 266629 115910 266879 115912
rect 266629 115907 266695 115910
rect 266813 115907 266879 115910
rect 583520 111482 584960 111572
rect 583342 111422 584960 111482
rect 473302 111012 473308 111076
rect 473372 111074 473378 111076
rect 482921 111074 482987 111077
rect 473372 111072 482987 111074
rect 473372 111016 482926 111072
rect 482982 111016 482987 111072
rect 473372 111014 482987 111016
rect 473372 111012 473378 111014
rect 482921 111011 482987 111014
rect 307702 110876 307708 110940
rect 307772 110938 307778 110940
rect 405406 110938 405412 110940
rect 307772 110878 312002 110938
rect 307772 110876 307778 110878
rect 244038 110740 244044 110804
rect 244108 110802 244114 110804
rect 278773 110802 278839 110805
rect 244108 110742 254042 110802
rect 244108 110740 244114 110742
rect 253982 110666 254042 110742
rect 278773 110800 288266 110802
rect 278773 110744 278778 110800
rect 278834 110744 288266 110800
rect 278773 110742 288266 110744
rect 278773 110739 278839 110742
rect 278773 110666 278839 110669
rect 253982 110664 278839 110666
rect 253982 110608 278778 110664
rect 278834 110608 278839 110664
rect 253982 110606 278839 110608
rect 288206 110666 288266 110742
rect 307518 110666 307524 110668
rect 288206 110606 307524 110666
rect 278773 110603 278839 110606
rect 307518 110604 307524 110606
rect 307588 110604 307594 110668
rect 311942 110666 312002 110878
rect 398606 110878 405412 110938
rect 328269 110802 328335 110805
rect 317278 110800 328335 110802
rect 317278 110744 328274 110800
rect 328330 110744 328335 110800
rect 317278 110742 328335 110744
rect 317278 110666 317338 110742
rect 328269 110739 328335 110742
rect 328453 110802 328519 110805
rect 357341 110802 357407 110805
rect 376661 110802 376727 110805
rect 328453 110800 340890 110802
rect 328453 110744 328458 110800
rect 328514 110744 340890 110800
rect 328453 110742 340890 110744
rect 328453 110739 328519 110742
rect 311942 110606 317338 110666
rect 340830 110530 340890 110742
rect 357341 110800 360210 110802
rect 357341 110744 357346 110800
rect 357402 110744 360210 110800
rect 357341 110742 360210 110744
rect 357341 110739 357407 110742
rect 347773 110530 347839 110533
rect 340830 110528 347839 110530
rect 340830 110472 347778 110528
rect 347834 110472 347839 110528
rect 340830 110470 347839 110472
rect 360150 110530 360210 110742
rect 376661 110800 379530 110802
rect 376661 110744 376666 110800
rect 376722 110744 379530 110800
rect 376661 110742 379530 110744
rect 376661 110739 376727 110742
rect 368197 110530 368263 110533
rect 360150 110528 368263 110530
rect 360150 110472 368202 110528
rect 368258 110472 368263 110528
rect 360150 110470 368263 110472
rect 379470 110530 379530 110742
rect 398606 110666 398666 110878
rect 405406 110876 405412 110878
rect 405476 110876 405482 110940
rect 487797 110938 487863 110941
rect 483062 110936 487863 110938
rect 483062 110880 487802 110936
rect 487858 110880 487863 110936
rect 483062 110878 487863 110880
rect 473302 110802 473308 110804
rect 466502 110742 473308 110802
rect 414013 110666 414079 110669
rect 437197 110666 437263 110669
rect 389222 110606 398666 110666
rect 408542 110664 414079 110666
rect 408542 110608 414018 110664
rect 414074 110608 414079 110664
rect 408542 110606 414079 110608
rect 389222 110530 389282 110606
rect 379470 110470 389282 110530
rect 347773 110467 347839 110470
rect 368197 110467 368263 110470
rect 405590 110468 405596 110532
rect 405660 110530 405666 110532
rect 408542 110530 408602 110606
rect 414013 110603 414079 110606
rect 427862 110664 437263 110666
rect 427862 110608 437202 110664
rect 437258 110608 437263 110664
rect 427862 110606 437263 110608
rect 405660 110470 408602 110530
rect 423489 110530 423555 110533
rect 427862 110530 427922 110606
rect 437197 110603 437263 110606
rect 437473 110666 437539 110669
rect 456517 110666 456583 110669
rect 437473 110664 444298 110666
rect 437473 110608 437478 110664
rect 437534 110608 444298 110664
rect 437473 110606 444298 110608
rect 437473 110603 437539 110606
rect 423489 110528 427922 110530
rect 423489 110472 423494 110528
rect 423550 110472 427922 110528
rect 423489 110470 427922 110472
rect 444238 110530 444298 110606
rect 447182 110664 456583 110666
rect 447182 110608 456522 110664
rect 456578 110608 456583 110664
rect 447182 110606 456583 110608
rect 447182 110530 447242 110606
rect 456517 110603 456583 110606
rect 458817 110666 458883 110669
rect 458817 110664 463618 110666
rect 458817 110608 458822 110664
rect 458878 110608 463618 110664
rect 458817 110606 463618 110608
rect 458817 110603 458883 110606
rect 444238 110470 447242 110530
rect 463558 110530 463618 110606
rect 466502 110530 466562 110742
rect 473302 110740 473308 110742
rect 473372 110740 473378 110804
rect 482921 110666 482987 110669
rect 483062 110666 483122 110878
rect 487797 110875 487863 110878
rect 492622 110740 492628 110804
rect 492692 110802 492698 110804
rect 492692 110742 509250 110802
rect 492692 110740 492698 110742
rect 482921 110664 483122 110666
rect 482921 110608 482926 110664
rect 482982 110608 483122 110664
rect 482921 110606 483122 110608
rect 509190 110666 509250 110742
rect 518942 110742 528570 110802
rect 509190 110606 518818 110666
rect 482921 110603 482987 110606
rect 463558 110470 466562 110530
rect 487797 110530 487863 110533
rect 492622 110530 492628 110532
rect 487797 110528 492628 110530
rect 487797 110472 487802 110528
rect 487858 110472 492628 110528
rect 487797 110470 492628 110472
rect 405660 110468 405666 110470
rect 423489 110467 423555 110470
rect 487797 110467 487863 110470
rect 492622 110468 492628 110470
rect 492692 110468 492698 110532
rect 518758 110530 518818 110606
rect 518942 110530 519002 110742
rect 528510 110666 528570 110742
rect 538262 110742 547890 110802
rect 528510 110606 538138 110666
rect 518758 110470 519002 110530
rect 538078 110530 538138 110606
rect 538262 110530 538322 110742
rect 547830 110666 547890 110742
rect 557582 110742 567210 110802
rect 547830 110606 557458 110666
rect 538078 110470 538322 110530
rect 557398 110530 557458 110606
rect 557582 110530 557642 110742
rect 567150 110666 567210 110742
rect 583342 110666 583402 111422
rect 583520 111332 584960 111422
rect 567150 110606 576778 110666
rect 557398 110470 557642 110530
rect 576718 110530 576778 110606
rect 576902 110606 583402 110666
rect 576902 110530 576962 110606
rect 576718 110470 576962 110530
rect 389449 108900 389515 108901
rect 389398 108898 389404 108900
rect 389358 108838 389404 108898
rect 389468 108896 389515 108900
rect 389510 108840 389515 108896
rect 389398 108836 389404 108838
rect 389468 108836 389515 108840
rect 389449 108835 389515 108836
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 341241 106314 341307 106317
rect 341425 106314 341491 106317
rect 341241 106312 341491 106314
rect 341241 106256 341246 106312
rect 341302 106256 341430 106312
rect 341486 106256 341491 106312
rect 341241 106254 341491 106256
rect 341241 106251 341307 106254
rect 341425 106251 341491 106254
rect 366817 106314 366883 106317
rect 367001 106314 367067 106317
rect 366817 106312 367067 106314
rect 366817 106256 366822 106312
rect 366878 106256 367006 106312
rect 367062 106256 367067 106312
rect 366817 106254 367067 106256
rect 366817 106251 366883 106254
rect 367001 106251 367067 106254
rect 290089 102098 290155 102101
rect 290089 102096 290290 102098
rect 290089 102040 290094 102096
rect 290150 102040 290290 102096
rect 290089 102038 290290 102040
rect 290089 102035 290155 102038
rect 289905 101962 289971 101965
rect 290230 101962 290290 102038
rect 289905 101960 290290 101962
rect 289905 101904 289910 101960
rect 289966 101904 290290 101960
rect 289905 101902 290290 101904
rect 289905 101899 289971 101902
rect 583520 99636 584960 99876
rect 367001 96932 367067 96933
rect 366950 96930 366956 96932
rect 366910 96870 366956 96930
rect 367020 96928 367067 96932
rect 367062 96872 367067 96928
rect 366950 96868 366956 96870
rect 367020 96868 367067 96872
rect 367001 96867 367067 96868
rect 266721 96794 266787 96797
rect 266494 96792 266787 96794
rect 266494 96736 266726 96792
rect 266782 96736 266787 96792
rect 266494 96734 266787 96736
rect 236269 96658 236335 96661
rect 236637 96658 236703 96661
rect 236269 96656 236703 96658
rect 236269 96600 236274 96656
rect 236330 96600 236642 96656
rect 236698 96600 236703 96656
rect 236269 96598 236703 96600
rect 236269 96595 236335 96598
rect 236637 96595 236703 96598
rect 239121 96658 239187 96661
rect 239305 96658 239371 96661
rect 239121 96656 239371 96658
rect 239121 96600 239126 96656
rect 239182 96600 239310 96656
rect 239366 96600 239371 96656
rect 239121 96598 239371 96600
rect 239121 96595 239187 96598
rect 239305 96595 239371 96598
rect 259545 96658 259611 96661
rect 259729 96658 259795 96661
rect 259545 96656 259795 96658
rect 259545 96600 259550 96656
rect 259606 96600 259734 96656
rect 259790 96600 259795 96656
rect 259545 96598 259795 96600
rect 266494 96658 266554 96734
rect 266721 96731 266787 96734
rect 266629 96658 266695 96661
rect 367001 96660 367067 96661
rect 366950 96658 366956 96660
rect 266494 96656 266695 96658
rect 266494 96600 266634 96656
rect 266690 96600 266695 96656
rect 266494 96598 266695 96600
rect 366910 96598 366956 96658
rect 367020 96656 367067 96660
rect 367062 96600 367067 96656
rect 259545 96595 259611 96598
rect 259729 96595 259795 96598
rect 266629 96595 266695 96598
rect 366950 96596 366956 96598
rect 367020 96596 367067 96600
rect 367001 96595 367067 96596
rect 360469 95298 360535 95301
rect 360334 95296 360535 95298
rect 360334 95240 360474 95296
rect 360530 95240 360535 95296
rect 360334 95238 360535 95240
rect 360334 95165 360394 95238
rect 360469 95235 360535 95238
rect 360334 95160 360443 95165
rect 360334 95104 360382 95160
rect 360438 95104 360443 95160
rect 360334 95102 360443 95104
rect 360377 95099 360443 95102
rect 296805 93802 296871 93805
rect 296670 93800 296871 93802
rect 296670 93744 296810 93800
rect 296866 93744 296871 93800
rect 296670 93742 296871 93744
rect 296670 93666 296730 93742
rect 296805 93739 296871 93742
rect 297173 93666 297239 93669
rect 296670 93664 297239 93666
rect 296670 93608 297178 93664
rect 297234 93608 297239 93664
rect 296670 93606 297239 93608
rect 297173 93603 297239 93606
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 241462 87484 241468 87548
rect 241532 87546 241538 87548
rect 251081 87546 251147 87549
rect 241532 87544 251147 87546
rect 241532 87488 251086 87544
rect 251142 87488 251147 87544
rect 241532 87486 251147 87488
rect 241532 87484 241538 87486
rect 251081 87483 251147 87486
rect 396022 87484 396028 87548
rect 396092 87546 396098 87548
rect 405590 87546 405596 87548
rect 396092 87486 405596 87546
rect 396092 87484 396098 87486
rect 405590 87484 405596 87486
rect 405660 87484 405666 87548
rect 260782 87348 260788 87412
rect 260852 87410 260858 87412
rect 277342 87410 277348 87412
rect 260852 87350 277348 87410
rect 260852 87348 260858 87350
rect 277342 87348 277348 87350
rect 277412 87348 277418 87412
rect 308998 87350 317338 87410
rect 251081 87274 251147 87277
rect 251214 87274 251220 87276
rect 251081 87272 251220 87274
rect 251081 87216 251086 87272
rect 251142 87216 251220 87272
rect 251081 87214 251220 87216
rect 251081 87211 251147 87214
rect 251214 87212 251220 87214
rect 251284 87212 251290 87276
rect 251173 87140 251239 87141
rect 239990 87076 239996 87140
rect 240060 87138 240066 87140
rect 241462 87138 241468 87140
rect 240060 87078 241468 87138
rect 240060 87076 240066 87078
rect 241462 87076 241468 87078
rect 241532 87076 241538 87140
rect 251173 87136 251220 87140
rect 251284 87138 251290 87140
rect 260649 87138 260715 87141
rect 260782 87138 260788 87140
rect 251173 87080 251178 87136
rect 251173 87076 251220 87080
rect 251284 87078 251330 87138
rect 260649 87136 260788 87138
rect 260649 87080 260654 87136
rect 260710 87080 260788 87136
rect 260649 87078 260788 87080
rect 251284 87076 251290 87078
rect 251173 87075 251239 87076
rect 260649 87075 260715 87078
rect 260782 87076 260788 87078
rect 260852 87076 260858 87140
rect 277342 87076 277348 87140
rect 277412 87138 277418 87140
rect 283465 87138 283531 87141
rect 277412 87136 283531 87138
rect 277412 87080 283470 87136
rect 283526 87080 283531 87136
rect 277412 87078 283531 87080
rect 277412 87076 277418 87078
rect 283465 87075 283531 87078
rect 283649 87138 283715 87141
rect 297541 87138 297607 87141
rect 283649 87136 297607 87138
rect 283649 87080 283654 87136
rect 283710 87080 297546 87136
rect 297602 87080 297607 87136
rect 283649 87078 297607 87080
rect 283649 87075 283715 87078
rect 297541 87075 297607 87078
rect 306281 87002 306347 87005
rect 308998 87002 309058 87350
rect 317278 87274 317338 87350
rect 481582 87348 481588 87412
rect 481652 87410 481658 87412
rect 491201 87410 491267 87413
rect 481652 87408 491267 87410
rect 481652 87352 491206 87408
rect 491262 87352 491267 87408
rect 481652 87350 491267 87352
rect 481652 87348 481658 87350
rect 491201 87347 491267 87350
rect 357341 87274 357407 87277
rect 476021 87274 476087 87277
rect 317278 87214 340706 87274
rect 340646 87138 340706 87214
rect 357341 87272 360210 87274
rect 357341 87216 357346 87272
rect 357402 87216 360210 87272
rect 357341 87214 360210 87216
rect 357341 87211 357407 87214
rect 346301 87138 346367 87141
rect 340646 87136 346367 87138
rect 340646 87080 346306 87136
rect 346362 87080 346367 87136
rect 340646 87078 346367 87080
rect 346301 87075 346367 87078
rect 306281 87000 309058 87002
rect 306281 86944 306286 87000
rect 306342 86944 309058 87000
rect 306281 86942 309058 86944
rect 346301 87002 346367 87005
rect 347773 87002 347839 87005
rect 346301 87000 347839 87002
rect 346301 86944 346306 87000
rect 346362 86944 347778 87000
rect 347834 86944 347839 87000
rect 346301 86942 347839 86944
rect 360150 87002 360210 87214
rect 466502 87272 476087 87274
rect 466502 87216 476026 87272
rect 476082 87216 476087 87272
rect 466502 87214 476087 87216
rect 376753 87138 376819 87141
rect 369902 87136 376819 87138
rect 369902 87080 376758 87136
rect 376814 87080 376819 87136
rect 369902 87078 376819 87080
rect 369902 87002 369962 87078
rect 376753 87075 376819 87078
rect 395981 87140 396047 87141
rect 395981 87136 396028 87140
rect 396092 87138 396098 87140
rect 437197 87138 437263 87141
rect 395981 87080 395986 87136
rect 395981 87076 396028 87080
rect 396092 87078 396174 87138
rect 408542 87078 424978 87138
rect 396092 87076 396098 87078
rect 395981 87075 396047 87076
rect 360150 86942 369962 87002
rect 386229 87002 386295 87005
rect 386413 87002 386479 87005
rect 386229 87000 386479 87002
rect 386229 86944 386234 87000
rect 386290 86944 386418 87000
rect 386474 86944 386479 87000
rect 386229 86942 386479 86944
rect 306281 86939 306347 86942
rect 346301 86939 346367 86942
rect 347773 86939 347839 86942
rect 386229 86939 386295 86942
rect 386413 86939 386479 86942
rect 405590 86940 405596 87004
rect 405660 87002 405666 87004
rect 408542 87002 408602 87078
rect 405660 86942 408602 87002
rect 424918 87002 424978 87078
rect 427862 87136 437263 87138
rect 427862 87080 437202 87136
rect 437258 87080 437263 87136
rect 427862 87078 437263 87080
rect 427862 87002 427922 87078
rect 437197 87075 437263 87078
rect 437473 87138 437539 87141
rect 456517 87138 456583 87141
rect 437473 87136 444298 87138
rect 437473 87080 437478 87136
rect 437534 87080 444298 87136
rect 437473 87078 444298 87080
rect 437473 87075 437539 87078
rect 424918 86942 427922 87002
rect 444238 87002 444298 87078
rect 447182 87136 456583 87138
rect 447182 87080 456522 87136
rect 456578 87080 456583 87136
rect 447182 87078 456583 87080
rect 447182 87002 447242 87078
rect 456517 87075 456583 87078
rect 456977 87138 457043 87141
rect 456977 87136 463618 87138
rect 456977 87080 456982 87136
rect 457038 87080 463618 87136
rect 456977 87078 463618 87080
rect 456977 87075 457043 87078
rect 444238 86942 447242 87002
rect 463558 87002 463618 87078
rect 466502 87002 466562 87214
rect 476021 87211 476087 87214
rect 502241 87274 502307 87277
rect 502241 87272 509250 87274
rect 502241 87216 502246 87272
rect 502302 87216 509250 87272
rect 502241 87214 509250 87216
rect 502241 87211 502307 87214
rect 476205 87138 476271 87141
rect 481582 87138 481588 87140
rect 476205 87136 481588 87138
rect 476205 87080 476210 87136
rect 476266 87080 481588 87136
rect 476205 87078 481588 87080
rect 476205 87075 476271 87078
rect 481582 87076 481588 87078
rect 481652 87076 481658 87140
rect 509190 87138 509250 87214
rect 518942 87214 528570 87274
rect 509190 87078 518818 87138
rect 463558 86942 466562 87002
rect 491201 87002 491267 87005
rect 494605 87002 494671 87005
rect 491201 87000 494671 87002
rect 491201 86944 491206 87000
rect 491262 86944 494610 87000
rect 494666 86944 494671 87000
rect 491201 86942 494671 86944
rect 518758 87002 518818 87078
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 538262 87214 547890 87274
rect 528510 87078 538138 87138
rect 518758 86942 519002 87002
rect 538078 87002 538138 87078
rect 538262 87002 538322 87214
rect 547830 87138 547890 87214
rect 557582 87214 567210 87274
rect 547830 87078 557458 87138
rect 538078 86942 538322 87002
rect 557398 87002 557458 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 557398 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 405660 86940 405666 86942
rect 491201 86939 491267 86942
rect 494605 86939 494671 86942
rect 358629 85642 358695 85645
rect 358629 85640 358922 85642
rect 358629 85584 358634 85640
rect 358690 85584 358922 85640
rect 358629 85582 358922 85584
rect 358629 85579 358695 85582
rect 358862 85370 358922 85582
rect 358997 85370 359063 85373
rect 358862 85368 359063 85370
rect 358862 85312 359002 85368
rect 359058 85312 359063 85368
rect 358862 85310 359063 85312
rect 358997 85307 359063 85310
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 386413 76530 386479 76533
rect 395838 76530 395844 76532
rect 386413 76528 395844 76530
rect 386413 76472 386418 76528
rect 386474 76472 395844 76528
rect 386413 76470 395844 76472
rect 386413 76467 386479 76470
rect 395838 76468 395844 76470
rect 395908 76468 395914 76532
rect 473302 76468 473308 76532
rect 473372 76530 473378 76532
rect 482921 76530 482987 76533
rect 473372 76528 482987 76530
rect 473372 76472 482926 76528
rect 482982 76472 482987 76528
rect 473372 76470 482987 76472
rect 473372 76468 473378 76470
rect 482921 76467 482987 76470
rect 487797 76394 487863 76397
rect 483062 76392 487863 76394
rect 483062 76336 487802 76392
rect 487858 76336 487863 76392
rect 483062 76334 487863 76336
rect 269062 76196 269068 76260
rect 269132 76258 269138 76260
rect 296529 76258 296595 76261
rect 269132 76256 296595 76258
rect 269132 76200 296534 76256
rect 296590 76200 296595 76256
rect 269132 76198 296595 76200
rect 269132 76196 269138 76198
rect 296529 76195 296595 76198
rect 327022 76196 327028 76260
rect 327092 76258 327098 76260
rect 376661 76258 376727 76261
rect 386413 76258 386479 76261
rect 473302 76258 473308 76260
rect 327092 76198 340890 76258
rect 327092 76196 327098 76198
rect 251081 76122 251147 76125
rect 251081 76120 254042 76122
rect 251081 76064 251086 76120
rect 251142 76064 254042 76120
rect 251081 76062 254042 76064
rect 251081 76059 251147 76062
rect 241094 75924 241100 75988
rect 241164 75986 241170 75988
rect 241462 75986 241468 75988
rect 241164 75926 241468 75986
rect 241164 75924 241170 75926
rect 241462 75924 241468 75926
rect 241532 75924 241538 75988
rect 253982 75986 254042 76062
rect 269062 75986 269068 75988
rect 253982 75926 269068 75986
rect 269062 75924 269068 75926
rect 269132 75924 269138 75988
rect 306373 75986 306439 75989
rect 301454 75984 306439 75986
rect 301454 75928 306378 75984
rect 306434 75928 306439 75984
rect 301454 75926 306439 75928
rect 296529 75850 296595 75853
rect 301454 75850 301514 75926
rect 306373 75923 306439 75926
rect 311249 75986 311315 75989
rect 327022 75986 327028 75988
rect 311249 75984 327028 75986
rect 311249 75928 311254 75984
rect 311310 75928 327028 75984
rect 311249 75926 327028 75928
rect 311249 75923 311315 75926
rect 327022 75924 327028 75926
rect 327092 75924 327098 75988
rect 340830 75986 340890 76198
rect 376661 76256 386479 76258
rect 376661 76200 376666 76256
rect 376722 76200 386418 76256
rect 386474 76200 386479 76256
rect 376661 76198 386479 76200
rect 376661 76195 376727 76198
rect 386413 76195 386479 76198
rect 466502 76198 473308 76258
rect 367093 76122 367159 76125
rect 350582 76120 367159 76122
rect 350582 76064 367098 76120
rect 367154 76064 367159 76120
rect 350582 76062 367159 76064
rect 350582 75986 350642 76062
rect 367093 76059 367159 76062
rect 395838 76060 395844 76124
rect 395908 76122 395914 76124
rect 396073 76122 396139 76125
rect 395908 76120 396139 76122
rect 395908 76064 396078 76120
rect 396134 76064 396139 76120
rect 395908 76062 396139 76064
rect 395908 76060 395914 76062
rect 396073 76059 396139 76062
rect 399385 76122 399451 76125
rect 437197 76122 437263 76125
rect 399385 76120 405658 76122
rect 399385 76064 399390 76120
rect 399446 76064 405658 76120
rect 399385 76062 405658 76064
rect 399385 76059 399451 76062
rect 340830 75926 350642 75986
rect 405598 75986 405658 76062
rect 408542 76062 427738 76122
rect 408542 75986 408602 76062
rect 405598 75926 408602 75986
rect 427678 75986 427738 76062
rect 427862 76120 437263 76122
rect 427862 76064 437202 76120
rect 437258 76064 437263 76120
rect 427862 76062 437263 76064
rect 427862 75986 427922 76062
rect 437197 76059 437263 76062
rect 437473 76122 437539 76125
rect 456517 76122 456583 76125
rect 437473 76120 444298 76122
rect 437473 76064 437478 76120
rect 437534 76064 444298 76120
rect 437473 76062 444298 76064
rect 437473 76059 437539 76062
rect 427678 75926 427922 75986
rect 444238 75986 444298 76062
rect 447182 76120 456583 76122
rect 447182 76064 456522 76120
rect 456578 76064 456583 76120
rect 447182 76062 456583 76064
rect 447182 75986 447242 76062
rect 456517 76059 456583 76062
rect 456793 76122 456859 76125
rect 456793 76120 463618 76122
rect 456793 76064 456798 76120
rect 456854 76064 463618 76120
rect 456793 76062 463618 76064
rect 456793 76059 456859 76062
rect 444238 75926 447242 75986
rect 463558 75986 463618 76062
rect 466502 75986 466562 76198
rect 473302 76196 473308 76198
rect 473372 76196 473378 76260
rect 482921 76122 482987 76125
rect 483062 76122 483122 76334
rect 487797 76331 487863 76334
rect 492622 76196 492628 76260
rect 492692 76258 492698 76260
rect 583520 76258 584960 76348
rect 492692 76198 509250 76258
rect 492692 76196 492698 76198
rect 482921 76120 483122 76122
rect 482921 76064 482926 76120
rect 482982 76064 483122 76120
rect 482921 76062 483122 76064
rect 509190 76122 509250 76198
rect 518942 76198 528570 76258
rect 509190 76062 518818 76122
rect 482921 76059 482987 76062
rect 463558 75926 466562 75986
rect 487797 75986 487863 75989
rect 492622 75986 492628 75988
rect 487797 75984 492628 75986
rect 487797 75928 487802 75984
rect 487858 75928 492628 75984
rect 487797 75926 492628 75928
rect 487797 75923 487863 75926
rect 492622 75924 492628 75926
rect 492692 75924 492698 75988
rect 518758 75986 518818 76062
rect 518942 75986 519002 76198
rect 528510 76122 528570 76198
rect 538262 76198 547890 76258
rect 528510 76062 538138 76122
rect 518758 75926 519002 75986
rect 538078 75986 538138 76062
rect 538262 75986 538322 76198
rect 547830 76122 547890 76198
rect 557582 76198 567210 76258
rect 547830 76062 557458 76122
rect 538078 75926 538322 75986
rect 557398 75986 557458 76062
rect 557582 75986 557642 76198
rect 567150 76122 567210 76198
rect 583342 76198 584960 76258
rect 583342 76122 583402 76198
rect 567150 76062 576778 76122
rect 557398 75926 557642 75986
rect 576718 75986 576778 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 576718 75926 576962 75986
rect 296529 75848 301514 75850
rect 296529 75792 296534 75848
rect 296590 75792 301514 75848
rect 296529 75790 301514 75792
rect 296529 75787 296595 75790
rect 241462 75652 241468 75716
rect 241532 75714 241538 75716
rect 251081 75714 251147 75717
rect 241532 75712 251147 75714
rect 241532 75656 251086 75712
rect 251142 75656 251147 75712
rect 241532 75654 251147 75656
rect 241532 75652 241538 75654
rect 251081 75651 251147 75654
rect 421005 67690 421071 67693
rect 421189 67690 421255 67693
rect 421005 67688 421255 67690
rect 421005 67632 421010 67688
rect 421066 67632 421194 67688
rect 421250 67632 421255 67688
rect 421005 67630 421255 67632
rect 421005 67627 421071 67630
rect 421189 67627 421255 67630
rect 337193 66196 337259 66197
rect 337142 66132 337148 66196
rect 337212 66194 337259 66196
rect 337212 66192 337304 66194
rect 337254 66136 337304 66192
rect 337212 66134 337304 66136
rect 337212 66132 337259 66134
rect 337193 66131 337259 66132
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect 583520 64562 584960 64652
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 583342 64502 584960 64562
rect 249742 63956 249748 64020
rect 249812 64018 249818 64020
rect 259361 64018 259427 64021
rect 405406 64018 405412 64020
rect 249812 64016 259427 64018
rect 249812 63960 259366 64016
rect 259422 63960 259427 64016
rect 249812 63958 259427 63960
rect 249812 63956 249818 63958
rect 259361 63955 259427 63958
rect 398606 63958 405412 64018
rect 275553 63882 275619 63885
rect 280102 63882 280108 63884
rect 275553 63880 280108 63882
rect 275553 63824 275558 63880
rect 275614 63824 280108 63880
rect 275553 63822 280108 63824
rect 275553 63819 275619 63822
rect 280102 63820 280108 63822
rect 280172 63820 280178 63884
rect 327022 63820 327028 63884
rect 327092 63882 327098 63884
rect 327092 63822 340890 63882
rect 327092 63820 327098 63822
rect 237230 63684 237236 63748
rect 237300 63746 237306 63748
rect 249742 63746 249748 63748
rect 237300 63686 249748 63746
rect 237300 63684 237306 63686
rect 249742 63684 249748 63686
rect 249812 63684 249818 63748
rect 285078 63686 317338 63746
rect 259361 63610 259427 63613
rect 275553 63610 275619 63613
rect 259361 63608 275619 63610
rect 259361 63552 259366 63608
rect 259422 63552 275558 63608
rect 275614 63552 275619 63608
rect 259361 63550 275619 63552
rect 259361 63547 259427 63550
rect 275553 63547 275619 63550
rect 280102 63548 280108 63612
rect 280172 63610 280178 63612
rect 285078 63610 285138 63686
rect 280172 63550 285138 63610
rect 317278 63610 317338 63686
rect 327022 63610 327028 63612
rect 317278 63550 327028 63610
rect 280172 63548 280178 63550
rect 327022 63548 327028 63550
rect 327092 63548 327098 63612
rect 340830 63610 340890 63822
rect 398606 63746 398666 63958
rect 405406 63956 405412 63958
rect 405476 63956 405482 64020
rect 470550 63822 480178 63882
rect 414013 63746 414079 63749
rect 389222 63686 398666 63746
rect 408542 63744 414079 63746
rect 408542 63688 414018 63744
rect 414074 63688 414079 63744
rect 408542 63686 414079 63688
rect 389222 63610 389282 63686
rect 340830 63550 389282 63610
rect 405590 63548 405596 63612
rect 405660 63610 405666 63612
rect 408542 63610 408602 63686
rect 414013 63683 414079 63686
rect 418889 63746 418955 63749
rect 437197 63746 437263 63749
rect 418889 63744 427738 63746
rect 418889 63688 418894 63744
rect 418950 63688 427738 63744
rect 418889 63686 427738 63688
rect 418889 63683 418955 63686
rect 405660 63550 408602 63610
rect 427678 63610 427738 63686
rect 427862 63744 437263 63746
rect 427862 63688 437202 63744
rect 437258 63688 437263 63744
rect 427862 63686 437263 63688
rect 427862 63610 427922 63686
rect 437197 63683 437263 63686
rect 437473 63746 437539 63749
rect 456517 63746 456583 63749
rect 437473 63744 444298 63746
rect 437473 63688 437478 63744
rect 437534 63688 444298 63744
rect 437473 63686 444298 63688
rect 437473 63683 437539 63686
rect 427678 63550 427922 63610
rect 444238 63610 444298 63686
rect 447182 63744 456583 63746
rect 447182 63688 456522 63744
rect 456578 63688 456583 63744
rect 447182 63686 456583 63688
rect 447182 63610 447242 63686
rect 456517 63683 456583 63686
rect 456885 63746 456951 63749
rect 456885 63744 466378 63746
rect 456885 63688 456890 63744
rect 456946 63688 466378 63744
rect 456885 63686 466378 63688
rect 456885 63683 456951 63686
rect 444238 63550 447242 63610
rect 466318 63610 466378 63686
rect 470550 63610 470610 63822
rect 466318 63550 470610 63610
rect 480118 63610 480178 63822
rect 480302 63822 489930 63882
rect 480302 63610 480362 63822
rect 489870 63746 489930 63822
rect 499622 63822 509250 63882
rect 489870 63686 499498 63746
rect 480118 63550 480362 63610
rect 499438 63610 499498 63686
rect 499622 63610 499682 63822
rect 509190 63746 509250 63822
rect 518942 63822 528570 63882
rect 509190 63686 518818 63746
rect 499438 63550 499682 63610
rect 518758 63610 518818 63686
rect 518942 63610 519002 63822
rect 528510 63746 528570 63822
rect 538262 63822 547890 63882
rect 528510 63686 538138 63746
rect 518758 63550 519002 63610
rect 538078 63610 538138 63686
rect 538262 63610 538322 63822
rect 547830 63746 547890 63822
rect 557582 63822 567210 63882
rect 547830 63686 557458 63746
rect 538078 63550 538322 63610
rect 557398 63610 557458 63686
rect 557582 63610 557642 63822
rect 567150 63746 567210 63822
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 567150 63686 576778 63746
rect 557398 63550 557642 63610
rect 576718 63610 576778 63686
rect 576902 63686 583402 63746
rect 576902 63610 576962 63686
rect 576718 63550 576962 63610
rect 405660 63548 405666 63550
rect 337142 56612 337148 56676
rect 337212 56674 337218 56676
rect 337285 56674 337351 56677
rect 337212 56672 337351 56674
rect 337212 56616 337290 56672
rect 337346 56616 337351 56672
rect 337212 56614 337351 56616
rect 337212 56612 337218 56614
rect 337285 56611 337351 56614
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 2773 50146 2839 50149
rect -960 50144 2839 50146
rect -960 50088 2778 50144
rect 2834 50088 2839 50144
rect -960 50086 2839 50088
rect -960 49996 480 50086
rect 2773 50083 2839 50086
rect 251449 48514 251515 48517
rect 251222 48512 251515 48514
rect 251222 48456 251454 48512
rect 251510 48456 251515 48512
rect 251222 48454 251515 48456
rect 245561 48378 245627 48381
rect 251222 48378 251282 48454
rect 251449 48451 251515 48454
rect 341241 48514 341307 48517
rect 341241 48512 341626 48514
rect 341241 48456 341246 48512
rect 341302 48456 341626 48512
rect 341241 48454 341626 48456
rect 341241 48451 341307 48454
rect 251357 48378 251423 48381
rect 245561 48376 245762 48378
rect 245561 48320 245566 48376
rect 245622 48320 245762 48376
rect 245561 48318 245762 48320
rect 251222 48376 251423 48378
rect 251222 48320 251362 48376
rect 251418 48320 251423 48376
rect 251222 48318 251423 48320
rect 245561 48315 245627 48318
rect 245561 48242 245627 48245
rect 245702 48242 245762 48318
rect 251357 48315 251423 48318
rect 341425 48378 341491 48381
rect 341566 48378 341626 48454
rect 341425 48376 341626 48378
rect 341425 48320 341430 48376
rect 341486 48320 341626 48376
rect 341425 48318 341626 48320
rect 341425 48315 341491 48318
rect 245561 48240 245762 48242
rect 245561 48184 245566 48240
rect 245622 48184 245762 48240
rect 245561 48182 245762 48184
rect 388989 48242 389055 48245
rect 389173 48242 389239 48245
rect 388989 48240 389239 48242
rect 388989 48184 388994 48240
rect 389050 48184 389178 48240
rect 389234 48184 389239 48240
rect 388989 48182 389239 48184
rect 245561 48179 245627 48182
rect 388989 48179 389055 48182
rect 389173 48179 389239 48182
rect 288893 44162 288959 44165
rect 289077 44162 289143 44165
rect 288893 44160 289143 44162
rect 288893 44104 288898 44160
rect 288954 44104 289082 44160
rect 289138 44104 289143 44160
rect 288893 44102 289143 44104
rect 288893 44099 288959 44102
rect 289077 44099 289143 44102
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 232998 40292 233004 40356
rect 233068 40354 233074 40356
rect 279969 40354 280035 40357
rect 233068 40294 234538 40354
rect 233068 40292 233074 40294
rect 234478 40082 234538 40294
rect 275326 40352 280035 40354
rect 275326 40296 279974 40352
rect 280030 40296 280035 40352
rect 275326 40294 280035 40296
rect 234662 40158 254042 40218
rect 234662 40082 234722 40158
rect 234478 40022 234722 40082
rect 253982 40082 254042 40158
rect 275326 40082 275386 40294
rect 279969 40291 280035 40294
rect 280153 40354 280219 40357
rect 280153 40352 283666 40354
rect 280153 40296 280158 40352
rect 280214 40296 283666 40352
rect 280153 40294 283666 40296
rect 280153 40291 280219 40294
rect 283606 40218 283666 40294
rect 327022 40292 327028 40356
rect 327092 40354 327098 40356
rect 327092 40294 340890 40354
rect 327092 40292 327098 40294
rect 306373 40218 306439 40221
rect 283606 40216 306439 40218
rect 283606 40160 306378 40216
rect 306434 40160 306439 40216
rect 283606 40158 306439 40160
rect 306373 40155 306439 40158
rect 253982 40022 275386 40082
rect 315941 40082 316007 40085
rect 327022 40082 327028 40084
rect 315941 40080 327028 40082
rect 315941 40024 315946 40080
rect 316002 40024 327028 40080
rect 315941 40022 327028 40024
rect 315941 40019 316007 40022
rect 327022 40020 327028 40022
rect 327092 40020 327098 40084
rect 340830 40082 340890 40294
rect 470550 40294 480178 40354
rect 396073 40218 396139 40221
rect 389222 40216 396139 40218
rect 389222 40160 396078 40216
rect 396134 40160 396139 40216
rect 389222 40158 396139 40160
rect 389222 40082 389282 40158
rect 396073 40155 396139 40158
rect 399017 40218 399083 40221
rect 417877 40218 417943 40221
rect 399017 40216 405658 40218
rect 399017 40160 399022 40216
rect 399078 40160 405658 40216
rect 399017 40158 405658 40160
rect 399017 40155 399083 40158
rect 340830 40022 389282 40082
rect 405598 40082 405658 40158
rect 408542 40216 417943 40218
rect 408542 40160 417882 40216
rect 417938 40160 417943 40216
rect 408542 40158 417943 40160
rect 408542 40082 408602 40158
rect 417877 40155 417943 40158
rect 418245 40218 418311 40221
rect 437197 40218 437263 40221
rect 418245 40216 427738 40218
rect 418245 40160 418250 40216
rect 418306 40160 427738 40216
rect 418245 40158 427738 40160
rect 418245 40155 418311 40158
rect 405598 40022 408602 40082
rect 427678 40082 427738 40158
rect 427862 40216 437263 40218
rect 427862 40160 437202 40216
rect 437258 40160 437263 40216
rect 427862 40158 437263 40160
rect 427862 40082 427922 40158
rect 437197 40155 437263 40158
rect 437473 40218 437539 40221
rect 456517 40218 456583 40221
rect 437473 40216 444298 40218
rect 437473 40160 437478 40216
rect 437534 40160 444298 40216
rect 437473 40158 444298 40160
rect 437473 40155 437539 40158
rect 427678 40022 427922 40082
rect 444238 40082 444298 40158
rect 447182 40216 456583 40218
rect 447182 40160 456522 40216
rect 456578 40160 456583 40216
rect 447182 40158 456583 40160
rect 447182 40082 447242 40158
rect 456517 40155 456583 40158
rect 456885 40218 456951 40221
rect 456885 40216 466378 40218
rect 456885 40160 456890 40216
rect 456946 40160 466378 40216
rect 456885 40158 466378 40160
rect 456885 40155 456951 40158
rect 444238 40022 447242 40082
rect 466318 40082 466378 40158
rect 470550 40082 470610 40294
rect 466318 40022 470610 40082
rect 480118 40082 480178 40294
rect 480302 40294 489930 40354
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect -960 35866 480 35956
rect 3141 35866 3207 35869
rect -960 35864 3207 35866
rect -960 35808 3146 35864
rect 3202 35808 3207 35864
rect -960 35806 3207 35808
rect -960 35716 480 35806
rect 3141 35803 3207 35806
rect 288382 29412 288388 29476
rect 288452 29474 288458 29476
rect 298001 29474 298067 29477
rect 405590 29474 405596 29476
rect 288452 29472 298067 29474
rect 288452 29416 298006 29472
rect 298062 29416 298067 29472
rect 288452 29414 298067 29416
rect 288452 29412 288458 29414
rect 298001 29411 298067 29414
rect 398606 29414 405596 29474
rect 257981 29338 258047 29341
rect 263409 29338 263475 29341
rect 257981 29336 263475 29338
rect 257981 29280 257986 29336
rect 258042 29280 263414 29336
rect 263470 29280 263475 29336
rect 257981 29278 263475 29280
rect 257981 29275 258047 29278
rect 263409 29275 263475 29278
rect 263593 29338 263659 29341
rect 277301 29338 277367 29341
rect 280102 29338 280108 29340
rect 263593 29336 263978 29338
rect 263593 29280 263598 29336
rect 263654 29280 263978 29336
rect 263593 29278 263978 29280
rect 263593 29275 263659 29278
rect 235758 29140 235764 29204
rect 235828 29202 235834 29204
rect 238753 29202 238819 29205
rect 235828 29200 238819 29202
rect 235828 29144 238758 29200
rect 238814 29144 238819 29200
rect 235828 29142 238819 29144
rect 263918 29202 263978 29278
rect 277301 29336 280108 29338
rect 277301 29280 277306 29336
rect 277362 29280 280108 29336
rect 277301 29278 280108 29280
rect 277301 29275 277367 29278
rect 280102 29276 280108 29278
rect 280172 29276 280178 29340
rect 317321 29338 317387 29341
rect 325734 29338 325740 29340
rect 317321 29336 325740 29338
rect 317321 29280 317326 29336
rect 317382 29280 325740 29336
rect 317321 29278 325740 29280
rect 317321 29275 317387 29278
rect 325734 29276 325740 29278
rect 325804 29276 325810 29340
rect 330477 29338 330543 29341
rect 357341 29338 357407 29341
rect 330477 29336 340890 29338
rect 330477 29280 330482 29336
rect 330538 29280 340890 29336
rect 330477 29278 340890 29280
rect 330477 29275 330543 29278
rect 267733 29202 267799 29205
rect 288382 29202 288388 29204
rect 263918 29200 267799 29202
rect 263918 29144 267738 29200
rect 267794 29144 267799 29200
rect 263918 29142 267799 29144
rect 235828 29140 235834 29142
rect 238753 29139 238819 29142
rect 267733 29139 267799 29142
rect 280294 29142 288388 29202
rect 256601 29066 256667 29069
rect 257981 29066 258047 29069
rect 256601 29064 258047 29066
rect 256601 29008 256606 29064
rect 256662 29008 257986 29064
rect 258042 29008 258047 29064
rect 256601 29006 258047 29008
rect 256601 29003 256667 29006
rect 257981 29003 258047 29006
rect 280102 29004 280108 29068
rect 280172 29066 280178 29068
rect 280294 29066 280354 29142
rect 288382 29140 288388 29142
rect 288452 29140 288458 29204
rect 298001 29202 298067 29205
rect 298001 29200 298202 29202
rect 298001 29144 298006 29200
rect 298062 29144 298202 29200
rect 298001 29142 298202 29144
rect 298001 29139 298067 29142
rect 280172 29006 280354 29066
rect 298142 29066 298202 29142
rect 302785 29066 302851 29069
rect 298142 29064 302851 29066
rect 298142 29008 302790 29064
rect 302846 29008 302851 29064
rect 298142 29006 302851 29008
rect 280172 29004 280178 29006
rect 302785 29003 302851 29006
rect 325734 29004 325740 29068
rect 325804 29066 325810 29068
rect 330477 29066 330543 29069
rect 325804 29064 330543 29066
rect 325804 29008 330482 29064
rect 330538 29008 330543 29064
rect 325804 29006 330543 29008
rect 340830 29066 340890 29278
rect 357341 29336 360210 29338
rect 357341 29280 357346 29336
rect 357402 29280 360210 29336
rect 357341 29278 360210 29280
rect 357341 29275 357407 29278
rect 347773 29066 347839 29069
rect 340830 29064 347839 29066
rect 340830 29008 347778 29064
rect 347834 29008 347839 29064
rect 340830 29006 347839 29008
rect 360150 29066 360210 29278
rect 367142 29278 379530 29338
rect 367142 29205 367202 29278
rect 367093 29200 367202 29205
rect 367093 29144 367098 29200
rect 367154 29144 367202 29200
rect 367093 29142 367202 29144
rect 367093 29139 367159 29142
rect 367093 29066 367159 29069
rect 360150 29064 367159 29066
rect 360150 29008 367098 29064
rect 367154 29008 367159 29064
rect 360150 29006 367159 29008
rect 325804 29004 325810 29006
rect 330477 29003 330543 29006
rect 347773 29003 347839 29006
rect 367093 29003 367159 29006
rect 377121 29066 377187 29069
rect 377305 29066 377371 29069
rect 377121 29064 377371 29066
rect 377121 29008 377126 29064
rect 377182 29008 377310 29064
rect 377366 29008 377371 29064
rect 377121 29006 377371 29008
rect 379470 29066 379530 29278
rect 398606 29202 398666 29414
rect 405590 29412 405596 29414
rect 405660 29412 405666 29476
rect 481582 29412 481588 29476
rect 481652 29474 481658 29476
rect 491201 29474 491267 29477
rect 481652 29472 491267 29474
rect 481652 29416 491206 29472
rect 491262 29416 491267 29472
rect 481652 29414 491267 29416
rect 481652 29412 481658 29414
rect 491201 29411 491267 29414
rect 476021 29338 476087 29341
rect 466502 29336 476087 29338
rect 466502 29280 476026 29336
rect 476082 29280 476087 29336
rect 466502 29278 476087 29280
rect 437197 29202 437263 29205
rect 389222 29142 398666 29202
rect 408542 29142 420194 29202
rect 389222 29066 389282 29142
rect 379470 29006 389282 29066
rect 377121 29003 377187 29006
rect 377305 29003 377371 29006
rect 405590 29004 405596 29068
rect 405660 29066 405666 29068
rect 408542 29066 408602 29142
rect 405660 29006 408602 29066
rect 420134 29066 420194 29142
rect 427862 29200 437263 29202
rect 427862 29144 437202 29200
rect 437258 29144 437263 29200
rect 427862 29142 437263 29144
rect 427862 29066 427922 29142
rect 437197 29139 437263 29142
rect 437473 29202 437539 29205
rect 456517 29202 456583 29205
rect 437473 29200 444298 29202
rect 437473 29144 437478 29200
rect 437534 29144 444298 29200
rect 437473 29142 444298 29144
rect 437473 29139 437539 29142
rect 420134 29006 427922 29066
rect 444238 29066 444298 29142
rect 447182 29200 456583 29202
rect 447182 29144 456522 29200
rect 456578 29144 456583 29200
rect 447182 29142 456583 29144
rect 447182 29066 447242 29142
rect 456517 29139 456583 29142
rect 456977 29202 457043 29205
rect 456977 29200 463618 29202
rect 456977 29144 456982 29200
rect 457038 29144 463618 29200
rect 456977 29142 463618 29144
rect 456977 29139 457043 29142
rect 444238 29006 447242 29066
rect 463558 29066 463618 29142
rect 466502 29066 466562 29278
rect 476021 29275 476087 29278
rect 502241 29338 502307 29341
rect 583520 29338 584960 29428
rect 502241 29336 509250 29338
rect 502241 29280 502246 29336
rect 502302 29280 509250 29336
rect 502241 29278 509250 29280
rect 502241 29275 502307 29278
rect 476205 29202 476271 29205
rect 481582 29202 481588 29204
rect 476205 29200 481588 29202
rect 476205 29144 476210 29200
rect 476266 29144 481588 29200
rect 476205 29142 481588 29144
rect 476205 29139 476271 29142
rect 481582 29140 481588 29142
rect 481652 29140 481658 29204
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 463558 29006 466562 29066
rect 491201 29066 491267 29069
rect 492765 29066 492831 29069
rect 491201 29064 492831 29066
rect 491201 29008 491206 29064
rect 491262 29008 492770 29064
rect 492826 29008 492831 29064
rect 491201 29006 492831 29008
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 405660 29004 405666 29006
rect 491201 29003 491267 29006
rect 492765 29003 492831 29006
rect 315941 28930 316007 28933
rect 317321 28930 317387 28933
rect 330109 28930 330175 28933
rect 315941 28928 317387 28930
rect 315941 28872 315946 28928
rect 316002 28872 317326 28928
rect 317382 28872 317387 28928
rect 315941 28870 317387 28872
rect 315941 28867 316007 28870
rect 317321 28867 317387 28870
rect 329974 28928 330175 28930
rect 329974 28872 330114 28928
rect 330170 28872 330175 28928
rect 329974 28870 330175 28872
rect 302785 28794 302851 28797
rect 306373 28794 306439 28797
rect 302785 28792 306439 28794
rect 302785 28736 302790 28792
rect 302846 28736 306378 28792
rect 306434 28736 306439 28792
rect 302785 28734 306439 28736
rect 329974 28794 330034 28870
rect 330109 28867 330175 28870
rect 330201 28794 330267 28797
rect 329974 28792 330267 28794
rect 329974 28736 330206 28792
rect 330262 28736 330267 28792
rect 329974 28734 330267 28736
rect 302785 28731 302851 28734
rect 306373 28731 306439 28734
rect 330201 28731 330267 28734
rect 294137 27706 294203 27709
rect 294137 27704 294338 27706
rect 294137 27648 294142 27704
rect 294198 27648 294338 27704
rect 294137 27646 294338 27648
rect 294137 27643 294203 27646
rect 294137 27570 294203 27573
rect 294278 27570 294338 27646
rect 294137 27568 294338 27570
rect 294137 27512 294142 27568
rect 294198 27512 294338 27568
rect 294137 27510 294338 27512
rect 294137 27507 294203 27510
rect 251357 26346 251423 26349
rect 251357 26344 251466 26346
rect 251357 26288 251362 26344
rect 251418 26288 251466 26344
rect 251357 26283 251466 26288
rect 251406 26210 251466 26283
rect 251633 26210 251699 26213
rect 251406 26208 251699 26210
rect 251406 26152 251638 26208
rect 251694 26152 251699 26208
rect 251406 26150 251699 26152
rect 251633 26147 251699 26150
rect 465574 21994 465580 21996
rect 614 21934 465580 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 465574 21932 465580 21934
rect 465644 21932 465650 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 231710 17308 231716 17372
rect 231780 17370 231786 17372
rect 239806 17370 239812 17372
rect 231780 17310 239812 17370
rect 231780 17308 231786 17310
rect 239806 17308 239812 17310
rect 239876 17308 239882 17372
rect 473302 17172 473308 17236
rect 473372 17234 473378 17236
rect 482921 17234 482987 17237
rect 473372 17232 482987 17234
rect 473372 17176 482926 17232
rect 482982 17176 482987 17232
rect 473372 17174 482987 17176
rect 473372 17172 473378 17174
rect 482921 17171 482987 17174
rect 298461 17098 298527 17101
rect 306373 17098 306439 17101
rect 336641 17098 336707 17101
rect 298461 17096 306439 17098
rect 298461 17040 298466 17096
rect 298522 17040 306378 17096
rect 306434 17040 306439 17096
rect 298461 17038 306439 17040
rect 298461 17035 298527 17038
rect 306373 17035 306439 17038
rect 327030 17096 336707 17098
rect 327030 17040 336646 17096
rect 336702 17040 336707 17096
rect 327030 17038 336707 17040
rect 244966 16766 254594 16826
rect 239990 16628 239996 16692
rect 240060 16690 240066 16692
rect 244966 16690 245026 16766
rect 240060 16630 245026 16690
rect 254534 16690 254594 16766
rect 260966 16764 260972 16828
rect 261036 16826 261042 16828
rect 288341 16826 288407 16829
rect 289261 16826 289327 16829
rect 327030 16826 327090 17038
rect 336641 17035 336707 17038
rect 395889 17098 395955 17101
rect 396022 17098 396028 17100
rect 395889 17096 396028 17098
rect 395889 17040 395894 17096
rect 395950 17040 396028 17096
rect 395889 17038 396028 17040
rect 395889 17035 395955 17038
rect 396022 17036 396028 17038
rect 396092 17036 396098 17100
rect 487797 17098 487863 17101
rect 483062 17096 487863 17098
rect 483062 17040 487802 17096
rect 487858 17040 487863 17096
rect 483062 17038 487863 17040
rect 347773 16962 347839 16965
rect 473302 16962 473308 16964
rect 261036 16766 273178 16826
rect 261036 16764 261042 16766
rect 260782 16690 260788 16692
rect 254534 16630 260788 16690
rect 240060 16628 240066 16630
rect 260782 16628 260788 16630
rect 260852 16628 260858 16692
rect 273118 16690 273178 16766
rect 288341 16824 289327 16826
rect 288341 16768 288346 16824
rect 288402 16768 289266 16824
rect 289322 16768 289327 16824
rect 288341 16766 289327 16768
rect 288341 16763 288407 16766
rect 289261 16763 289327 16766
rect 322246 16766 327090 16826
rect 340830 16960 347839 16962
rect 340830 16904 347778 16960
rect 347834 16904 347839 16960
rect 340830 16902 347839 16904
rect 315941 16690 316007 16693
rect 322246 16690 322306 16766
rect 273118 16630 273362 16690
rect 273302 16554 273362 16630
rect 315941 16688 322306 16690
rect 315941 16632 315946 16688
rect 316002 16632 322306 16688
rect 315941 16630 322306 16632
rect 336641 16690 336707 16693
rect 340830 16690 340890 16902
rect 347773 16899 347839 16902
rect 466502 16902 473308 16962
rect 376526 16826 376770 16860
rect 379286 16826 379714 16860
rect 385125 16826 385191 16829
rect 417877 16826 417943 16829
rect 366958 16824 385191 16826
rect 366958 16800 385130 16824
rect 366958 16766 376586 16800
rect 376710 16766 379346 16800
rect 379654 16768 385130 16800
rect 385186 16768 385191 16824
rect 379654 16766 385191 16768
rect 336641 16688 340890 16690
rect 336641 16632 336646 16688
rect 336702 16632 340890 16688
rect 336641 16630 340890 16632
rect 352649 16690 352715 16693
rect 366958 16690 367018 16766
rect 385125 16763 385191 16766
rect 408542 16824 417943 16826
rect 408542 16768 417882 16824
rect 417938 16768 417943 16824
rect 408542 16766 417943 16768
rect 352649 16688 367018 16690
rect 352649 16632 352654 16688
rect 352710 16632 367018 16688
rect 352649 16630 367018 16632
rect 315941 16627 316007 16630
rect 336641 16627 336707 16630
rect 352649 16627 352715 16630
rect 396022 16628 396028 16692
rect 396092 16690 396098 16692
rect 398741 16690 398807 16693
rect 396092 16688 398807 16690
rect 396092 16632 398746 16688
rect 398802 16632 398807 16688
rect 396092 16630 398807 16632
rect 396092 16628 396098 16630
rect 398741 16627 398807 16630
rect 398925 16690 398991 16693
rect 408542 16690 408602 16766
rect 417877 16763 417943 16766
rect 418245 16826 418311 16829
rect 437197 16826 437263 16829
rect 418245 16824 427738 16826
rect 418245 16768 418250 16824
rect 418306 16768 427738 16824
rect 418245 16766 427738 16768
rect 418245 16763 418311 16766
rect 398925 16688 408602 16690
rect 398925 16632 398930 16688
rect 398986 16632 408602 16688
rect 398925 16630 408602 16632
rect 427678 16690 427738 16766
rect 427862 16824 437263 16826
rect 427862 16768 437202 16824
rect 437258 16768 437263 16824
rect 427862 16766 437263 16768
rect 427862 16690 427922 16766
rect 437197 16763 437263 16766
rect 437473 16826 437539 16829
rect 456517 16826 456583 16829
rect 437473 16824 444298 16826
rect 437473 16768 437478 16824
rect 437534 16768 444298 16824
rect 437473 16766 444298 16768
rect 437473 16763 437539 16766
rect 427678 16630 427922 16690
rect 444238 16690 444298 16766
rect 447182 16824 456583 16826
rect 447182 16768 456522 16824
rect 456578 16768 456583 16824
rect 447182 16766 456583 16768
rect 447182 16690 447242 16766
rect 456517 16763 456583 16766
rect 458817 16826 458883 16829
rect 458817 16824 463618 16826
rect 458817 16768 458822 16824
rect 458878 16768 463618 16824
rect 458817 16766 463618 16768
rect 458817 16763 458883 16766
rect 444238 16630 447242 16690
rect 463558 16690 463618 16766
rect 466502 16690 466562 16902
rect 473302 16900 473308 16902
rect 473372 16900 473378 16964
rect 482921 16826 482987 16829
rect 483062 16826 483122 17038
rect 487797 17035 487863 17038
rect 492622 16900 492628 16964
rect 492692 16962 492698 16964
rect 492692 16902 509250 16962
rect 492692 16900 492698 16902
rect 482921 16824 483122 16826
rect 482921 16768 482926 16824
rect 482982 16768 483122 16824
rect 482921 16766 483122 16768
rect 509190 16826 509250 16902
rect 518942 16902 528570 16962
rect 509190 16766 518818 16826
rect 482921 16763 482987 16766
rect 463558 16630 466562 16690
rect 487797 16690 487863 16693
rect 492622 16690 492628 16692
rect 487797 16688 492628 16690
rect 487797 16632 487802 16688
rect 487858 16632 492628 16688
rect 487797 16630 492628 16632
rect 398925 16627 398991 16630
rect 487797 16627 487863 16630
rect 492622 16628 492628 16630
rect 492692 16628 492698 16692
rect 518758 16690 518818 16766
rect 518942 16690 519002 16902
rect 528510 16826 528570 16902
rect 538262 16902 547890 16962
rect 528510 16766 538138 16826
rect 518758 16630 519002 16690
rect 538078 16690 538138 16766
rect 538262 16690 538322 16902
rect 547830 16826 547890 16902
rect 557582 16902 567210 16962
rect 547830 16766 557458 16826
rect 538078 16630 538322 16690
rect 557398 16690 557458 16766
rect 557582 16690 557642 16902
rect 567150 16826 567210 16902
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 567150 16766 576778 16826
rect 557398 16630 557642 16690
rect 576718 16690 576778 16766
rect 576902 16766 583402 16826
rect 576902 16690 576962 16766
rect 576718 16630 576962 16690
rect 278814 16554 278820 16556
rect 273302 16494 278820 16554
rect 278814 16492 278820 16494
rect 278884 16492 278890 16556
rect 289905 16554 289971 16557
rect 298093 16554 298159 16557
rect 289905 16552 298159 16554
rect 289905 16496 289910 16552
rect 289966 16496 298098 16552
rect 298154 16496 298159 16552
rect 289905 16494 298159 16496
rect 289905 16491 289971 16494
rect 298093 16491 298159 16494
rect 307569 16554 307635 16557
rect 310789 16554 310855 16557
rect 307569 16552 310855 16554
rect 307569 16496 307574 16552
rect 307630 16496 310794 16552
rect 310850 16496 310855 16552
rect 307569 16494 310855 16496
rect 307569 16491 307635 16494
rect 310789 16491 310855 16494
rect 278814 16220 278820 16284
rect 278884 16282 278890 16284
rect 288341 16282 288407 16285
rect 278884 16280 288407 16282
rect 278884 16224 288346 16280
rect 288402 16224 288407 16280
rect 278884 16222 288407 16224
rect 278884 16220 278890 16222
rect 288341 16219 288407 16222
rect 3141 11658 3207 11661
rect 466494 11658 466500 11660
rect 3141 11656 466500 11658
rect 3141 11600 3146 11656
rect 3202 11600 466500 11656
rect 3141 11598 466500 11600
rect 3141 11595 3207 11598
rect 466494 11596 466500 11598
rect 466564 11596 466570 11660
rect 265249 9618 265315 9621
rect 265433 9618 265499 9621
rect 265249 9616 265499 9618
rect 265249 9560 265254 9616
rect 265310 9560 265438 9616
rect 265494 9560 265499 9616
rect 265249 9558 265499 9560
rect 265249 9555 265315 9558
rect 265433 9555 265499 9558
rect 132585 8938 132651 8941
rect 284477 8938 284543 8941
rect 132585 8936 284543 8938
rect 132585 8880 132590 8936
rect 132646 8880 284482 8936
rect 284538 8880 284543 8936
rect 132585 8878 284543 8880
rect 132585 8875 132651 8878
rect 284477 8875 284543 8878
rect 128997 7578 129063 7581
rect 283097 7578 283163 7581
rect 128997 7576 283163 7578
rect 128997 7520 129002 7576
rect 129058 7520 283102 7576
rect 283158 7520 283163 7576
rect 128997 7518 283163 7520
rect 128997 7515 129063 7518
rect 283097 7515 283163 7518
rect -960 7170 480 7260
rect 3141 7170 3207 7173
rect -960 7168 3207 7170
rect -960 7112 3146 7168
rect 3202 7112 3207 7168
rect -960 7110 3207 7112
rect -960 7020 480 7110
rect 3141 7107 3207 7110
rect 51625 6218 51691 6221
rect 249977 6218 250043 6221
rect 51625 6216 250043 6218
rect 51625 6160 51630 6216
rect 51686 6160 249982 6216
rect 250038 6160 250043 6216
rect 51625 6158 250043 6160
rect 51625 6155 51691 6158
rect 249977 6155 250043 6158
rect 583520 5796 584960 6036
rect 208669 4858 208735 4861
rect 314653 4858 314719 4861
rect 208669 4856 314719 4858
rect 208669 4800 208674 4856
rect 208730 4800 314658 4856
rect 314714 4800 314719 4856
rect 208669 4798 314719 4800
rect 208669 4795 208735 4798
rect 314653 4795 314719 4798
rect 467741 4858 467807 4861
rect 576209 4858 576275 4861
rect 467741 4856 576275 4858
rect 467741 4800 467746 4856
rect 467802 4800 576214 4856
rect 576270 4800 576275 4856
rect 467741 4798 576275 4800
rect 467741 4795 467807 4798
rect 576209 4795 576275 4798
rect 460105 3770 460171 3773
rect 463509 3770 463575 3773
rect 460105 3768 463575 3770
rect 460105 3712 460110 3768
rect 460166 3712 463514 3768
rect 463570 3712 463575 3768
rect 460105 3710 463575 3712
rect 460105 3707 460171 3710
rect 463509 3707 463575 3710
rect 421373 3498 421439 3501
rect 421557 3498 421623 3501
rect 421373 3496 421623 3498
rect 421373 3440 421378 3496
rect 421434 3440 421562 3496
rect 421618 3440 421623 3496
rect 421373 3438 421623 3440
rect 421373 3435 421439 3438
rect 421557 3435 421623 3438
rect 6453 3362 6519 3365
rect 232037 3362 232103 3365
rect 6453 3360 232103 3362
rect 6453 3304 6458 3360
rect 6514 3304 232042 3360
rect 232098 3304 232103 3360
rect 6453 3302 232103 3304
rect 6453 3299 6519 3302
rect 232037 3299 232103 3302
rect 307385 3362 307451 3365
rect 356237 3362 356303 3365
rect 307385 3360 356303 3362
rect 307385 3304 307390 3360
rect 307446 3304 356242 3360
rect 356298 3304 356303 3360
rect 307385 3302 356303 3304
rect 307385 3299 307451 3302
rect 356237 3299 356303 3302
rect 468753 3362 468819 3365
rect 580993 3362 581059 3365
rect 468753 3360 581059 3362
rect 468753 3304 468758 3360
rect 468814 3304 580998 3360
rect 581054 3304 581059 3360
rect 468753 3302 581059 3304
rect 468753 3299 468819 3302
rect 580993 3299 581059 3302
<< via3 >>
rect 465948 583340 466012 583404
rect 465764 583204 465828 583268
rect 242756 583068 242820 583132
rect 239260 582932 239324 582996
rect 465580 579668 465644 579732
rect 231716 579260 231780 579324
rect 233004 579320 233068 579324
rect 233004 579264 233018 579320
rect 233018 579264 233068 579320
rect 233004 579260 233068 579264
rect 235764 579260 235828 579324
rect 237236 579320 237300 579324
rect 237236 579264 237250 579320
rect 237250 579264 237300 579320
rect 237236 579260 237300 579264
rect 239996 579260 240060 579324
rect 241284 579260 241348 579324
rect 244044 579260 244108 579324
rect 249564 579320 249628 579324
rect 249564 579264 249578 579320
rect 249578 579264 249628 579320
rect 249564 579260 249628 579264
rect 466500 579320 466564 579324
rect 466500 579264 466514 579320
rect 466514 579264 466564 579320
rect 466500 579260 466564 579264
rect 465948 533020 466012 533084
rect 465764 486100 465828 486164
rect 243676 340580 243740 340644
rect 249564 340580 249628 340644
rect 242756 337996 242820 338060
rect 249564 336636 249628 336700
rect 249196 316100 249260 316164
rect 249196 312020 249260 312084
rect 249380 311748 249444 311812
rect 251404 307668 251468 307732
rect 249380 306308 249444 306372
rect 341380 299372 341444 299436
rect 251404 298148 251468 298212
rect 249196 296788 249260 296852
rect 239260 295156 239324 295220
rect 341380 289852 341444 289916
rect 341380 280060 341444 280124
rect 249196 275028 249260 275092
rect 341380 270540 341444 270604
rect 249380 267880 249444 267884
rect 249380 267824 249430 267880
rect 249430 267824 249444 267880
rect 249380 267820 249444 267824
rect 341380 260748 341444 260812
rect 249196 257952 249260 257956
rect 249196 257896 249246 257952
rect 249246 257896 249260 257952
rect 249196 257892 249260 257896
rect 341380 251228 341444 251292
rect 249012 248372 249076 248436
rect 249012 230556 249076 230620
rect 249380 230420 249444 230484
rect 249380 219268 249444 219332
rect 249748 219132 249812 219196
rect 249748 209612 249812 209676
rect 249564 200152 249628 200156
rect 249564 200096 249614 200152
rect 249614 200096 249628 200152
rect 249564 200092 249628 200096
rect 421236 196556 421300 196620
rect 249564 193156 249628 193220
rect 421236 183696 421300 183700
rect 421236 183640 421250 183696
rect 421250 183640 421300 183696
rect 421236 183636 421300 183640
rect 249012 182140 249076 182204
rect 285628 157932 285692 157996
rect 277348 157660 277412 157724
rect 285628 157660 285692 157724
rect 249564 157524 249628 157588
rect 277348 157388 277412 157452
rect 405412 157796 405476 157860
rect 405596 157388 405660 157452
rect 239076 138136 239140 138140
rect 239076 138080 239126 138136
rect 239126 138080 239140 138136
rect 239076 138076 239140 138080
rect 239076 135280 239140 135284
rect 239076 135224 239126 135280
rect 239126 135224 239140 135280
rect 239076 135220 239140 135224
rect 389404 118764 389468 118828
rect 473308 111012 473372 111076
rect 307708 110876 307772 110940
rect 244044 110740 244108 110804
rect 307524 110604 307588 110668
rect 405412 110876 405476 110940
rect 405596 110468 405660 110532
rect 473308 110740 473372 110804
rect 492628 110740 492692 110804
rect 492628 110468 492692 110532
rect 389404 108896 389468 108900
rect 389404 108840 389454 108896
rect 389454 108840 389468 108896
rect 389404 108836 389468 108840
rect 366956 96928 367020 96932
rect 366956 96872 367006 96928
rect 367006 96872 367020 96928
rect 366956 96868 367020 96872
rect 366956 96656 367020 96660
rect 366956 96600 367006 96656
rect 367006 96600 367020 96656
rect 366956 96596 367020 96600
rect 241468 87484 241532 87548
rect 396028 87484 396092 87548
rect 405596 87484 405660 87548
rect 260788 87348 260852 87412
rect 277348 87348 277412 87412
rect 251220 87212 251284 87276
rect 239996 87076 240060 87140
rect 241468 87076 241532 87140
rect 251220 87136 251284 87140
rect 251220 87080 251234 87136
rect 251234 87080 251284 87136
rect 251220 87076 251284 87080
rect 260788 87076 260852 87140
rect 277348 87076 277412 87140
rect 481588 87348 481652 87412
rect 396028 87136 396092 87140
rect 396028 87080 396042 87136
rect 396042 87080 396092 87136
rect 396028 87076 396092 87080
rect 405596 86940 405660 87004
rect 481588 87076 481652 87140
rect 395844 76468 395908 76532
rect 473308 76468 473372 76532
rect 269068 76196 269132 76260
rect 327028 76196 327092 76260
rect 241100 75924 241164 75988
rect 241468 75924 241532 75988
rect 269068 75924 269132 75988
rect 327028 75924 327092 75988
rect 395844 76060 395908 76124
rect 473308 76196 473372 76260
rect 492628 76196 492692 76260
rect 492628 75924 492692 75988
rect 241468 75652 241532 75716
rect 337148 66192 337212 66196
rect 337148 66136 337198 66192
rect 337198 66136 337212 66192
rect 337148 66132 337212 66136
rect 249748 63956 249812 64020
rect 280108 63820 280172 63884
rect 327028 63820 327092 63884
rect 237236 63684 237300 63748
rect 249748 63684 249812 63748
rect 280108 63548 280172 63612
rect 327028 63548 327092 63612
rect 405412 63956 405476 64020
rect 405596 63548 405660 63612
rect 337148 56612 337212 56676
rect 233004 40292 233068 40356
rect 327028 40292 327092 40356
rect 327028 40020 327092 40084
rect 288388 29412 288452 29476
rect 235764 29140 235828 29204
rect 280108 29276 280172 29340
rect 325740 29276 325804 29340
rect 280108 29004 280172 29068
rect 288388 29140 288452 29204
rect 325740 29004 325804 29068
rect 405596 29412 405660 29476
rect 481588 29412 481652 29476
rect 405596 29004 405660 29068
rect 481588 29140 481652 29204
rect 465580 21932 465644 21996
rect 231716 17308 231780 17372
rect 239812 17308 239876 17372
rect 473308 17172 473372 17236
rect 239996 16628 240060 16692
rect 260972 16764 261036 16828
rect 396028 17036 396092 17100
rect 260788 16628 260852 16692
rect 396028 16628 396092 16692
rect 473308 16900 473372 16964
rect 492628 16900 492692 16964
rect 492628 16628 492692 16692
rect 278820 16492 278884 16556
rect 278820 16220 278884 16284
rect 466500 11596 466564 11660
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 231715 579324 231781 579325
rect 231715 579260 231716 579324
rect 231780 579260 231781 579324
rect 231715 579259 231781 579260
rect 233003 579324 233069 579325
rect 233003 579260 233004 579324
rect 233068 579260 233069 579324
rect 233003 579259 233069 579260
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 17373 231778 579259
rect 233006 40357 233066 579259
rect 234804 560454 235404 595898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 235763 579324 235829 579325
rect 235763 579260 235764 579324
rect 235828 579260 235829 579324
rect 235763 579259 235829 579260
rect 237235 579324 237301 579325
rect 237235 579260 237236 579324
rect 237300 579260 237301 579324
rect 237235 579259 237301 579260
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 233003 40356 233069 40357
rect 233003 40292 233004 40356
rect 233068 40292 233069 40356
rect 233003 40291 233069 40292
rect 234804 20454 235404 55898
rect 235766 29205 235826 579259
rect 237238 63749 237298 579259
rect 238404 564054 239004 599498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 239259 582996 239325 582997
rect 239259 582932 239260 582996
rect 239324 582932 239325 582996
rect 239259 582931 239325 582932
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 239262 295221 239322 582931
rect 239995 579324 240061 579325
rect 239995 579260 239996 579324
rect 240060 579260 240061 579324
rect 239995 579259 240061 579260
rect 241283 579324 241349 579325
rect 241283 579260 241284 579324
rect 241348 579260 241349 579324
rect 241283 579259 241349 579260
rect 239259 295220 239325 295221
rect 239259 295156 239260 295220
rect 239324 295156 239325 295220
rect 239259 295155 239325 295156
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 239075 138140 239141 138141
rect 239075 138076 239076 138140
rect 239140 138076 239141 138140
rect 239075 138075 239141 138076
rect 239078 135285 239138 138075
rect 239075 135284 239141 135285
rect 239075 135220 239076 135284
rect 239140 135220 239141 135284
rect 239075 135219 239141 135220
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 237235 63748 237301 63749
rect 237235 63684 237236 63748
rect 237300 63684 237301 63748
rect 237235 63683 237301 63684
rect 238404 60054 239004 95498
rect 239998 87141 240058 579259
rect 239995 87140 240061 87141
rect 239995 87076 239996 87140
rect 240060 87076 240061 87140
rect 239995 87075 240061 87076
rect 241286 77210 241346 579259
rect 242004 567654 242604 603098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 242755 583132 242821 583133
rect 242755 583068 242756 583132
rect 242820 583068 242821 583132
rect 242755 583067 242821 583068
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242758 338061 242818 583067
rect 244043 579324 244109 579325
rect 244043 579260 244044 579324
rect 244108 579260 244109 579324
rect 244043 579259 244109 579260
rect 243678 413898 243738 432702
rect 243126 407098 243186 412982
rect 243678 397490 243738 406182
rect 243310 397430 243738 397490
rect 243310 396218 243370 397430
rect 243678 340645 243738 395982
rect 243675 340644 243741 340645
rect 243675 340580 243676 340644
rect 243740 340580 243741 340644
rect 243675 340579 243741 340580
rect 242755 338060 242821 338061
rect 242755 337996 242756 338060
rect 242820 337996 242821 338060
rect 242755 337995 242821 337996
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 244046 110805 244106 579259
rect 245604 571254 246204 606698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 249563 579324 249629 579325
rect 249563 579260 249564 579324
rect 249628 579260 249629 579324
rect 249563 579259 249629 579260
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 249566 432170 249626 579259
rect 249382 432110 249626 432170
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 249382 431578 249442 432110
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 249563 340644 249629 340645
rect 249563 340580 249564 340644
rect 249628 340580 249629 340644
rect 249563 340579 249629 340580
rect 249566 336701 249626 340579
rect 249563 336700 249629 336701
rect 249563 336636 249564 336700
rect 249628 336636 249629 336700
rect 249563 336635 249629 336636
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 249195 316164 249261 316165
rect 249195 316100 249196 316164
rect 249260 316100 249261 316164
rect 249195 316099 249261 316100
rect 249198 312085 249258 316099
rect 249195 312084 249261 312085
rect 249195 312020 249196 312084
rect 249260 312020 249261 312084
rect 249195 312019 249261 312020
rect 249379 311812 249445 311813
rect 249379 311748 249380 311812
rect 249444 311748 249445 311812
rect 249379 311747 249445 311748
rect 249382 306373 249442 311747
rect 251403 307732 251469 307733
rect 251403 307668 251404 307732
rect 251468 307668 251469 307732
rect 251403 307667 251469 307668
rect 249379 306372 249445 306373
rect 249379 306308 249380 306372
rect 249444 306308 249445 306372
rect 249379 306307 249445 306308
rect 251406 298213 251466 307667
rect 251403 298212 251469 298213
rect 251403 298148 251404 298212
rect 251468 298148 251469 298212
rect 251403 298147 251469 298148
rect 249195 296852 249261 296853
rect 249195 296788 249196 296852
rect 249260 296788 249261 296852
rect 249195 296787 249261 296788
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 249198 275093 249258 296787
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 249195 275092 249261 275093
rect 249195 275028 249196 275092
rect 249260 275028 249261 275092
rect 249195 275027 249261 275028
rect 249379 267884 249445 267885
rect 249379 267820 249380 267884
rect 249444 267820 249445 267884
rect 249379 267819 249445 267820
rect 249382 265570 249442 267819
rect 249198 265510 249442 265570
rect 249198 257957 249258 265510
rect 249195 257956 249261 257957
rect 249195 257892 249196 257956
rect 249260 257892 249261 257956
rect 249195 257891 249261 257892
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 249011 248436 249077 248437
rect 249011 248372 249012 248436
rect 249076 248372 249077 248436
rect 249011 248371 249077 248372
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 249014 230621 249074 248371
rect 249011 230620 249077 230621
rect 249011 230556 249012 230620
rect 249076 230556 249077 230620
rect 249011 230555 249077 230556
rect 249379 230484 249445 230485
rect 249379 230420 249380 230484
rect 249444 230420 249445 230484
rect 249379 230419 249445 230420
rect 249382 219333 249442 230419
rect 249379 219332 249445 219333
rect 249379 219268 249380 219332
rect 249444 219268 249445 219332
rect 249379 219267 249445 219268
rect 249747 219196 249813 219197
rect 249747 219132 249748 219196
rect 249812 219132 249813 219196
rect 249747 219131 249813 219132
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 249750 209677 249810 219131
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 249747 209676 249813 209677
rect 249747 209612 249748 209676
rect 249812 209612 249813 209676
rect 249747 209611 249813 209612
rect 249563 200156 249629 200157
rect 249563 200092 249564 200156
rect 249628 200092 249629 200156
rect 249563 200091 249629 200092
rect 249566 193221 249626 200091
rect 249563 193220 249629 193221
rect 249563 193156 249564 193220
rect 249628 193156 249629 193220
rect 249563 193155 249629 193156
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 249011 182204 249077 182205
rect 249011 182140 249012 182204
rect 249076 182140 249077 182204
rect 249011 182139 249077 182140
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 249014 166970 249074 182139
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 249014 166910 249626 166970
rect 249566 157589 249626 166910
rect 249563 157588 249629 157589
rect 249563 157524 249564 157588
rect 249628 157524 249629 157588
rect 249563 157523 249629 157524
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 244043 110804 244109 110805
rect 244043 110740 244044 110804
rect 244108 110740 244109 110804
rect 244043 110739 244109 110740
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 241467 87548 241533 87549
rect 241467 87484 241468 87548
rect 241532 87484 241533 87548
rect 241467 87483 241533 87484
rect 241470 87141 241530 87483
rect 241467 87140 241533 87141
rect 241467 87076 241468 87140
rect 241532 87076 241533 87140
rect 241467 87075 241533 87076
rect 241102 77150 241346 77210
rect 241102 75989 241162 77150
rect 241099 75988 241165 75989
rect 241099 75924 241100 75988
rect 241164 75924 241165 75988
rect 241099 75923 241165 75924
rect 241467 75988 241533 75989
rect 241467 75924 241468 75988
rect 241532 75924 241533 75988
rect 241467 75923 241533 75924
rect 241470 75717 241530 75923
rect 241467 75716 241533 75717
rect 241467 75652 241468 75716
rect 241532 75652 241533 75716
rect 241467 75651 241533 75652
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 235763 29204 235829 29205
rect 235763 29140 235764 29204
rect 235828 29140 235829 29204
rect 235763 29139 235829 29140
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 231715 17372 231781 17373
rect 231715 17308 231716 17372
rect 231780 17308 231781 17372
rect 231715 17307 231781 17308
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 239811 17372 239877 17373
rect 239811 17308 239812 17372
rect 239876 17308 239877 17372
rect 239811 17307 239877 17308
rect 239814 16690 239874 17307
rect 239995 16692 240061 16693
rect 239995 16690 239996 16692
rect 239814 16630 239996 16690
rect 239995 16628 239996 16630
rect 240060 16628 240061 16692
rect 239995 16627 240061 16628
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 251219 87276 251285 87277
rect 251219 87212 251220 87276
rect 251284 87212 251285 87276
rect 251219 87211 251285 87212
rect 251222 87141 251282 87211
rect 251219 87140 251285 87141
rect 251219 87076 251220 87140
rect 251284 87076 251285 87140
rect 251219 87075 251285 87076
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 249747 64020 249813 64021
rect 249747 63956 249748 64020
rect 249812 63956 249813 64020
rect 249747 63955 249813 63956
rect 249750 63749 249810 63955
rect 249747 63748 249813 63749
rect 249747 63684 249748 63748
rect 249812 63684 249813 63748
rect 249747 63683 249813 63684
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 260787 87412 260853 87413
rect 260787 87348 260788 87412
rect 260852 87348 260853 87412
rect 260787 87347 260853 87348
rect 260790 87141 260850 87347
rect 260787 87140 260853 87141
rect 260787 87076 260788 87140
rect 260852 87076 260853 87140
rect 260787 87075 260853 87076
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 269067 76260 269133 76261
rect 269067 76196 269068 76260
rect 269132 76196 269133 76260
rect 269067 76195 269133 76196
rect 269070 75989 269130 76195
rect 269067 75988 269133 75989
rect 269067 75924 269068 75988
rect 269132 75924 269133 75988
rect 269067 75923 269133 75924
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 260971 16828 261037 16829
rect 260971 16764 260972 16828
rect 261036 16764 261037 16828
rect 260971 16763 261037 16764
rect 260787 16692 260853 16693
rect 260787 16628 260788 16692
rect 260852 16690 260853 16692
rect 260974 16690 261034 16763
rect 260852 16630 261034 16690
rect 260852 16628 260853 16630
rect 260787 16627 260853 16628
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 277347 157724 277413 157725
rect 277347 157660 277348 157724
rect 277412 157660 277413 157724
rect 277347 157659 277413 157660
rect 277350 157453 277410 157659
rect 277347 157452 277413 157453
rect 277347 157388 277348 157452
rect 277412 157388 277413 157452
rect 277347 157387 277413 157388
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 277347 87412 277413 87413
rect 277347 87348 277348 87412
rect 277412 87348 277413 87412
rect 277347 87347 277413 87348
rect 277350 87141 277410 87347
rect 277347 87140 277413 87141
rect 277347 87076 277348 87140
rect 277412 87076 277413 87140
rect 277347 87075 277413 87076
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 63654 278604 99098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 285627 157996 285693 157997
rect 285627 157932 285628 157996
rect 285692 157932 285693 157996
rect 285627 157931 285693 157932
rect 285630 157725 285690 157931
rect 285627 157724 285693 157725
rect 285627 157660 285628 157724
rect 285692 157660 285693 157724
rect 285627 157659 285693 157660
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 280107 63884 280173 63885
rect 280107 63820 280108 63884
rect 280172 63820 280173 63884
rect 280107 63819 280173 63820
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 280110 63613 280170 63819
rect 280107 63612 280173 63613
rect 280107 63548 280108 63612
rect 280172 63548 280173 63612
rect 280107 63547 280173 63548
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 280107 29340 280173 29341
rect 280107 29276 280108 29340
rect 280172 29276 280173 29340
rect 280107 29275 280173 29276
rect 280110 29069 280170 29275
rect 280107 29068 280173 29069
rect 280107 29004 280108 29068
rect 280172 29004 280173 29068
rect 280107 29003 280173 29004
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278819 16556 278885 16557
rect 278819 16492 278820 16556
rect 278884 16492 278885 16556
rect 278819 16491 278885 16492
rect 278822 16285 278882 16491
rect 278819 16284 278885 16285
rect 278819 16220 278820 16284
rect 278884 16220 278885 16284
rect 278819 16219 278885 16220
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288387 29476 288453 29477
rect 288387 29412 288388 29476
rect 288452 29412 288453 29476
rect 288387 29411 288453 29412
rect 288390 29205 288450 29411
rect 288387 29204 288453 29205
rect 288387 29140 288388 29204
rect 288452 29140 288453 29204
rect 288387 29139 288453 29140
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 307707 110940 307773 110941
rect 307707 110876 307708 110940
rect 307772 110876 307773 110940
rect 307707 110875 307773 110876
rect 307523 110668 307589 110669
rect 307523 110604 307524 110668
rect 307588 110604 307589 110668
rect 307523 110603 307589 110604
rect 307526 110530 307586 110603
rect 307710 110530 307770 110875
rect 307526 110470 307770 110530
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 327027 76260 327093 76261
rect 327027 76196 327028 76260
rect 327092 76196 327093 76260
rect 327027 76195 327093 76196
rect 327030 75989 327090 76195
rect 327027 75988 327093 75989
rect 327027 75924 327028 75988
rect 327092 75924 327093 75988
rect 327027 75923 327093 75924
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 327027 63884 327093 63885
rect 327027 63820 327028 63884
rect 327092 63820 327093 63884
rect 327027 63819 327093 63820
rect 327030 63613 327090 63819
rect 327027 63612 327093 63613
rect 327027 63548 327028 63612
rect 327092 63548 327093 63612
rect 327027 63547 327093 63548
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 327027 40356 327093 40357
rect 327027 40292 327028 40356
rect 327092 40292 327093 40356
rect 327027 40291 327093 40292
rect 327030 40085 327090 40291
rect 327027 40084 327093 40085
rect 327027 40020 327028 40084
rect 327092 40020 327093 40084
rect 327027 40019 327093 40020
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 325739 29340 325805 29341
rect 325739 29276 325740 29340
rect 325804 29276 325805 29340
rect 325739 29275 325805 29276
rect 325742 29069 325802 29275
rect 325739 29068 325805 29069
rect 325739 29004 325740 29068
rect 325804 29004 325805 29068
rect 325739 29003 325805 29004
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 341379 299436 341445 299437
rect 341379 299372 341380 299436
rect 341444 299372 341445 299436
rect 341379 299371 341445 299372
rect 341382 289917 341442 299371
rect 341379 289916 341445 289917
rect 341379 289852 341380 289916
rect 341444 289852 341445 289916
rect 341379 289851 341445 289852
rect 341379 280124 341445 280125
rect 341379 280060 341380 280124
rect 341444 280060 341445 280124
rect 341379 280059 341445 280060
rect 341382 270605 341442 280059
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 341379 270604 341445 270605
rect 341379 270540 341380 270604
rect 341444 270540 341445 270604
rect 341379 270539 341445 270540
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 341379 260812 341445 260813
rect 341379 260748 341380 260812
rect 341444 260748 341445 260812
rect 341379 260747 341445 260748
rect 341382 251293 341442 260747
rect 341379 251292 341445 251293
rect 341379 251228 341380 251292
rect 341444 251228 341445 251292
rect 341379 251227 341445 251228
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 337147 66196 337213 66197
rect 337147 66132 337148 66196
rect 337212 66132 337213 66196
rect 337147 66131 337213 66132
rect 337150 56677 337210 66131
rect 337147 56676 337213 56677
rect 337147 56612 337148 56676
rect 337212 56612 337213 56676
rect 337147 56611 337213 56612
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 366955 96932 367021 96933
rect 366955 96868 366956 96932
rect 367020 96868 367021 96932
rect 366955 96867 367021 96868
rect 366958 96661 367018 96867
rect 366955 96660 367021 96661
rect 366955 96596 366956 96660
rect 367020 96596 367021 96660
rect 366955 96595 367021 96596
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389403 118828 389469 118829
rect 389403 118764 389404 118828
rect 389468 118764 389469 118828
rect 389403 118763 389469 118764
rect 389406 108901 389466 118763
rect 389403 108900 389469 108901
rect 389403 108836 389404 108900
rect 389468 108836 389469 108900
rect 389403 108835 389469 108836
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396027 87548 396093 87549
rect 396027 87484 396028 87548
rect 396092 87484 396093 87548
rect 396027 87483 396093 87484
rect 396030 87141 396090 87483
rect 396027 87140 396093 87141
rect 396027 87076 396028 87140
rect 396092 87076 396093 87140
rect 396027 87075 396093 87076
rect 395843 76532 395909 76533
rect 395843 76468 395844 76532
rect 395908 76468 395909 76532
rect 395843 76467 395909 76468
rect 395846 76125 395906 76467
rect 395843 76124 395909 76125
rect 395843 76060 395844 76124
rect 395908 76060 395909 76124
rect 395843 76059 395909 76060
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396027 17100 396093 17101
rect 396027 17036 396028 17100
rect 396092 17036 396093 17100
rect 396027 17035 396093 17036
rect 396030 16693 396090 17035
rect 396027 16692 396093 16693
rect 396027 16628 396028 16692
rect 396092 16628 396093 16692
rect 396027 16627 396093 16628
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 405411 157860 405477 157861
rect 405411 157796 405412 157860
rect 405476 157796 405477 157860
rect 405411 157795 405477 157796
rect 405414 157450 405474 157795
rect 405595 157452 405661 157453
rect 405595 157450 405596 157452
rect 405414 157390 405596 157450
rect 405595 157388 405596 157390
rect 405660 157388 405661 157452
rect 405595 157387 405661 157388
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 405411 110940 405477 110941
rect 405411 110876 405412 110940
rect 405476 110876 405477 110940
rect 405411 110875 405477 110876
rect 405414 110530 405474 110875
rect 405595 110532 405661 110533
rect 405595 110530 405596 110532
rect 405414 110470 405596 110530
rect 405595 110468 405596 110470
rect 405660 110468 405661 110532
rect 405595 110467 405661 110468
rect 405595 87548 405661 87549
rect 405595 87484 405596 87548
rect 405660 87484 405661 87548
rect 405595 87483 405661 87484
rect 405598 87005 405658 87483
rect 405595 87004 405661 87005
rect 405595 86940 405596 87004
rect 405660 86940 405661 87004
rect 405595 86939 405661 86940
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 405411 64020 405477 64021
rect 405411 63956 405412 64020
rect 405476 63956 405477 64020
rect 405411 63955 405477 63956
rect 405414 63610 405474 63955
rect 405595 63612 405661 63613
rect 405595 63610 405596 63612
rect 405414 63550 405596 63610
rect 405595 63548 405596 63550
rect 405660 63548 405661 63612
rect 405595 63547 405661 63548
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 405595 29476 405661 29477
rect 405595 29412 405596 29476
rect 405660 29412 405661 29476
rect 405595 29411 405661 29412
rect 405598 29069 405658 29411
rect 405595 29068 405661 29069
rect 405595 29004 405596 29068
rect 405660 29004 405661 29068
rect 405595 29003 405661 29004
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 421235 196620 421301 196621
rect 421235 196556 421236 196620
rect 421300 196556 421301 196620
rect 421235 196555 421301 196556
rect 421238 183701 421298 196555
rect 421235 183700 421301 183701
rect 421235 183636 421236 183700
rect 421300 183636 421301 183700
rect 421235 183635 421301 183636
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 465947 583404 466013 583405
rect 465947 583340 465948 583404
rect 466012 583340 466013 583404
rect 465947 583339 466013 583340
rect 465763 583268 465829 583269
rect 465763 583204 465764 583268
rect 465828 583204 465829 583268
rect 465763 583203 465829 583204
rect 465579 579732 465645 579733
rect 465579 579668 465580 579732
rect 465644 579668 465645 579732
rect 465579 579667 465645 579668
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 465582 21997 465642 579667
rect 465766 486165 465826 583203
rect 465950 533085 466010 583339
rect 466499 579324 466565 579325
rect 466499 579260 466500 579324
rect 466564 579260 466565 579324
rect 466499 579259 466565 579260
rect 465947 533084 466013 533085
rect 465947 533020 465948 533084
rect 466012 533020 466013 533084
rect 465947 533019 466013 533020
rect 465763 486164 465829 486165
rect 465763 486100 465764 486164
rect 465828 486100 465829 486164
rect 465763 486099 465829 486100
rect 465579 21996 465645 21997
rect 465579 21932 465580 21996
rect 465644 21932 465645 21996
rect 465579 21931 465645 21932
rect 466502 11661 466562 579259
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 466499 11660 466565 11661
rect 466499 11596 466500 11660
rect 466564 11596 466565 11660
rect 466499 11595 466565 11596
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 473307 111076 473373 111077
rect 473307 111012 473308 111076
rect 473372 111012 473373 111076
rect 473307 111011 473373 111012
rect 473310 110805 473370 111011
rect 473307 110804 473373 110805
rect 473307 110740 473308 110804
rect 473372 110740 473373 110804
rect 473307 110739 473373 110740
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 473307 76532 473373 76533
rect 473307 76468 473308 76532
rect 473372 76468 473373 76532
rect 473307 76467 473373 76468
rect 473310 76261 473370 76467
rect 473307 76260 473373 76261
rect 473307 76196 473308 76260
rect 473372 76196 473373 76260
rect 473307 76195 473373 76196
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 473307 17236 473373 17237
rect 473307 17172 473308 17236
rect 473372 17172 473373 17236
rect 473307 17171 473373 17172
rect 473310 16965 473370 17171
rect 473307 16964 473373 16965
rect 473307 16900 473308 16964
rect 473372 16900 473373 16964
rect 473307 16899 473373 16900
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 481587 87412 481653 87413
rect 481587 87348 481588 87412
rect 481652 87348 481653 87412
rect 481587 87347 481653 87348
rect 481590 87141 481650 87347
rect 481587 87140 481653 87141
rect 481587 87076 481588 87140
rect 481652 87076 481653 87140
rect 481587 87075 481653 87076
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 481587 29476 481653 29477
rect 481587 29412 481588 29476
rect 481652 29412 481653 29476
rect 481587 29411 481653 29412
rect 481590 29205 481650 29411
rect 481587 29204 481653 29205
rect 481587 29140 481588 29204
rect 481652 29140 481653 29204
rect 481587 29139 481653 29140
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 492627 110804 492693 110805
rect 492627 110740 492628 110804
rect 492692 110740 492693 110804
rect 492627 110739 492693 110740
rect 492630 110533 492690 110739
rect 492627 110532 492693 110533
rect 492627 110468 492628 110532
rect 492692 110468 492693 110532
rect 492627 110467 492693 110468
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 492627 76260 492693 76261
rect 492627 76196 492628 76260
rect 492692 76196 492693 76260
rect 492627 76195 492693 76196
rect 492630 75989 492690 76195
rect 492627 75988 492693 75989
rect 492627 75924 492628 75988
rect 492692 75924 492693 75988
rect 492627 75923 492693 75924
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 492627 16964 492693 16965
rect 492627 16900 492628 16964
rect 492692 16900 492693 16964
rect 492627 16899 492693 16900
rect 492630 16693 492690 16899
rect 492627 16692 492693 16693
rect 492627 16628 492628 16692
rect 492692 16628 492693 16692
rect 492627 16627 492693 16628
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 243590 432702 243826 432938
rect 243590 413662 243826 413898
rect 243038 412982 243274 413218
rect 243038 406862 243274 407098
rect 243590 406182 243826 406418
rect 243222 395982 243458 396218
rect 243590 395982 243826 396218
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 249294 431342 249530 431578
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 252986 181898 253222 182134
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect 243548 432938 248468 432980
rect 243548 432702 243590 432938
rect 243826 432702 248468 432938
rect 243548 432660 248468 432702
rect 248148 431620 248468 432660
rect 248148 431578 249572 431620
rect 248148 431342 249294 431578
rect 249530 431342 249572 431578
rect 248148 431300 249572 431342
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect 243548 413898 243868 413940
rect 243548 413662 243590 413898
rect 243826 413662 243868 413898
rect 243548 413260 243868 413662
rect 242996 413218 243868 413260
rect 242996 412982 243038 413218
rect 243274 412982 243868 413218
rect 242996 412940 243868 412982
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect 242996 407098 243316 407140
rect 242996 406862 243038 407098
rect 243274 406862 243316 407098
rect 242996 406460 243316 406862
rect 242996 406418 243868 406460
rect 242996 406182 243590 406418
rect 243826 406182 243868 406418
rect 242996 406140 243868 406182
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect 243180 396218 243868 396260
rect 243180 395982 243222 396218
rect 243458 395982 243590 396218
rect 243826 395982 243868 396218
rect 243180 395940 243868 395982
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1607998175
transform 1 0 230000 0 1 340000
box 0 0 239540 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
