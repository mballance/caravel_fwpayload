magic
tech sky130A
magscale 1 2
timestamp 1607632543
<< obsli1 >>
rect 814 2159 298526 297585
<< obsm1 >>
rect 0 892 299432 297616
<< metal2 >>
rect 1016 299200 1072 300000
rect 3592 299200 3648 300000
rect 6260 299200 6316 300000
rect 8836 299200 8892 300000
rect 11504 299200 11560 300000
rect 14172 299200 14228 300000
rect 16748 299200 16804 300000
rect 19416 299200 19472 300000
rect 21992 299200 22048 300000
rect 24660 299200 24716 300000
rect 27328 299200 27384 300000
rect 29904 299200 29960 300000
rect 32572 299200 32628 300000
rect 35148 299200 35204 300000
rect 37816 299200 37872 300000
rect 40484 299200 40540 300000
rect 43060 299200 43116 300000
rect 45728 299200 45784 300000
rect 48304 299200 48360 300000
rect 50972 299200 51028 300000
rect 53640 299200 53696 300000
rect 56216 299200 56272 300000
rect 58884 299200 58940 300000
rect 61460 299200 61516 300000
rect 64128 299200 64184 300000
rect 66796 299200 66852 300000
rect 69372 299200 69428 300000
rect 72040 299200 72096 300000
rect 74616 299200 74672 300000
rect 77284 299200 77340 300000
rect 79952 299200 80008 300000
rect 82528 299200 82584 300000
rect 85196 299200 85252 300000
rect 87772 299200 87828 300000
rect 90440 299200 90496 300000
rect 93108 299200 93164 300000
rect 95684 299200 95740 300000
rect 98352 299200 98408 300000
rect 101020 299200 101076 300000
rect 103596 299200 103652 300000
rect 106264 299200 106320 300000
rect 108840 299200 108896 300000
rect 111508 299200 111564 300000
rect 114176 299200 114232 300000
rect 116752 299200 116808 300000
rect 119420 299200 119476 300000
rect 121996 299200 122052 300000
rect 124664 299200 124720 300000
rect 127332 299200 127388 300000
rect 129908 299200 129964 300000
rect 132576 299200 132632 300000
rect 135152 299200 135208 300000
rect 137820 299200 137876 300000
rect 140488 299200 140544 300000
rect 143064 299200 143120 300000
rect 145732 299200 145788 300000
rect 148308 299200 148364 300000
rect 150976 299200 151032 300000
rect 153644 299200 153700 300000
rect 156220 299200 156276 300000
rect 158888 299200 158944 300000
rect 161464 299200 161520 300000
rect 164132 299200 164188 300000
rect 166800 299200 166856 300000
rect 169376 299200 169432 300000
rect 172044 299200 172100 300000
rect 174620 299200 174676 300000
rect 177288 299200 177344 300000
rect 179956 299200 180012 300000
rect 182532 299200 182588 300000
rect 185200 299200 185256 300000
rect 187776 299200 187832 300000
rect 190444 299200 190500 300000
rect 193112 299200 193168 300000
rect 195688 299200 195744 300000
rect 198356 299200 198412 300000
rect 201024 299200 201080 300000
rect 203600 299200 203656 300000
rect 206268 299200 206324 300000
rect 208844 299200 208900 300000
rect 211512 299200 211568 300000
rect 214180 299200 214236 300000
rect 216756 299200 216812 300000
rect 219424 299200 219480 300000
rect 222000 299200 222056 300000
rect 224668 299200 224724 300000
rect 227336 299200 227392 300000
rect 229912 299200 229968 300000
rect 232580 299200 232636 300000
rect 235156 299200 235212 300000
rect 237824 299200 237880 300000
rect 240492 299200 240548 300000
rect 243068 299200 243124 300000
rect 245736 299200 245792 300000
rect 248312 299200 248368 300000
rect 250980 299200 251036 300000
rect 253648 299200 253704 300000
rect 256224 299200 256280 300000
rect 258892 299200 258948 300000
rect 261468 299200 261524 300000
rect 264136 299200 264192 300000
rect 266804 299200 266860 300000
rect 269380 299200 269436 300000
rect 272048 299200 272104 300000
rect 274624 299200 274680 300000
rect 277292 299200 277348 300000
rect 279960 299200 280016 300000
rect 282536 299200 282592 300000
rect 285204 299200 285260 300000
rect 287780 299200 287836 300000
rect 290448 299200 290504 300000
rect 293116 299200 293172 300000
rect 295692 299200 295748 300000
rect 298360 299200 298416 300000
rect 4 0 60 800
rect 556 0 612 800
rect 1200 0 1256 800
rect 1752 0 1808 800
rect 2396 0 2452 800
rect 3040 0 3096 800
rect 3592 0 3648 800
rect 4236 0 4292 800
rect 4880 0 4936 800
rect 5432 0 5488 800
rect 6076 0 6132 800
rect 6720 0 6776 800
rect 7272 0 7328 800
rect 7916 0 7972 800
rect 8560 0 8616 800
rect 9112 0 9168 800
rect 9756 0 9812 800
rect 10400 0 10456 800
rect 10952 0 11008 800
rect 11596 0 11652 800
rect 12240 0 12296 800
rect 12792 0 12848 800
rect 13436 0 13492 800
rect 14080 0 14136 800
rect 14632 0 14688 800
rect 15276 0 15332 800
rect 15920 0 15976 800
rect 16472 0 16528 800
rect 17116 0 17172 800
rect 17668 0 17724 800
rect 18312 0 18368 800
rect 18956 0 19012 800
rect 19508 0 19564 800
rect 20152 0 20208 800
rect 20796 0 20852 800
rect 21348 0 21404 800
rect 21992 0 22048 800
rect 22636 0 22692 800
rect 23188 0 23244 800
rect 23832 0 23888 800
rect 24476 0 24532 800
rect 25028 0 25084 800
rect 25672 0 25728 800
rect 26316 0 26372 800
rect 26868 0 26924 800
rect 27512 0 27568 800
rect 28156 0 28212 800
rect 28708 0 28764 800
rect 29352 0 29408 800
rect 29996 0 30052 800
rect 30548 0 30604 800
rect 31192 0 31248 800
rect 31836 0 31892 800
rect 32388 0 32444 800
rect 33032 0 33088 800
rect 33676 0 33732 800
rect 34228 0 34284 800
rect 34872 0 34928 800
rect 35424 0 35480 800
rect 36068 0 36124 800
rect 36712 0 36768 800
rect 37264 0 37320 800
rect 37908 0 37964 800
rect 38552 0 38608 800
rect 39104 0 39160 800
rect 39748 0 39804 800
rect 40392 0 40448 800
rect 40944 0 41000 800
rect 41588 0 41644 800
rect 42232 0 42288 800
rect 42784 0 42840 800
rect 43428 0 43484 800
rect 44072 0 44128 800
rect 44624 0 44680 800
rect 45268 0 45324 800
rect 45912 0 45968 800
rect 46464 0 46520 800
rect 47108 0 47164 800
rect 47752 0 47808 800
rect 48304 0 48360 800
rect 48948 0 49004 800
rect 49592 0 49648 800
rect 50144 0 50200 800
rect 50788 0 50844 800
rect 51432 0 51488 800
rect 51984 0 52040 800
rect 52628 0 52684 800
rect 53180 0 53236 800
rect 53824 0 53880 800
rect 54468 0 54524 800
rect 55020 0 55076 800
rect 55664 0 55720 800
rect 56308 0 56364 800
rect 56860 0 56916 800
rect 57504 0 57560 800
rect 58148 0 58204 800
rect 58700 0 58756 800
rect 59344 0 59400 800
rect 59988 0 60044 800
rect 60540 0 60596 800
rect 61184 0 61240 800
rect 61828 0 61884 800
rect 62380 0 62436 800
rect 63024 0 63080 800
rect 63668 0 63724 800
rect 64220 0 64276 800
rect 64864 0 64920 800
rect 65508 0 65564 800
rect 66060 0 66116 800
rect 66704 0 66760 800
rect 67348 0 67404 800
rect 67900 0 67956 800
rect 68544 0 68600 800
rect 69188 0 69244 800
rect 69740 0 69796 800
rect 70384 0 70440 800
rect 70936 0 70992 800
rect 71580 0 71636 800
rect 72224 0 72280 800
rect 72776 0 72832 800
rect 73420 0 73476 800
rect 74064 0 74120 800
rect 74616 0 74672 800
rect 75260 0 75316 800
rect 75904 0 75960 800
rect 76456 0 76512 800
rect 77100 0 77156 800
rect 77744 0 77800 800
rect 78296 0 78352 800
rect 78940 0 78996 800
rect 79584 0 79640 800
rect 80136 0 80192 800
rect 80780 0 80836 800
rect 81424 0 81480 800
rect 81976 0 82032 800
rect 82620 0 82676 800
rect 83264 0 83320 800
rect 83816 0 83872 800
rect 84460 0 84516 800
rect 85104 0 85160 800
rect 85656 0 85712 800
rect 86300 0 86356 800
rect 86944 0 87000 800
rect 87496 0 87552 800
rect 88140 0 88196 800
rect 88692 0 88748 800
rect 89336 0 89392 800
rect 89980 0 90036 800
rect 90532 0 90588 800
rect 91176 0 91232 800
rect 91820 0 91876 800
rect 92372 0 92428 800
rect 93016 0 93072 800
rect 93660 0 93716 800
rect 94212 0 94268 800
rect 94856 0 94912 800
rect 95500 0 95556 800
rect 96052 0 96108 800
rect 96696 0 96752 800
rect 97340 0 97396 800
rect 97892 0 97948 800
rect 98536 0 98592 800
rect 99180 0 99236 800
rect 99732 0 99788 800
rect 100376 0 100432 800
rect 101020 0 101076 800
rect 101572 0 101628 800
rect 102216 0 102272 800
rect 102860 0 102916 800
rect 103412 0 103468 800
rect 104056 0 104112 800
rect 104700 0 104756 800
rect 105252 0 105308 800
rect 105896 0 105952 800
rect 106448 0 106504 800
rect 107092 0 107148 800
rect 107736 0 107792 800
rect 108288 0 108344 800
rect 108932 0 108988 800
rect 109576 0 109632 800
rect 110128 0 110184 800
rect 110772 0 110828 800
rect 111416 0 111472 800
rect 111968 0 112024 800
rect 112612 0 112668 800
rect 113256 0 113312 800
rect 113808 0 113864 800
rect 114452 0 114508 800
rect 115096 0 115152 800
rect 115648 0 115704 800
rect 116292 0 116348 800
rect 116936 0 116992 800
rect 117488 0 117544 800
rect 118132 0 118188 800
rect 118776 0 118832 800
rect 119328 0 119384 800
rect 119972 0 120028 800
rect 120616 0 120672 800
rect 121168 0 121224 800
rect 121812 0 121868 800
rect 122456 0 122512 800
rect 123008 0 123064 800
rect 123652 0 123708 800
rect 124204 0 124260 800
rect 124848 0 124904 800
rect 125492 0 125548 800
rect 126044 0 126100 800
rect 126688 0 126744 800
rect 127332 0 127388 800
rect 127884 0 127940 800
rect 128528 0 128584 800
rect 129172 0 129228 800
rect 129724 0 129780 800
rect 130368 0 130424 800
rect 131012 0 131068 800
rect 131564 0 131620 800
rect 132208 0 132264 800
rect 132852 0 132908 800
rect 133404 0 133460 800
rect 134048 0 134104 800
rect 134692 0 134748 800
rect 135244 0 135300 800
rect 135888 0 135944 800
rect 136532 0 136588 800
rect 137084 0 137140 800
rect 137728 0 137784 800
rect 138372 0 138428 800
rect 138924 0 138980 800
rect 139568 0 139624 800
rect 140212 0 140268 800
rect 140764 0 140820 800
rect 141408 0 141464 800
rect 141960 0 142016 800
rect 142604 0 142660 800
rect 143248 0 143304 800
rect 143800 0 143856 800
rect 144444 0 144500 800
rect 145088 0 145144 800
rect 145640 0 145696 800
rect 146284 0 146340 800
rect 146928 0 146984 800
rect 147480 0 147536 800
rect 148124 0 148180 800
rect 148768 0 148824 800
rect 149320 0 149376 800
rect 149964 0 150020 800
rect 150608 0 150664 800
rect 151160 0 151216 800
rect 151804 0 151860 800
rect 152448 0 152504 800
rect 153000 0 153056 800
rect 153644 0 153700 800
rect 154288 0 154344 800
rect 154840 0 154896 800
rect 155484 0 155540 800
rect 156128 0 156184 800
rect 156680 0 156736 800
rect 157324 0 157380 800
rect 157968 0 158024 800
rect 158520 0 158576 800
rect 159164 0 159220 800
rect 159716 0 159772 800
rect 160360 0 160416 800
rect 161004 0 161060 800
rect 161556 0 161612 800
rect 162200 0 162256 800
rect 162844 0 162900 800
rect 163396 0 163452 800
rect 164040 0 164096 800
rect 164684 0 164740 800
rect 165236 0 165292 800
rect 165880 0 165936 800
rect 166524 0 166580 800
rect 167076 0 167132 800
rect 167720 0 167776 800
rect 168364 0 168420 800
rect 168916 0 168972 800
rect 169560 0 169616 800
rect 170204 0 170260 800
rect 170756 0 170812 800
rect 171400 0 171456 800
rect 172044 0 172100 800
rect 172596 0 172652 800
rect 173240 0 173296 800
rect 173884 0 173940 800
rect 174436 0 174492 800
rect 175080 0 175136 800
rect 175724 0 175780 800
rect 176276 0 176332 800
rect 176920 0 176976 800
rect 177472 0 177528 800
rect 178116 0 178172 800
rect 178760 0 178816 800
rect 179312 0 179368 800
rect 179956 0 180012 800
rect 180600 0 180656 800
rect 181152 0 181208 800
rect 181796 0 181852 800
rect 182440 0 182496 800
rect 182992 0 183048 800
rect 183636 0 183692 800
rect 184280 0 184336 800
rect 184832 0 184888 800
rect 185476 0 185532 800
rect 186120 0 186176 800
rect 186672 0 186728 800
rect 187316 0 187372 800
rect 187960 0 188016 800
rect 188512 0 188568 800
rect 189156 0 189212 800
rect 189800 0 189856 800
rect 190352 0 190408 800
rect 190996 0 191052 800
rect 191640 0 191696 800
rect 192192 0 192248 800
rect 192836 0 192892 800
rect 193480 0 193536 800
rect 194032 0 194088 800
rect 194676 0 194732 800
rect 195228 0 195284 800
rect 195872 0 195928 800
rect 196516 0 196572 800
rect 197068 0 197124 800
rect 197712 0 197768 800
rect 198356 0 198412 800
rect 198908 0 198964 800
rect 199552 0 199608 800
rect 200196 0 200252 800
rect 200748 0 200804 800
rect 201392 0 201448 800
rect 202036 0 202092 800
rect 202588 0 202644 800
rect 203232 0 203288 800
rect 203876 0 203932 800
rect 204428 0 204484 800
rect 205072 0 205128 800
rect 205716 0 205772 800
rect 206268 0 206324 800
rect 206912 0 206968 800
rect 207556 0 207612 800
rect 208108 0 208164 800
rect 208752 0 208808 800
rect 209396 0 209452 800
rect 209948 0 210004 800
rect 210592 0 210648 800
rect 211236 0 211292 800
rect 211788 0 211844 800
rect 212432 0 212488 800
rect 212984 0 213040 800
rect 213628 0 213684 800
rect 214272 0 214328 800
rect 214824 0 214880 800
rect 215468 0 215524 800
rect 216112 0 216168 800
rect 216664 0 216720 800
rect 217308 0 217364 800
rect 217952 0 218008 800
rect 218504 0 218560 800
rect 219148 0 219204 800
rect 219792 0 219848 800
rect 220344 0 220400 800
rect 220988 0 221044 800
rect 221632 0 221688 800
rect 222184 0 222240 800
rect 222828 0 222884 800
rect 223472 0 223528 800
rect 224024 0 224080 800
rect 224668 0 224724 800
rect 225312 0 225368 800
rect 225864 0 225920 800
rect 226508 0 226564 800
rect 227152 0 227208 800
rect 227704 0 227760 800
rect 228348 0 228404 800
rect 228992 0 229048 800
rect 229544 0 229600 800
rect 230188 0 230244 800
rect 230740 0 230796 800
rect 231384 0 231440 800
rect 232028 0 232084 800
rect 232580 0 232636 800
rect 233224 0 233280 800
rect 233868 0 233924 800
rect 234420 0 234476 800
rect 235064 0 235120 800
rect 235708 0 235764 800
rect 236260 0 236316 800
rect 236904 0 236960 800
rect 237548 0 237604 800
rect 238100 0 238156 800
rect 238744 0 238800 800
rect 239388 0 239444 800
rect 239940 0 239996 800
rect 240584 0 240640 800
rect 241228 0 241284 800
rect 241780 0 241836 800
rect 242424 0 242480 800
rect 243068 0 243124 800
rect 243620 0 243676 800
rect 244264 0 244320 800
rect 244908 0 244964 800
rect 245460 0 245516 800
rect 246104 0 246160 800
rect 246748 0 246804 800
rect 247300 0 247356 800
rect 247944 0 248000 800
rect 248496 0 248552 800
rect 249140 0 249196 800
rect 249784 0 249840 800
rect 250336 0 250392 800
rect 250980 0 251036 800
rect 251624 0 251680 800
rect 252176 0 252232 800
rect 252820 0 252876 800
rect 253464 0 253520 800
rect 254016 0 254072 800
rect 254660 0 254716 800
rect 255304 0 255360 800
rect 255856 0 255912 800
rect 256500 0 256556 800
rect 257144 0 257200 800
rect 257696 0 257752 800
rect 258340 0 258396 800
rect 258984 0 259040 800
rect 259536 0 259592 800
rect 260180 0 260236 800
rect 260824 0 260880 800
rect 261376 0 261432 800
rect 262020 0 262076 800
rect 262664 0 262720 800
rect 263216 0 263272 800
rect 263860 0 263916 800
rect 264504 0 264560 800
rect 265056 0 265112 800
rect 265700 0 265756 800
rect 266252 0 266308 800
rect 266896 0 266952 800
rect 267540 0 267596 800
rect 268092 0 268148 800
rect 268736 0 268792 800
rect 269380 0 269436 800
rect 269932 0 269988 800
rect 270576 0 270632 800
rect 271220 0 271276 800
rect 271772 0 271828 800
rect 272416 0 272472 800
rect 273060 0 273116 800
rect 273612 0 273668 800
rect 274256 0 274312 800
rect 274900 0 274956 800
rect 275452 0 275508 800
rect 276096 0 276152 800
rect 276740 0 276796 800
rect 277292 0 277348 800
rect 277936 0 277992 800
rect 278580 0 278636 800
rect 279132 0 279188 800
rect 279776 0 279832 800
rect 280420 0 280476 800
rect 280972 0 281028 800
rect 281616 0 281672 800
rect 282260 0 282316 800
rect 282812 0 282868 800
rect 283456 0 283512 800
rect 284008 0 284064 800
rect 284652 0 284708 800
rect 285296 0 285352 800
rect 285848 0 285904 800
rect 286492 0 286548 800
rect 287136 0 287192 800
rect 287688 0 287744 800
rect 288332 0 288388 800
rect 288976 0 289032 800
rect 289528 0 289584 800
rect 290172 0 290228 800
rect 290816 0 290872 800
rect 291368 0 291424 800
rect 292012 0 292068 800
rect 292656 0 292712 800
rect 293208 0 293264 800
rect 293852 0 293908 800
rect 294496 0 294552 800
rect 295048 0 295104 800
rect 295692 0 295748 800
rect 296336 0 296392 800
rect 296888 0 296944 800
rect 297532 0 297588 800
rect 298176 0 298232 800
rect 298728 0 298784 800
rect 299372 0 299428 800
<< obsm2 >>
rect 6 299144 960 299200
rect 1128 299144 3536 299200
rect 3704 299144 6204 299200
rect 6372 299144 8780 299200
rect 8948 299144 11448 299200
rect 11616 299144 14116 299200
rect 14284 299144 16692 299200
rect 16860 299144 19360 299200
rect 19528 299144 21936 299200
rect 22104 299144 24604 299200
rect 24772 299144 27272 299200
rect 27440 299144 29848 299200
rect 30016 299144 32516 299200
rect 32684 299144 35092 299200
rect 35260 299144 37760 299200
rect 37928 299144 40428 299200
rect 40596 299144 43004 299200
rect 43172 299144 45672 299200
rect 45840 299144 48248 299200
rect 48416 299144 50916 299200
rect 51084 299144 53584 299200
rect 53752 299144 56160 299200
rect 56328 299144 58828 299200
rect 58996 299144 61404 299200
rect 61572 299144 64072 299200
rect 64240 299144 66740 299200
rect 66908 299144 69316 299200
rect 69484 299144 71984 299200
rect 72152 299144 74560 299200
rect 74728 299144 77228 299200
rect 77396 299144 79896 299200
rect 80064 299144 82472 299200
rect 82640 299144 85140 299200
rect 85308 299144 87716 299200
rect 87884 299144 90384 299200
rect 90552 299144 93052 299200
rect 93220 299144 95628 299200
rect 95796 299144 98296 299200
rect 98464 299144 100964 299200
rect 101132 299144 103540 299200
rect 103708 299144 106208 299200
rect 106376 299144 108784 299200
rect 108952 299144 111452 299200
rect 111620 299144 114120 299200
rect 114288 299144 116696 299200
rect 116864 299144 119364 299200
rect 119532 299144 121940 299200
rect 122108 299144 124608 299200
rect 124776 299144 127276 299200
rect 127444 299144 129852 299200
rect 130020 299144 132520 299200
rect 132688 299144 135096 299200
rect 135264 299144 137764 299200
rect 137932 299144 140432 299200
rect 140600 299144 143008 299200
rect 143176 299144 145676 299200
rect 145844 299144 148252 299200
rect 148420 299144 150920 299200
rect 151088 299144 153588 299200
rect 153756 299144 156164 299200
rect 156332 299144 158832 299200
rect 159000 299144 161408 299200
rect 161576 299144 164076 299200
rect 164244 299144 166744 299200
rect 166912 299144 169320 299200
rect 169488 299144 171988 299200
rect 172156 299144 174564 299200
rect 174732 299144 177232 299200
rect 177400 299144 179900 299200
rect 180068 299144 182476 299200
rect 182644 299144 185144 299200
rect 185312 299144 187720 299200
rect 187888 299144 190388 299200
rect 190556 299144 193056 299200
rect 193224 299144 195632 299200
rect 195800 299144 198300 299200
rect 198468 299144 200968 299200
rect 201136 299144 203544 299200
rect 203712 299144 206212 299200
rect 206380 299144 208788 299200
rect 208956 299144 211456 299200
rect 211624 299144 214124 299200
rect 214292 299144 216700 299200
rect 216868 299144 219368 299200
rect 219536 299144 221944 299200
rect 222112 299144 224612 299200
rect 224780 299144 227280 299200
rect 227448 299144 229856 299200
rect 230024 299144 232524 299200
rect 232692 299144 235100 299200
rect 235268 299144 237768 299200
rect 237936 299144 240436 299200
rect 240604 299144 243012 299200
rect 243180 299144 245680 299200
rect 245848 299144 248256 299200
rect 248424 299144 250924 299200
rect 251092 299144 253592 299200
rect 253760 299144 256168 299200
rect 256336 299144 258836 299200
rect 259004 299144 261412 299200
rect 261580 299144 264080 299200
rect 264248 299144 266748 299200
rect 266916 299144 269324 299200
rect 269492 299144 271992 299200
rect 272160 299144 274568 299200
rect 274736 299144 277236 299200
rect 277404 299144 279904 299200
rect 280072 299144 282480 299200
rect 282648 299144 285148 299200
rect 285316 299144 287724 299200
rect 287892 299144 290392 299200
rect 290560 299144 293060 299200
rect 293228 299144 295636 299200
rect 295804 299144 298304 299200
rect 298472 299144 299426 299200
rect 6 856 299426 299144
rect 116 800 500 856
rect 668 800 1144 856
rect 1312 800 1696 856
rect 1864 800 2340 856
rect 2508 800 2984 856
rect 3152 800 3536 856
rect 3704 800 4180 856
rect 4348 800 4824 856
rect 4992 800 5376 856
rect 5544 800 6020 856
rect 6188 800 6664 856
rect 6832 800 7216 856
rect 7384 800 7860 856
rect 8028 800 8504 856
rect 8672 800 9056 856
rect 9224 800 9700 856
rect 9868 800 10344 856
rect 10512 800 10896 856
rect 11064 800 11540 856
rect 11708 800 12184 856
rect 12352 800 12736 856
rect 12904 800 13380 856
rect 13548 800 14024 856
rect 14192 800 14576 856
rect 14744 800 15220 856
rect 15388 800 15864 856
rect 16032 800 16416 856
rect 16584 800 17060 856
rect 17228 800 17612 856
rect 17780 800 18256 856
rect 18424 800 18900 856
rect 19068 800 19452 856
rect 19620 800 20096 856
rect 20264 800 20740 856
rect 20908 800 21292 856
rect 21460 800 21936 856
rect 22104 800 22580 856
rect 22748 800 23132 856
rect 23300 800 23776 856
rect 23944 800 24420 856
rect 24588 800 24972 856
rect 25140 800 25616 856
rect 25784 800 26260 856
rect 26428 800 26812 856
rect 26980 800 27456 856
rect 27624 800 28100 856
rect 28268 800 28652 856
rect 28820 800 29296 856
rect 29464 800 29940 856
rect 30108 800 30492 856
rect 30660 800 31136 856
rect 31304 800 31780 856
rect 31948 800 32332 856
rect 32500 800 32976 856
rect 33144 800 33620 856
rect 33788 800 34172 856
rect 34340 800 34816 856
rect 34984 800 35368 856
rect 35536 800 36012 856
rect 36180 800 36656 856
rect 36824 800 37208 856
rect 37376 800 37852 856
rect 38020 800 38496 856
rect 38664 800 39048 856
rect 39216 800 39692 856
rect 39860 800 40336 856
rect 40504 800 40888 856
rect 41056 800 41532 856
rect 41700 800 42176 856
rect 42344 800 42728 856
rect 42896 800 43372 856
rect 43540 800 44016 856
rect 44184 800 44568 856
rect 44736 800 45212 856
rect 45380 800 45856 856
rect 46024 800 46408 856
rect 46576 800 47052 856
rect 47220 800 47696 856
rect 47864 800 48248 856
rect 48416 800 48892 856
rect 49060 800 49536 856
rect 49704 800 50088 856
rect 50256 800 50732 856
rect 50900 800 51376 856
rect 51544 800 51928 856
rect 52096 800 52572 856
rect 52740 800 53124 856
rect 53292 800 53768 856
rect 53936 800 54412 856
rect 54580 800 54964 856
rect 55132 800 55608 856
rect 55776 800 56252 856
rect 56420 800 56804 856
rect 56972 800 57448 856
rect 57616 800 58092 856
rect 58260 800 58644 856
rect 58812 800 59288 856
rect 59456 800 59932 856
rect 60100 800 60484 856
rect 60652 800 61128 856
rect 61296 800 61772 856
rect 61940 800 62324 856
rect 62492 800 62968 856
rect 63136 800 63612 856
rect 63780 800 64164 856
rect 64332 800 64808 856
rect 64976 800 65452 856
rect 65620 800 66004 856
rect 66172 800 66648 856
rect 66816 800 67292 856
rect 67460 800 67844 856
rect 68012 800 68488 856
rect 68656 800 69132 856
rect 69300 800 69684 856
rect 69852 800 70328 856
rect 70496 800 70880 856
rect 71048 800 71524 856
rect 71692 800 72168 856
rect 72336 800 72720 856
rect 72888 800 73364 856
rect 73532 800 74008 856
rect 74176 800 74560 856
rect 74728 800 75204 856
rect 75372 800 75848 856
rect 76016 800 76400 856
rect 76568 800 77044 856
rect 77212 800 77688 856
rect 77856 800 78240 856
rect 78408 800 78884 856
rect 79052 800 79528 856
rect 79696 800 80080 856
rect 80248 800 80724 856
rect 80892 800 81368 856
rect 81536 800 81920 856
rect 82088 800 82564 856
rect 82732 800 83208 856
rect 83376 800 83760 856
rect 83928 800 84404 856
rect 84572 800 85048 856
rect 85216 800 85600 856
rect 85768 800 86244 856
rect 86412 800 86888 856
rect 87056 800 87440 856
rect 87608 800 88084 856
rect 88252 800 88636 856
rect 88804 800 89280 856
rect 89448 800 89924 856
rect 90092 800 90476 856
rect 90644 800 91120 856
rect 91288 800 91764 856
rect 91932 800 92316 856
rect 92484 800 92960 856
rect 93128 800 93604 856
rect 93772 800 94156 856
rect 94324 800 94800 856
rect 94968 800 95444 856
rect 95612 800 95996 856
rect 96164 800 96640 856
rect 96808 800 97284 856
rect 97452 800 97836 856
rect 98004 800 98480 856
rect 98648 800 99124 856
rect 99292 800 99676 856
rect 99844 800 100320 856
rect 100488 800 100964 856
rect 101132 800 101516 856
rect 101684 800 102160 856
rect 102328 800 102804 856
rect 102972 800 103356 856
rect 103524 800 104000 856
rect 104168 800 104644 856
rect 104812 800 105196 856
rect 105364 800 105840 856
rect 106008 800 106392 856
rect 106560 800 107036 856
rect 107204 800 107680 856
rect 107848 800 108232 856
rect 108400 800 108876 856
rect 109044 800 109520 856
rect 109688 800 110072 856
rect 110240 800 110716 856
rect 110884 800 111360 856
rect 111528 800 111912 856
rect 112080 800 112556 856
rect 112724 800 113200 856
rect 113368 800 113752 856
rect 113920 800 114396 856
rect 114564 800 115040 856
rect 115208 800 115592 856
rect 115760 800 116236 856
rect 116404 800 116880 856
rect 117048 800 117432 856
rect 117600 800 118076 856
rect 118244 800 118720 856
rect 118888 800 119272 856
rect 119440 800 119916 856
rect 120084 800 120560 856
rect 120728 800 121112 856
rect 121280 800 121756 856
rect 121924 800 122400 856
rect 122568 800 122952 856
rect 123120 800 123596 856
rect 123764 800 124148 856
rect 124316 800 124792 856
rect 124960 800 125436 856
rect 125604 800 125988 856
rect 126156 800 126632 856
rect 126800 800 127276 856
rect 127444 800 127828 856
rect 127996 800 128472 856
rect 128640 800 129116 856
rect 129284 800 129668 856
rect 129836 800 130312 856
rect 130480 800 130956 856
rect 131124 800 131508 856
rect 131676 800 132152 856
rect 132320 800 132796 856
rect 132964 800 133348 856
rect 133516 800 133992 856
rect 134160 800 134636 856
rect 134804 800 135188 856
rect 135356 800 135832 856
rect 136000 800 136476 856
rect 136644 800 137028 856
rect 137196 800 137672 856
rect 137840 800 138316 856
rect 138484 800 138868 856
rect 139036 800 139512 856
rect 139680 800 140156 856
rect 140324 800 140708 856
rect 140876 800 141352 856
rect 141520 800 141904 856
rect 142072 800 142548 856
rect 142716 800 143192 856
rect 143360 800 143744 856
rect 143912 800 144388 856
rect 144556 800 145032 856
rect 145200 800 145584 856
rect 145752 800 146228 856
rect 146396 800 146872 856
rect 147040 800 147424 856
rect 147592 800 148068 856
rect 148236 800 148712 856
rect 148880 800 149264 856
rect 149432 800 149908 856
rect 150076 800 150552 856
rect 150720 800 151104 856
rect 151272 800 151748 856
rect 151916 800 152392 856
rect 152560 800 152944 856
rect 153112 800 153588 856
rect 153756 800 154232 856
rect 154400 800 154784 856
rect 154952 800 155428 856
rect 155596 800 156072 856
rect 156240 800 156624 856
rect 156792 800 157268 856
rect 157436 800 157912 856
rect 158080 800 158464 856
rect 158632 800 159108 856
rect 159276 800 159660 856
rect 159828 800 160304 856
rect 160472 800 160948 856
rect 161116 800 161500 856
rect 161668 800 162144 856
rect 162312 800 162788 856
rect 162956 800 163340 856
rect 163508 800 163984 856
rect 164152 800 164628 856
rect 164796 800 165180 856
rect 165348 800 165824 856
rect 165992 800 166468 856
rect 166636 800 167020 856
rect 167188 800 167664 856
rect 167832 800 168308 856
rect 168476 800 168860 856
rect 169028 800 169504 856
rect 169672 800 170148 856
rect 170316 800 170700 856
rect 170868 800 171344 856
rect 171512 800 171988 856
rect 172156 800 172540 856
rect 172708 800 173184 856
rect 173352 800 173828 856
rect 173996 800 174380 856
rect 174548 800 175024 856
rect 175192 800 175668 856
rect 175836 800 176220 856
rect 176388 800 176864 856
rect 177032 800 177416 856
rect 177584 800 178060 856
rect 178228 800 178704 856
rect 178872 800 179256 856
rect 179424 800 179900 856
rect 180068 800 180544 856
rect 180712 800 181096 856
rect 181264 800 181740 856
rect 181908 800 182384 856
rect 182552 800 182936 856
rect 183104 800 183580 856
rect 183748 800 184224 856
rect 184392 800 184776 856
rect 184944 800 185420 856
rect 185588 800 186064 856
rect 186232 800 186616 856
rect 186784 800 187260 856
rect 187428 800 187904 856
rect 188072 800 188456 856
rect 188624 800 189100 856
rect 189268 800 189744 856
rect 189912 800 190296 856
rect 190464 800 190940 856
rect 191108 800 191584 856
rect 191752 800 192136 856
rect 192304 800 192780 856
rect 192948 800 193424 856
rect 193592 800 193976 856
rect 194144 800 194620 856
rect 194788 800 195172 856
rect 195340 800 195816 856
rect 195984 800 196460 856
rect 196628 800 197012 856
rect 197180 800 197656 856
rect 197824 800 198300 856
rect 198468 800 198852 856
rect 199020 800 199496 856
rect 199664 800 200140 856
rect 200308 800 200692 856
rect 200860 800 201336 856
rect 201504 800 201980 856
rect 202148 800 202532 856
rect 202700 800 203176 856
rect 203344 800 203820 856
rect 203988 800 204372 856
rect 204540 800 205016 856
rect 205184 800 205660 856
rect 205828 800 206212 856
rect 206380 800 206856 856
rect 207024 800 207500 856
rect 207668 800 208052 856
rect 208220 800 208696 856
rect 208864 800 209340 856
rect 209508 800 209892 856
rect 210060 800 210536 856
rect 210704 800 211180 856
rect 211348 800 211732 856
rect 211900 800 212376 856
rect 212544 800 212928 856
rect 213096 800 213572 856
rect 213740 800 214216 856
rect 214384 800 214768 856
rect 214936 800 215412 856
rect 215580 800 216056 856
rect 216224 800 216608 856
rect 216776 800 217252 856
rect 217420 800 217896 856
rect 218064 800 218448 856
rect 218616 800 219092 856
rect 219260 800 219736 856
rect 219904 800 220288 856
rect 220456 800 220932 856
rect 221100 800 221576 856
rect 221744 800 222128 856
rect 222296 800 222772 856
rect 222940 800 223416 856
rect 223584 800 223968 856
rect 224136 800 224612 856
rect 224780 800 225256 856
rect 225424 800 225808 856
rect 225976 800 226452 856
rect 226620 800 227096 856
rect 227264 800 227648 856
rect 227816 800 228292 856
rect 228460 800 228936 856
rect 229104 800 229488 856
rect 229656 800 230132 856
rect 230300 800 230684 856
rect 230852 800 231328 856
rect 231496 800 231972 856
rect 232140 800 232524 856
rect 232692 800 233168 856
rect 233336 800 233812 856
rect 233980 800 234364 856
rect 234532 800 235008 856
rect 235176 800 235652 856
rect 235820 800 236204 856
rect 236372 800 236848 856
rect 237016 800 237492 856
rect 237660 800 238044 856
rect 238212 800 238688 856
rect 238856 800 239332 856
rect 239500 800 239884 856
rect 240052 800 240528 856
rect 240696 800 241172 856
rect 241340 800 241724 856
rect 241892 800 242368 856
rect 242536 800 243012 856
rect 243180 800 243564 856
rect 243732 800 244208 856
rect 244376 800 244852 856
rect 245020 800 245404 856
rect 245572 800 246048 856
rect 246216 800 246692 856
rect 246860 800 247244 856
rect 247412 800 247888 856
rect 248056 800 248440 856
rect 248608 800 249084 856
rect 249252 800 249728 856
rect 249896 800 250280 856
rect 250448 800 250924 856
rect 251092 800 251568 856
rect 251736 800 252120 856
rect 252288 800 252764 856
rect 252932 800 253408 856
rect 253576 800 253960 856
rect 254128 800 254604 856
rect 254772 800 255248 856
rect 255416 800 255800 856
rect 255968 800 256444 856
rect 256612 800 257088 856
rect 257256 800 257640 856
rect 257808 800 258284 856
rect 258452 800 258928 856
rect 259096 800 259480 856
rect 259648 800 260124 856
rect 260292 800 260768 856
rect 260936 800 261320 856
rect 261488 800 261964 856
rect 262132 800 262608 856
rect 262776 800 263160 856
rect 263328 800 263804 856
rect 263972 800 264448 856
rect 264616 800 265000 856
rect 265168 800 265644 856
rect 265812 800 266196 856
rect 266364 800 266840 856
rect 267008 800 267484 856
rect 267652 800 268036 856
rect 268204 800 268680 856
rect 268848 800 269324 856
rect 269492 800 269876 856
rect 270044 800 270520 856
rect 270688 800 271164 856
rect 271332 800 271716 856
rect 271884 800 272360 856
rect 272528 800 273004 856
rect 273172 800 273556 856
rect 273724 800 274200 856
rect 274368 800 274844 856
rect 275012 800 275396 856
rect 275564 800 276040 856
rect 276208 800 276684 856
rect 276852 800 277236 856
rect 277404 800 277880 856
rect 278048 800 278524 856
rect 278692 800 279076 856
rect 279244 800 279720 856
rect 279888 800 280364 856
rect 280532 800 280916 856
rect 281084 800 281560 856
rect 281728 800 282204 856
rect 282372 800 282756 856
rect 282924 800 283400 856
rect 283568 800 283952 856
rect 284120 800 284596 856
rect 284764 800 285240 856
rect 285408 800 285792 856
rect 285960 800 286436 856
rect 286604 800 287080 856
rect 287248 800 287632 856
rect 287800 800 288276 856
rect 288444 800 288920 856
rect 289088 800 289472 856
rect 289640 800 290116 856
rect 290284 800 290760 856
rect 290928 800 291312 856
rect 291480 800 291956 856
rect 292124 800 292600 856
rect 292768 800 293152 856
rect 293320 800 293796 856
rect 293964 800 294440 856
rect 294608 800 294992 856
rect 295160 800 295636 856
rect 295804 800 296280 856
rect 296448 800 296832 856
rect 297000 800 297476 856
rect 297644 800 298120 856
rect 298288 800 298672 856
rect 298840 800 299316 856
<< obsm3 >>
rect 2391 851 296765 297601
<< metal4 >>
rect 3918 2128 4238 297616
rect 19278 2128 19598 297616
<< obsm4 >>
rect 34638 2128 296078 297616
<< labels >>
rlabel metal2 s 1016 299200 1072 300000 6 io_in[0]
port 1 nsew default input
rlabel metal2 s 79952 299200 80008 300000 6 io_in[10]
port 2 nsew default input
rlabel metal2 s 87772 299200 87828 300000 6 io_in[11]
port 3 nsew default input
rlabel metal2 s 95684 299200 95740 300000 6 io_in[12]
port 4 nsew default input
rlabel metal2 s 103596 299200 103652 300000 6 io_in[13]
port 5 nsew default input
rlabel metal2 s 111508 299200 111564 300000 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 119420 299200 119476 300000 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 127332 299200 127388 300000 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 135152 299200 135208 300000 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 143064 299200 143120 300000 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 150976 299200 151032 300000 6 io_in[19]
port 11 nsew default input
rlabel metal2 s 8836 299200 8892 300000 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 158888 299200 158944 300000 6 io_in[20]
port 13 nsew default input
rlabel metal2 s 166800 299200 166856 300000 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 174620 299200 174676 300000 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 182532 299200 182588 300000 6 io_in[23]
port 16 nsew default input
rlabel metal2 s 190444 299200 190500 300000 6 io_in[24]
port 17 nsew default input
rlabel metal2 s 198356 299200 198412 300000 6 io_in[25]
port 18 nsew default input
rlabel metal2 s 206268 299200 206324 300000 6 io_in[26]
port 19 nsew default input
rlabel metal2 s 214180 299200 214236 300000 6 io_in[27]
port 20 nsew default input
rlabel metal2 s 222000 299200 222056 300000 6 io_in[28]
port 21 nsew default input
rlabel metal2 s 229912 299200 229968 300000 6 io_in[29]
port 22 nsew default input
rlabel metal2 s 16748 299200 16804 300000 6 io_in[2]
port 23 nsew default input
rlabel metal2 s 237824 299200 237880 300000 6 io_in[30]
port 24 nsew default input
rlabel metal2 s 245736 299200 245792 300000 6 io_in[31]
port 25 nsew default input
rlabel metal2 s 253648 299200 253704 300000 6 io_in[32]
port 26 nsew default input
rlabel metal2 s 261468 299200 261524 300000 6 io_in[33]
port 27 nsew default input
rlabel metal2 s 269380 299200 269436 300000 6 io_in[34]
port 28 nsew default input
rlabel metal2 s 277292 299200 277348 300000 6 io_in[35]
port 29 nsew default input
rlabel metal2 s 285204 299200 285260 300000 6 io_in[36]
port 30 nsew default input
rlabel metal2 s 293116 299200 293172 300000 6 io_in[37]
port 31 nsew default input
rlabel metal2 s 24660 299200 24716 300000 6 io_in[3]
port 32 nsew default input
rlabel metal2 s 32572 299200 32628 300000 6 io_in[4]
port 33 nsew default input
rlabel metal2 s 40484 299200 40540 300000 6 io_in[5]
port 34 nsew default input
rlabel metal2 s 48304 299200 48360 300000 6 io_in[6]
port 35 nsew default input
rlabel metal2 s 56216 299200 56272 300000 6 io_in[7]
port 36 nsew default input
rlabel metal2 s 64128 299200 64184 300000 6 io_in[8]
port 37 nsew default input
rlabel metal2 s 72040 299200 72096 300000 6 io_in[9]
port 38 nsew default input
rlabel metal2 s 3592 299200 3648 300000 6 io_oeb[0]
port 39 nsew default output
rlabel metal2 s 82528 299200 82584 300000 6 io_oeb[10]
port 40 nsew default output
rlabel metal2 s 90440 299200 90496 300000 6 io_oeb[11]
port 41 nsew default output
rlabel metal2 s 98352 299200 98408 300000 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 106264 299200 106320 300000 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 114176 299200 114232 300000 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 121996 299200 122052 300000 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 129908 299200 129964 300000 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 137820 299200 137876 300000 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 145732 299200 145788 300000 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 153644 299200 153700 300000 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 11504 299200 11560 300000 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 161464 299200 161520 300000 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 169376 299200 169432 300000 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 177288 299200 177344 300000 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 185200 299200 185256 300000 6 io_oeb[23]
port 54 nsew default output
rlabel metal2 s 193112 299200 193168 300000 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 201024 299200 201080 300000 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 208844 299200 208900 300000 6 io_oeb[26]
port 57 nsew default output
rlabel metal2 s 216756 299200 216812 300000 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 224668 299200 224724 300000 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 232580 299200 232636 300000 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 19416 299200 19472 300000 6 io_oeb[2]
port 61 nsew default output
rlabel metal2 s 240492 299200 240548 300000 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 248312 299200 248368 300000 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 256224 299200 256280 300000 6 io_oeb[32]
port 64 nsew default output
rlabel metal2 s 264136 299200 264192 300000 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 272048 299200 272104 300000 6 io_oeb[34]
port 66 nsew default output
rlabel metal2 s 279960 299200 280016 300000 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 287780 299200 287836 300000 6 io_oeb[36]
port 68 nsew default output
rlabel metal2 s 295692 299200 295748 300000 6 io_oeb[37]
port 69 nsew default output
rlabel metal2 s 27328 299200 27384 300000 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 35148 299200 35204 300000 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 43060 299200 43116 300000 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 50972 299200 51028 300000 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 58884 299200 58940 300000 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 66796 299200 66852 300000 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 74616 299200 74672 300000 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 6260 299200 6316 300000 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 85196 299200 85252 300000 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 93108 299200 93164 300000 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 101020 299200 101076 300000 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 108840 299200 108896 300000 6 io_out[13]
port 81 nsew default output
rlabel metal2 s 116752 299200 116808 300000 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 124664 299200 124720 300000 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 132576 299200 132632 300000 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 140488 299200 140544 300000 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 148308 299200 148364 300000 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 156220 299200 156276 300000 6 io_out[19]
port 87 nsew default output
rlabel metal2 s 14172 299200 14228 300000 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 164132 299200 164188 300000 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 172044 299200 172100 300000 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 179956 299200 180012 300000 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 187776 299200 187832 300000 6 io_out[23]
port 92 nsew default output
rlabel metal2 s 195688 299200 195744 300000 6 io_out[24]
port 93 nsew default output
rlabel metal2 s 203600 299200 203656 300000 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 211512 299200 211568 300000 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 219424 299200 219480 300000 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 227336 299200 227392 300000 6 io_out[28]
port 97 nsew default output
rlabel metal2 s 235156 299200 235212 300000 6 io_out[29]
port 98 nsew default output
rlabel metal2 s 21992 299200 22048 300000 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 243068 299200 243124 300000 6 io_out[30]
port 100 nsew default output
rlabel metal2 s 250980 299200 251036 300000 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 258892 299200 258948 300000 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 266804 299200 266860 300000 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 274624 299200 274680 300000 6 io_out[34]
port 104 nsew default output
rlabel metal2 s 282536 299200 282592 300000 6 io_out[35]
port 105 nsew default output
rlabel metal2 s 290448 299200 290504 300000 6 io_out[36]
port 106 nsew default output
rlabel metal2 s 298360 299200 298416 300000 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 29904 299200 29960 300000 6 io_out[3]
port 108 nsew default output
rlabel metal2 s 37816 299200 37872 300000 6 io_out[4]
port 109 nsew default output
rlabel metal2 s 45728 299200 45784 300000 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 53640 299200 53696 300000 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 61460 299200 61516 300000 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 69372 299200 69428 300000 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 77284 299200 77340 300000 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 64864 0 64920 800 6 la_data_in[0]
port 115 nsew default input
rlabel metal2 s 248496 0 248552 800 6 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 250336 0 250392 800 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 252176 0 252232 800 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 254016 0 254072 800 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 255856 0 255912 800 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 257696 0 257752 800 6 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 259536 0 259592 800 6 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 261376 0 261432 800 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 263216 0 263272 800 6 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 265056 0 265112 800 6 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 83264 0 83320 800 6 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 266896 0 266952 800 6 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 268736 0 268792 800 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 270576 0 270632 800 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 272416 0 272472 800 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 274256 0 274312 800 6 la_data_in[114]
port 131 nsew default input
rlabel metal2 s 276096 0 276152 800 6 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 277936 0 277992 800 6 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 279776 0 279832 800 6 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 281616 0 281672 800 6 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 283456 0 283512 800 6 la_data_in[119]
port 136 nsew default input
rlabel metal2 s 85104 0 85160 800 6 la_data_in[11]
port 137 nsew default input
rlabel metal2 s 285296 0 285352 800 6 la_data_in[120]
port 138 nsew default input
rlabel metal2 s 287136 0 287192 800 6 la_data_in[121]
port 139 nsew default input
rlabel metal2 s 288976 0 289032 800 6 la_data_in[122]
port 140 nsew default input
rlabel metal2 s 290816 0 290872 800 6 la_data_in[123]
port 141 nsew default input
rlabel metal2 s 292656 0 292712 800 6 la_data_in[124]
port 142 nsew default input
rlabel metal2 s 294496 0 294552 800 6 la_data_in[125]
port 143 nsew default input
rlabel metal2 s 296336 0 296392 800 6 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 298176 0 298232 800 6 la_data_in[127]
port 145 nsew default input
rlabel metal2 s 86944 0 87000 800 6 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 88692 0 88748 800 6 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 90532 0 90588 800 6 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 92372 0 92428 800 6 la_data_in[15]
port 149 nsew default input
rlabel metal2 s 94212 0 94268 800 6 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 96052 0 96108 800 6 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 97892 0 97948 800 6 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 99732 0 99788 800 6 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 66704 0 66760 800 6 la_data_in[1]
port 154 nsew default input
rlabel metal2 s 101572 0 101628 800 6 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 103412 0 103468 800 6 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 105252 0 105308 800 6 la_data_in[22]
port 157 nsew default input
rlabel metal2 s 107092 0 107148 800 6 la_data_in[23]
port 158 nsew default input
rlabel metal2 s 108932 0 108988 800 6 la_data_in[24]
port 159 nsew default input
rlabel metal2 s 110772 0 110828 800 6 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 112612 0 112668 800 6 la_data_in[26]
port 161 nsew default input
rlabel metal2 s 114452 0 114508 800 6 la_data_in[27]
port 162 nsew default input
rlabel metal2 s 116292 0 116348 800 6 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 118132 0 118188 800 6 la_data_in[29]
port 164 nsew default input
rlabel metal2 s 68544 0 68600 800 6 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 119972 0 120028 800 6 la_data_in[30]
port 166 nsew default input
rlabel metal2 s 121812 0 121868 800 6 la_data_in[31]
port 167 nsew default input
rlabel metal2 s 123652 0 123708 800 6 la_data_in[32]
port 168 nsew default input
rlabel metal2 s 125492 0 125548 800 6 la_data_in[33]
port 169 nsew default input
rlabel metal2 s 127332 0 127388 800 6 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 129172 0 129228 800 6 la_data_in[35]
port 171 nsew default input
rlabel metal2 s 131012 0 131068 800 6 la_data_in[36]
port 172 nsew default input
rlabel metal2 s 132852 0 132908 800 6 la_data_in[37]
port 173 nsew default input
rlabel metal2 s 134692 0 134748 800 6 la_data_in[38]
port 174 nsew default input
rlabel metal2 s 136532 0 136588 800 6 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 70384 0 70440 800 6 la_data_in[3]
port 176 nsew default input
rlabel metal2 s 138372 0 138428 800 6 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 140212 0 140268 800 6 la_data_in[41]
port 178 nsew default input
rlabel metal2 s 141960 0 142016 800 6 la_data_in[42]
port 179 nsew default input
rlabel metal2 s 143800 0 143856 800 6 la_data_in[43]
port 180 nsew default input
rlabel metal2 s 145640 0 145696 800 6 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 147480 0 147536 800 6 la_data_in[45]
port 182 nsew default input
rlabel metal2 s 149320 0 149376 800 6 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 151160 0 151216 800 6 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 153000 0 153056 800 6 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 154840 0 154896 800 6 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 72224 0 72280 800 6 la_data_in[4]
port 187 nsew default input
rlabel metal2 s 156680 0 156736 800 6 la_data_in[50]
port 188 nsew default input
rlabel metal2 s 158520 0 158576 800 6 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 160360 0 160416 800 6 la_data_in[52]
port 190 nsew default input
rlabel metal2 s 162200 0 162256 800 6 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 164040 0 164096 800 6 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 165880 0 165936 800 6 la_data_in[55]
port 193 nsew default input
rlabel metal2 s 167720 0 167776 800 6 la_data_in[56]
port 194 nsew default input
rlabel metal2 s 169560 0 169616 800 6 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 171400 0 171456 800 6 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 173240 0 173296 800 6 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 74064 0 74120 800 6 la_data_in[5]
port 198 nsew default input
rlabel metal2 s 175080 0 175136 800 6 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 176920 0 176976 800 6 la_data_in[61]
port 200 nsew default input
rlabel metal2 s 178760 0 178816 800 6 la_data_in[62]
port 201 nsew default input
rlabel metal2 s 180600 0 180656 800 6 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 182440 0 182496 800 6 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 184280 0 184336 800 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 186120 0 186176 800 6 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 187960 0 188016 800 6 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 189800 0 189856 800 6 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 191640 0 191696 800 6 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 75904 0 75960 800 6 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 193480 0 193536 800 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 195228 0 195284 800 6 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 197068 0 197124 800 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 198908 0 198964 800 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 200748 0 200804 800 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 202588 0 202644 800 6 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 204428 0 204484 800 6 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 206268 0 206324 800 6 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 208108 0 208164 800 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 209948 0 210004 800 6 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 77744 0 77800 800 6 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 211788 0 211844 800 6 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 213628 0 213684 800 6 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 215468 0 215524 800 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 217308 0 217364 800 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 219148 0 219204 800 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 220988 0 221044 800 6 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 222828 0 222884 800 6 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 224668 0 224724 800 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 226508 0 226564 800 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 228348 0 228404 800 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 79584 0 79640 800 6 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 230188 0 230244 800 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 232028 0 232084 800 6 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 233868 0 233924 800 6 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 235708 0 235764 800 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 237548 0 237604 800 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 239388 0 239444 800 6 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 241228 0 241284 800 6 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 243068 0 243124 800 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 244908 0 244964 800 6 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 246748 0 246804 800 6 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 81424 0 81480 800 6 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 65508 0 65564 800 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 249140 0 249196 800 6 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 250980 0 251036 800 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 252820 0 252876 800 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 254660 0 254716 800 6 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 256500 0 256556 800 6 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 258340 0 258396 800 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 260180 0 260236 800 6 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 262020 0 262076 800 6 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 263860 0 263916 800 6 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 265700 0 265756 800 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 83816 0 83872 800 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 267540 0 267596 800 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 269380 0 269436 800 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 271220 0 271276 800 6 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 273060 0 273116 800 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 274900 0 274956 800 6 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 276740 0 276796 800 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 278580 0 278636 800 6 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 280420 0 280476 800 6 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 282260 0 282316 800 6 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 284008 0 284064 800 6 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 85656 0 85712 800 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 285848 0 285904 800 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 287688 0 287744 800 6 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 289528 0 289584 800 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 291368 0 291424 800 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 293208 0 293264 800 6 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 295048 0 295104 800 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 296888 0 296944 800 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 298728 0 298784 800 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 87496 0 87552 800 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 89336 0 89392 800 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 91176 0 91232 800 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 93016 0 93072 800 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 94856 0 94912 800 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 96696 0 96752 800 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 98536 0 98592 800 6 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 100376 0 100432 800 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 67348 0 67404 800 6 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 102216 0 102272 800 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 104056 0 104112 800 6 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 105896 0 105952 800 6 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 107736 0 107792 800 6 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 109576 0 109632 800 6 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 111416 0 111472 800 6 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 113256 0 113312 800 6 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 115096 0 115152 800 6 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 116936 0 116992 800 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 118776 0 118832 800 6 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 69188 0 69244 800 6 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 120616 0 120672 800 6 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 122456 0 122512 800 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 124204 0 124260 800 6 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 126044 0 126100 800 6 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 127884 0 127940 800 6 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 129724 0 129780 800 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 131564 0 131620 800 6 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 133404 0 133460 800 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 135244 0 135300 800 6 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 137084 0 137140 800 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 70936 0 70992 800 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 138924 0 138980 800 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 140764 0 140820 800 6 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 142604 0 142660 800 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 144444 0 144500 800 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 146284 0 146340 800 6 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 148124 0 148180 800 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 149964 0 150020 800 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 151804 0 151860 800 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 153644 0 153700 800 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 155484 0 155540 800 6 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 72776 0 72832 800 6 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 157324 0 157380 800 6 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 159164 0 159220 800 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 161004 0 161060 800 6 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 162844 0 162900 800 6 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 164684 0 164740 800 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 166524 0 166580 800 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 168364 0 168420 800 6 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 170204 0 170260 800 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 172044 0 172100 800 6 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 173884 0 173940 800 6 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 74616 0 74672 800 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 175724 0 175780 800 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 177472 0 177528 800 6 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 179312 0 179368 800 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 181152 0 181208 800 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 182992 0 183048 800 6 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 184832 0 184888 800 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 186672 0 186728 800 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 188512 0 188568 800 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 190352 0 190408 800 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 192192 0 192248 800 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 76456 0 76512 800 6 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 194032 0 194088 800 6 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 195872 0 195928 800 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 197712 0 197768 800 6 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 199552 0 199608 800 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 201392 0 201448 800 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 203232 0 203288 800 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 205072 0 205128 800 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 206912 0 206968 800 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 208752 0 208808 800 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 210592 0 210648 800 6 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 78296 0 78352 800 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 212432 0 212488 800 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 214272 0 214328 800 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 216112 0 216168 800 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 217952 0 218008 800 6 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 219792 0 219848 800 6 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 221632 0 221688 800 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 223472 0 223528 800 6 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 225312 0 225368 800 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 227152 0 227208 800 6 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 228992 0 229048 800 6 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 80136 0 80192 800 6 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 230740 0 230796 800 6 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 232580 0 232636 800 6 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 234420 0 234476 800 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 236260 0 236316 800 6 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 238100 0 238156 800 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 239940 0 239996 800 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 241780 0 241836 800 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 243620 0 243676 800 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 245460 0 245516 800 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 247300 0 247356 800 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 81976 0 82032 800 6 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 66060 0 66116 800 6 la_oen[0]
port 371 nsew default input
rlabel metal2 s 249784 0 249840 800 6 la_oen[100]
port 372 nsew default input
rlabel metal2 s 251624 0 251680 800 6 la_oen[101]
port 373 nsew default input
rlabel metal2 s 253464 0 253520 800 6 la_oen[102]
port 374 nsew default input
rlabel metal2 s 255304 0 255360 800 6 la_oen[103]
port 375 nsew default input
rlabel metal2 s 257144 0 257200 800 6 la_oen[104]
port 376 nsew default input
rlabel metal2 s 258984 0 259040 800 6 la_oen[105]
port 377 nsew default input
rlabel metal2 s 260824 0 260880 800 6 la_oen[106]
port 378 nsew default input
rlabel metal2 s 262664 0 262720 800 6 la_oen[107]
port 379 nsew default input
rlabel metal2 s 264504 0 264560 800 6 la_oen[108]
port 380 nsew default input
rlabel metal2 s 266252 0 266308 800 6 la_oen[109]
port 381 nsew default input
rlabel metal2 s 84460 0 84516 800 6 la_oen[10]
port 382 nsew default input
rlabel metal2 s 268092 0 268148 800 6 la_oen[110]
port 383 nsew default input
rlabel metal2 s 269932 0 269988 800 6 la_oen[111]
port 384 nsew default input
rlabel metal2 s 271772 0 271828 800 6 la_oen[112]
port 385 nsew default input
rlabel metal2 s 273612 0 273668 800 6 la_oen[113]
port 386 nsew default input
rlabel metal2 s 275452 0 275508 800 6 la_oen[114]
port 387 nsew default input
rlabel metal2 s 277292 0 277348 800 6 la_oen[115]
port 388 nsew default input
rlabel metal2 s 279132 0 279188 800 6 la_oen[116]
port 389 nsew default input
rlabel metal2 s 280972 0 281028 800 6 la_oen[117]
port 390 nsew default input
rlabel metal2 s 282812 0 282868 800 6 la_oen[118]
port 391 nsew default input
rlabel metal2 s 284652 0 284708 800 6 la_oen[119]
port 392 nsew default input
rlabel metal2 s 86300 0 86356 800 6 la_oen[11]
port 393 nsew default input
rlabel metal2 s 286492 0 286548 800 6 la_oen[120]
port 394 nsew default input
rlabel metal2 s 288332 0 288388 800 6 la_oen[121]
port 395 nsew default input
rlabel metal2 s 290172 0 290228 800 6 la_oen[122]
port 396 nsew default input
rlabel metal2 s 292012 0 292068 800 6 la_oen[123]
port 397 nsew default input
rlabel metal2 s 293852 0 293908 800 6 la_oen[124]
port 398 nsew default input
rlabel metal2 s 295692 0 295748 800 6 la_oen[125]
port 399 nsew default input
rlabel metal2 s 297532 0 297588 800 6 la_oen[126]
port 400 nsew default input
rlabel metal2 s 299372 0 299428 800 6 la_oen[127]
port 401 nsew default input
rlabel metal2 s 88140 0 88196 800 6 la_oen[12]
port 402 nsew default input
rlabel metal2 s 89980 0 90036 800 6 la_oen[13]
port 403 nsew default input
rlabel metal2 s 91820 0 91876 800 6 la_oen[14]
port 404 nsew default input
rlabel metal2 s 93660 0 93716 800 6 la_oen[15]
port 405 nsew default input
rlabel metal2 s 95500 0 95556 800 6 la_oen[16]
port 406 nsew default input
rlabel metal2 s 97340 0 97396 800 6 la_oen[17]
port 407 nsew default input
rlabel metal2 s 99180 0 99236 800 6 la_oen[18]
port 408 nsew default input
rlabel metal2 s 101020 0 101076 800 6 la_oen[19]
port 409 nsew default input
rlabel metal2 s 67900 0 67956 800 6 la_oen[1]
port 410 nsew default input
rlabel metal2 s 102860 0 102916 800 6 la_oen[20]
port 411 nsew default input
rlabel metal2 s 104700 0 104756 800 6 la_oen[21]
port 412 nsew default input
rlabel metal2 s 106448 0 106504 800 6 la_oen[22]
port 413 nsew default input
rlabel metal2 s 108288 0 108344 800 6 la_oen[23]
port 414 nsew default input
rlabel metal2 s 110128 0 110184 800 6 la_oen[24]
port 415 nsew default input
rlabel metal2 s 111968 0 112024 800 6 la_oen[25]
port 416 nsew default input
rlabel metal2 s 113808 0 113864 800 6 la_oen[26]
port 417 nsew default input
rlabel metal2 s 115648 0 115704 800 6 la_oen[27]
port 418 nsew default input
rlabel metal2 s 117488 0 117544 800 6 la_oen[28]
port 419 nsew default input
rlabel metal2 s 119328 0 119384 800 6 la_oen[29]
port 420 nsew default input
rlabel metal2 s 69740 0 69796 800 6 la_oen[2]
port 421 nsew default input
rlabel metal2 s 121168 0 121224 800 6 la_oen[30]
port 422 nsew default input
rlabel metal2 s 123008 0 123064 800 6 la_oen[31]
port 423 nsew default input
rlabel metal2 s 124848 0 124904 800 6 la_oen[32]
port 424 nsew default input
rlabel metal2 s 126688 0 126744 800 6 la_oen[33]
port 425 nsew default input
rlabel metal2 s 128528 0 128584 800 6 la_oen[34]
port 426 nsew default input
rlabel metal2 s 130368 0 130424 800 6 la_oen[35]
port 427 nsew default input
rlabel metal2 s 132208 0 132264 800 6 la_oen[36]
port 428 nsew default input
rlabel metal2 s 134048 0 134104 800 6 la_oen[37]
port 429 nsew default input
rlabel metal2 s 135888 0 135944 800 6 la_oen[38]
port 430 nsew default input
rlabel metal2 s 137728 0 137784 800 6 la_oen[39]
port 431 nsew default input
rlabel metal2 s 71580 0 71636 800 6 la_oen[3]
port 432 nsew default input
rlabel metal2 s 139568 0 139624 800 6 la_oen[40]
port 433 nsew default input
rlabel metal2 s 141408 0 141464 800 6 la_oen[41]
port 434 nsew default input
rlabel metal2 s 143248 0 143304 800 6 la_oen[42]
port 435 nsew default input
rlabel metal2 s 145088 0 145144 800 6 la_oen[43]
port 436 nsew default input
rlabel metal2 s 146928 0 146984 800 6 la_oen[44]
port 437 nsew default input
rlabel metal2 s 148768 0 148824 800 6 la_oen[45]
port 438 nsew default input
rlabel metal2 s 150608 0 150664 800 6 la_oen[46]
port 439 nsew default input
rlabel metal2 s 152448 0 152504 800 6 la_oen[47]
port 440 nsew default input
rlabel metal2 s 154288 0 154344 800 6 la_oen[48]
port 441 nsew default input
rlabel metal2 s 156128 0 156184 800 6 la_oen[49]
port 442 nsew default input
rlabel metal2 s 73420 0 73476 800 6 la_oen[4]
port 443 nsew default input
rlabel metal2 s 157968 0 158024 800 6 la_oen[50]
port 444 nsew default input
rlabel metal2 s 159716 0 159772 800 6 la_oen[51]
port 445 nsew default input
rlabel metal2 s 161556 0 161612 800 6 la_oen[52]
port 446 nsew default input
rlabel metal2 s 163396 0 163452 800 6 la_oen[53]
port 447 nsew default input
rlabel metal2 s 165236 0 165292 800 6 la_oen[54]
port 448 nsew default input
rlabel metal2 s 167076 0 167132 800 6 la_oen[55]
port 449 nsew default input
rlabel metal2 s 168916 0 168972 800 6 la_oen[56]
port 450 nsew default input
rlabel metal2 s 170756 0 170812 800 6 la_oen[57]
port 451 nsew default input
rlabel metal2 s 172596 0 172652 800 6 la_oen[58]
port 452 nsew default input
rlabel metal2 s 174436 0 174492 800 6 la_oen[59]
port 453 nsew default input
rlabel metal2 s 75260 0 75316 800 6 la_oen[5]
port 454 nsew default input
rlabel metal2 s 176276 0 176332 800 6 la_oen[60]
port 455 nsew default input
rlabel metal2 s 178116 0 178172 800 6 la_oen[61]
port 456 nsew default input
rlabel metal2 s 179956 0 180012 800 6 la_oen[62]
port 457 nsew default input
rlabel metal2 s 181796 0 181852 800 6 la_oen[63]
port 458 nsew default input
rlabel metal2 s 183636 0 183692 800 6 la_oen[64]
port 459 nsew default input
rlabel metal2 s 185476 0 185532 800 6 la_oen[65]
port 460 nsew default input
rlabel metal2 s 187316 0 187372 800 6 la_oen[66]
port 461 nsew default input
rlabel metal2 s 189156 0 189212 800 6 la_oen[67]
port 462 nsew default input
rlabel metal2 s 190996 0 191052 800 6 la_oen[68]
port 463 nsew default input
rlabel metal2 s 192836 0 192892 800 6 la_oen[69]
port 464 nsew default input
rlabel metal2 s 77100 0 77156 800 6 la_oen[6]
port 465 nsew default input
rlabel metal2 s 194676 0 194732 800 6 la_oen[70]
port 466 nsew default input
rlabel metal2 s 196516 0 196572 800 6 la_oen[71]
port 467 nsew default input
rlabel metal2 s 198356 0 198412 800 6 la_oen[72]
port 468 nsew default input
rlabel metal2 s 200196 0 200252 800 6 la_oen[73]
port 469 nsew default input
rlabel metal2 s 202036 0 202092 800 6 la_oen[74]
port 470 nsew default input
rlabel metal2 s 203876 0 203932 800 6 la_oen[75]
port 471 nsew default input
rlabel metal2 s 205716 0 205772 800 6 la_oen[76]
port 472 nsew default input
rlabel metal2 s 207556 0 207612 800 6 la_oen[77]
port 473 nsew default input
rlabel metal2 s 209396 0 209452 800 6 la_oen[78]
port 474 nsew default input
rlabel metal2 s 211236 0 211292 800 6 la_oen[79]
port 475 nsew default input
rlabel metal2 s 78940 0 78996 800 6 la_oen[7]
port 476 nsew default input
rlabel metal2 s 212984 0 213040 800 6 la_oen[80]
port 477 nsew default input
rlabel metal2 s 214824 0 214880 800 6 la_oen[81]
port 478 nsew default input
rlabel metal2 s 216664 0 216720 800 6 la_oen[82]
port 479 nsew default input
rlabel metal2 s 218504 0 218560 800 6 la_oen[83]
port 480 nsew default input
rlabel metal2 s 220344 0 220400 800 6 la_oen[84]
port 481 nsew default input
rlabel metal2 s 222184 0 222240 800 6 la_oen[85]
port 482 nsew default input
rlabel metal2 s 224024 0 224080 800 6 la_oen[86]
port 483 nsew default input
rlabel metal2 s 225864 0 225920 800 6 la_oen[87]
port 484 nsew default input
rlabel metal2 s 227704 0 227760 800 6 la_oen[88]
port 485 nsew default input
rlabel metal2 s 229544 0 229600 800 6 la_oen[89]
port 486 nsew default input
rlabel metal2 s 80780 0 80836 800 6 la_oen[8]
port 487 nsew default input
rlabel metal2 s 231384 0 231440 800 6 la_oen[90]
port 488 nsew default input
rlabel metal2 s 233224 0 233280 800 6 la_oen[91]
port 489 nsew default input
rlabel metal2 s 235064 0 235120 800 6 la_oen[92]
port 490 nsew default input
rlabel metal2 s 236904 0 236960 800 6 la_oen[93]
port 491 nsew default input
rlabel metal2 s 238744 0 238800 800 6 la_oen[94]
port 492 nsew default input
rlabel metal2 s 240584 0 240640 800 6 la_oen[95]
port 493 nsew default input
rlabel metal2 s 242424 0 242480 800 6 la_oen[96]
port 494 nsew default input
rlabel metal2 s 244264 0 244320 800 6 la_oen[97]
port 495 nsew default input
rlabel metal2 s 246104 0 246160 800 6 la_oen[98]
port 496 nsew default input
rlabel metal2 s 247944 0 248000 800 6 la_oen[99]
port 497 nsew default input
rlabel metal2 s 82620 0 82676 800 6 la_oen[9]
port 498 nsew default input
rlabel metal2 s 4 0 60 800 6 wb_clk_i
port 499 nsew default input
rlabel metal2 s 556 0 612 800 6 wb_rst_i
port 500 nsew default input
rlabel metal2 s 1200 0 1256 800 6 wbs_ack_o
port 501 nsew default output
rlabel metal2 s 3592 0 3648 800 6 wbs_adr_i[0]
port 502 nsew default input
rlabel metal2 s 24476 0 24532 800 6 wbs_adr_i[10]
port 503 nsew default input
rlabel metal2 s 26316 0 26372 800 6 wbs_adr_i[11]
port 504 nsew default input
rlabel metal2 s 28156 0 28212 800 6 wbs_adr_i[12]
port 505 nsew default input
rlabel metal2 s 29996 0 30052 800 6 wbs_adr_i[13]
port 506 nsew default input
rlabel metal2 s 31836 0 31892 800 6 wbs_adr_i[14]
port 507 nsew default input
rlabel metal2 s 33676 0 33732 800 6 wbs_adr_i[15]
port 508 nsew default input
rlabel metal2 s 35424 0 35480 800 6 wbs_adr_i[16]
port 509 nsew default input
rlabel metal2 s 37264 0 37320 800 6 wbs_adr_i[17]
port 510 nsew default input
rlabel metal2 s 39104 0 39160 800 6 wbs_adr_i[18]
port 511 nsew default input
rlabel metal2 s 40944 0 41000 800 6 wbs_adr_i[19]
port 512 nsew default input
rlabel metal2 s 6076 0 6132 800 6 wbs_adr_i[1]
port 513 nsew default input
rlabel metal2 s 42784 0 42840 800 6 wbs_adr_i[20]
port 514 nsew default input
rlabel metal2 s 44624 0 44680 800 6 wbs_adr_i[21]
port 515 nsew default input
rlabel metal2 s 46464 0 46520 800 6 wbs_adr_i[22]
port 516 nsew default input
rlabel metal2 s 48304 0 48360 800 6 wbs_adr_i[23]
port 517 nsew default input
rlabel metal2 s 50144 0 50200 800 6 wbs_adr_i[24]
port 518 nsew default input
rlabel metal2 s 51984 0 52040 800 6 wbs_adr_i[25]
port 519 nsew default input
rlabel metal2 s 53824 0 53880 800 6 wbs_adr_i[26]
port 520 nsew default input
rlabel metal2 s 55664 0 55720 800 6 wbs_adr_i[27]
port 521 nsew default input
rlabel metal2 s 57504 0 57560 800 6 wbs_adr_i[28]
port 522 nsew default input
rlabel metal2 s 59344 0 59400 800 6 wbs_adr_i[29]
port 523 nsew default input
rlabel metal2 s 8560 0 8616 800 6 wbs_adr_i[2]
port 524 nsew default input
rlabel metal2 s 61184 0 61240 800 6 wbs_adr_i[30]
port 525 nsew default input
rlabel metal2 s 63024 0 63080 800 6 wbs_adr_i[31]
port 526 nsew default input
rlabel metal2 s 10952 0 11008 800 6 wbs_adr_i[3]
port 527 nsew default input
rlabel metal2 s 13436 0 13492 800 6 wbs_adr_i[4]
port 528 nsew default input
rlabel metal2 s 15276 0 15332 800 6 wbs_adr_i[5]
port 529 nsew default input
rlabel metal2 s 17116 0 17172 800 6 wbs_adr_i[6]
port 530 nsew default input
rlabel metal2 s 18956 0 19012 800 6 wbs_adr_i[7]
port 531 nsew default input
rlabel metal2 s 20796 0 20852 800 6 wbs_adr_i[8]
port 532 nsew default input
rlabel metal2 s 22636 0 22692 800 6 wbs_adr_i[9]
port 533 nsew default input
rlabel metal2 s 1752 0 1808 800 6 wbs_cyc_i
port 534 nsew default input
rlabel metal2 s 4236 0 4292 800 6 wbs_dat_i[0]
port 535 nsew default input
rlabel metal2 s 25028 0 25084 800 6 wbs_dat_i[10]
port 536 nsew default input
rlabel metal2 s 26868 0 26924 800 6 wbs_dat_i[11]
port 537 nsew default input
rlabel metal2 s 28708 0 28764 800 6 wbs_dat_i[12]
port 538 nsew default input
rlabel metal2 s 30548 0 30604 800 6 wbs_dat_i[13]
port 539 nsew default input
rlabel metal2 s 32388 0 32444 800 6 wbs_dat_i[14]
port 540 nsew default input
rlabel metal2 s 34228 0 34284 800 6 wbs_dat_i[15]
port 541 nsew default input
rlabel metal2 s 36068 0 36124 800 6 wbs_dat_i[16]
port 542 nsew default input
rlabel metal2 s 37908 0 37964 800 6 wbs_dat_i[17]
port 543 nsew default input
rlabel metal2 s 39748 0 39804 800 6 wbs_dat_i[18]
port 544 nsew default input
rlabel metal2 s 41588 0 41644 800 6 wbs_dat_i[19]
port 545 nsew default input
rlabel metal2 s 6720 0 6776 800 6 wbs_dat_i[1]
port 546 nsew default input
rlabel metal2 s 43428 0 43484 800 6 wbs_dat_i[20]
port 547 nsew default input
rlabel metal2 s 45268 0 45324 800 6 wbs_dat_i[21]
port 548 nsew default input
rlabel metal2 s 47108 0 47164 800 6 wbs_dat_i[22]
port 549 nsew default input
rlabel metal2 s 48948 0 49004 800 6 wbs_dat_i[23]
port 550 nsew default input
rlabel metal2 s 50788 0 50844 800 6 wbs_dat_i[24]
port 551 nsew default input
rlabel metal2 s 52628 0 52684 800 6 wbs_dat_i[25]
port 552 nsew default input
rlabel metal2 s 54468 0 54524 800 6 wbs_dat_i[26]
port 553 nsew default input
rlabel metal2 s 56308 0 56364 800 6 wbs_dat_i[27]
port 554 nsew default input
rlabel metal2 s 58148 0 58204 800 6 wbs_dat_i[28]
port 555 nsew default input
rlabel metal2 s 59988 0 60044 800 6 wbs_dat_i[29]
port 556 nsew default input
rlabel metal2 s 9112 0 9168 800 6 wbs_dat_i[2]
port 557 nsew default input
rlabel metal2 s 61828 0 61884 800 6 wbs_dat_i[30]
port 558 nsew default input
rlabel metal2 s 63668 0 63724 800 6 wbs_dat_i[31]
port 559 nsew default input
rlabel metal2 s 11596 0 11652 800 6 wbs_dat_i[3]
port 560 nsew default input
rlabel metal2 s 14080 0 14136 800 6 wbs_dat_i[4]
port 561 nsew default input
rlabel metal2 s 15920 0 15976 800 6 wbs_dat_i[5]
port 562 nsew default input
rlabel metal2 s 17668 0 17724 800 6 wbs_dat_i[6]
port 563 nsew default input
rlabel metal2 s 19508 0 19564 800 6 wbs_dat_i[7]
port 564 nsew default input
rlabel metal2 s 21348 0 21404 800 6 wbs_dat_i[8]
port 565 nsew default input
rlabel metal2 s 23188 0 23244 800 6 wbs_dat_i[9]
port 566 nsew default input
rlabel metal2 s 4880 0 4936 800 6 wbs_dat_o[0]
port 567 nsew default output
rlabel metal2 s 25672 0 25728 800 6 wbs_dat_o[10]
port 568 nsew default output
rlabel metal2 s 27512 0 27568 800 6 wbs_dat_o[11]
port 569 nsew default output
rlabel metal2 s 29352 0 29408 800 6 wbs_dat_o[12]
port 570 nsew default output
rlabel metal2 s 31192 0 31248 800 6 wbs_dat_o[13]
port 571 nsew default output
rlabel metal2 s 33032 0 33088 800 6 wbs_dat_o[14]
port 572 nsew default output
rlabel metal2 s 34872 0 34928 800 6 wbs_dat_o[15]
port 573 nsew default output
rlabel metal2 s 36712 0 36768 800 6 wbs_dat_o[16]
port 574 nsew default output
rlabel metal2 s 38552 0 38608 800 6 wbs_dat_o[17]
port 575 nsew default output
rlabel metal2 s 40392 0 40448 800 6 wbs_dat_o[18]
port 576 nsew default output
rlabel metal2 s 42232 0 42288 800 6 wbs_dat_o[19]
port 577 nsew default output
rlabel metal2 s 7272 0 7328 800 6 wbs_dat_o[1]
port 578 nsew default output
rlabel metal2 s 44072 0 44128 800 6 wbs_dat_o[20]
port 579 nsew default output
rlabel metal2 s 45912 0 45968 800 6 wbs_dat_o[21]
port 580 nsew default output
rlabel metal2 s 47752 0 47808 800 6 wbs_dat_o[22]
port 581 nsew default output
rlabel metal2 s 49592 0 49648 800 6 wbs_dat_o[23]
port 582 nsew default output
rlabel metal2 s 51432 0 51488 800 6 wbs_dat_o[24]
port 583 nsew default output
rlabel metal2 s 53180 0 53236 800 6 wbs_dat_o[25]
port 584 nsew default output
rlabel metal2 s 55020 0 55076 800 6 wbs_dat_o[26]
port 585 nsew default output
rlabel metal2 s 56860 0 56916 800 6 wbs_dat_o[27]
port 586 nsew default output
rlabel metal2 s 58700 0 58756 800 6 wbs_dat_o[28]
port 587 nsew default output
rlabel metal2 s 60540 0 60596 800 6 wbs_dat_o[29]
port 588 nsew default output
rlabel metal2 s 9756 0 9812 800 6 wbs_dat_o[2]
port 589 nsew default output
rlabel metal2 s 62380 0 62436 800 6 wbs_dat_o[30]
port 590 nsew default output
rlabel metal2 s 64220 0 64276 800 6 wbs_dat_o[31]
port 591 nsew default output
rlabel metal2 s 12240 0 12296 800 6 wbs_dat_o[3]
port 592 nsew default output
rlabel metal2 s 14632 0 14688 800 6 wbs_dat_o[4]
port 593 nsew default output
rlabel metal2 s 16472 0 16528 800 6 wbs_dat_o[5]
port 594 nsew default output
rlabel metal2 s 18312 0 18368 800 6 wbs_dat_o[6]
port 595 nsew default output
rlabel metal2 s 20152 0 20208 800 6 wbs_dat_o[7]
port 596 nsew default output
rlabel metal2 s 21992 0 22048 800 6 wbs_dat_o[8]
port 597 nsew default output
rlabel metal2 s 23832 0 23888 800 6 wbs_dat_o[9]
port 598 nsew default output
rlabel metal2 s 5432 0 5488 800 6 wbs_sel_i[0]
port 599 nsew default input
rlabel metal2 s 7916 0 7972 800 6 wbs_sel_i[1]
port 600 nsew default input
rlabel metal2 s 10400 0 10456 800 6 wbs_sel_i[2]
port 601 nsew default input
rlabel metal2 s 12792 0 12848 800 6 wbs_sel_i[3]
port 602 nsew default input
rlabel metal2 s 2396 0 2452 800 6 wbs_stb_i
port 603 nsew default input
rlabel metal2 s 3040 0 3096 800 6 wbs_we_i
port 604 nsew default input
rlabel metal4 s 3918 2128 4238 297616 6 VPWR
port 605 nsew power input
rlabel metal4 s 19278 2128 19598 297616 6 VGND
port 606 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 299432 300000
string LEFview TRUE
<< end >>
