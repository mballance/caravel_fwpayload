magic
tech sky130A
magscale 1 2
timestamp 1608061857
<< locali >>
rect 364533 676243 364567 685797
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 364533 608651 364567 618205
rect 429393 601715 429427 608549
rect 559113 601715 559147 608549
rect 364625 589339 364659 598893
rect 429577 589339 429611 598893
rect 559297 589339 559331 598893
rect 247969 578595 248003 579309
rect 254225 578663 254259 579309
rect 292129 579139 292163 579309
rect 415685 578527 415719 579309
rect 428381 578459 428415 579309
rect 441077 578391 441111 579309
rect 453589 578323 453623 579309
rect 455797 578255 455831 579309
rect 318935 338045 319085 338079
rect 96111 337977 96261 338011
rect 115431 337977 115581 338011
rect 134751 337977 134901 338011
rect 154071 337977 154221 338011
rect 173391 337977 173541 338011
rect 192711 337977 192861 338011
rect 212031 337977 212181 338011
rect 96295 337841 96445 337875
rect 115615 337841 115765 337875
rect 134935 337841 135085 337875
rect 154255 337841 154405 337875
rect 173575 337841 173725 337875
rect 192895 337841 193045 337875
rect 212215 337841 212365 337875
rect 302191 337773 302283 337807
rect 302249 337739 302283 337773
rect 230489 337705 230707 337739
rect 96387 337569 96537 337603
rect 115707 337569 115857 337603
rect 135027 337569 135177 337603
rect 154347 337569 154497 337603
rect 173667 337569 173817 337603
rect 192987 337569 193137 337603
rect 212307 337569 212457 337603
rect 230489 337535 230523 337705
rect 230673 337671 230707 337705
rect 96295 337501 96445 337535
rect 115615 337501 115765 337535
rect 134935 337501 135085 337535
rect 154255 337501 154405 337535
rect 173575 337501 173725 337535
rect 192895 337501 193045 337535
rect 212215 337501 212365 337535
rect 230673 337637 231225 337671
rect 230581 337535 230615 337637
rect 234445 337467 234479 337637
rect 241529 337535 241563 337705
rect 96203 337433 96353 337467
rect 115523 337433 115673 337467
rect 134843 337433 134993 337467
rect 154163 337433 154313 337467
rect 173483 337433 173633 337467
rect 192803 337433 192953 337467
rect 212123 337433 212273 337467
rect 259745 337399 259779 337637
rect 115431 337365 115857 337399
rect 134751 337365 135177 337399
rect 154071 337365 154497 337399
rect 173391 337365 173817 337399
rect 192711 337365 193137 337399
rect 212031 337365 212457 337399
rect 303997 337195 304031 337773
rect 315497 337331 315531 338045
rect 318935 337909 318993 337943
rect 318843 337773 318993 337807
rect 327089 337739 327123 338113
rect 318935 337569 318993 337603
rect 318843 337433 319085 337467
rect 115615 337161 115857 337195
rect 326353 337195 326387 337297
rect 115523 337093 115765 337127
rect 134843 337093 135085 337127
rect 154163 337093 154313 337127
rect 173483 337093 173633 337127
rect 192803 337093 192953 337127
rect 212123 337093 212273 337127
rect 134751 337025 134993 337059
rect 154071 337025 154405 337059
rect 173391 337025 173725 337059
rect 192711 337025 193045 337059
rect 212031 337025 212365 337059
rect 334725 336787 334759 337365
rect 335829 337059 335863 337501
rect 335921 337399 335955 337841
rect 336013 337671 336047 337841
rect 336657 337739 336691 338113
rect 346409 337739 346443 338657
rect 372721 337807 372755 338045
rect 344293 337637 344661 337671
rect 344293 337535 344327 337637
rect 336197 336923 336231 337365
rect 340797 337127 340831 337365
rect 340613 336787 340647 337025
rect 340889 336855 340923 337365
rect 341717 337263 341751 337501
rect 342821 337195 342855 337501
rect 345581 336923 345615 337365
rect 345857 336991 345891 337161
rect 354045 336991 354079 337365
rect 364993 337195 365027 337637
rect 365119 337501 365269 337535
rect 365361 337467 365395 337569
rect 369869 337195 369903 337365
rect 374561 337195 374595 337433
rect 374653 336991 374687 337909
rect 412465 337739 412499 338045
rect 430037 337739 430071 337977
rect 414121 337399 414155 337705
rect 432521 337535 432555 338045
rect 432613 337399 432647 337773
rect 423045 336991 423079 337229
rect 345523 336821 345765 336855
rect 429301 336787 429335 337093
rect 431417 337059 431451 337161
rect 432705 336991 432739 337637
rect 434085 337127 434119 337977
rect 442273 337943 442307 338045
rect 442365 337943 442399 338113
rect 483155 338045 483247 338079
rect 483213 338011 483247 338045
rect 434303 337841 434453 337875
rect 434545 337739 434579 337909
rect 432429 336855 432463 336889
rect 436109 336855 436143 337433
rect 432429 336821 432613 336855
rect 340613 336753 340797 336787
rect 341015 336753 341165 336787
rect 437305 336787 437339 337637
rect 444389 337603 444423 337977
rect 449449 337671 449483 337841
rect 452025 337807 452059 337977
rect 455889 337807 455923 337977
rect 437489 337501 437673 337535
rect 437489 337195 437523 337501
rect 451933 337467 451967 337773
rect 437581 336855 437615 337161
rect 437523 336821 437615 336855
rect 445769 336855 445803 337365
rect 450369 336855 450403 337365
rect 456717 336787 456751 337841
rect 461501 337671 461535 337909
rect 461409 337331 461443 337637
rect 437305 336753 437397 336787
rect 463709 337331 463743 337841
rect 466377 337331 466411 337909
rect 483155 337909 483305 337943
rect 459017 336719 459051 337297
rect 466193 336855 466227 337297
rect 469229 337263 469263 337909
rect 483155 337773 483305 337807
rect 483155 337637 483305 337671
rect 483063 337433 483213 337467
rect 466319 337229 466411 337263
rect 466377 336923 466411 337229
rect 284401 335223 284435 336685
rect 250177 328491 250211 334441
rect 259837 318835 259871 328389
rect 262689 317475 262723 322269
rect 265265 317475 265299 318869
rect 266645 318835 266679 321589
rect 267749 318835 267783 321589
rect 288817 319107 288851 336685
rect 302525 328491 302559 334713
rect 327273 327131 327307 336685
rect 299857 317475 299891 327029
rect 339785 318835 339819 336685
rect 341349 318835 341383 328389
rect 358737 318835 358771 328389
rect 421205 327131 421239 336685
rect 466285 336651 466319 336889
rect 469597 336719 469631 336753
rect 469447 336685 469631 336719
rect 359197 317747 359231 327029
rect 470609 318835 470643 328389
rect 244473 309179 244507 311797
rect 236285 299523 236319 309077
rect 259653 299591 259687 309077
rect 262689 306391 262723 315945
rect 265265 299523 265299 309077
rect 266645 296735 266679 298129
rect 272165 296735 272199 314585
rect 273453 301563 273487 309281
rect 284585 306391 284619 311865
rect 285965 306459 285999 311865
rect 251465 289867 251499 294661
rect 272165 285719 272199 295273
rect 288725 290003 288759 311933
rect 310897 307887 310931 311933
rect 310713 298163 310747 307717
rect 295533 287079 295567 288473
rect 236285 270555 236319 280109
rect 239137 270555 239171 280109
rect 251465 270555 251499 280109
rect 259561 273071 259595 280109
rect 266737 276063 266771 285617
rect 296821 276063 296855 286977
rect 310897 282795 310931 293029
rect 323317 288507 323351 299421
rect 324697 289867 324731 299421
rect 327273 298163 327307 302141
rect 337025 298231 337059 307717
rect 339877 299931 339911 309077
rect 341165 299523 341199 309077
rect 358737 307819 358771 317373
rect 372721 309179 372755 318733
rect 386797 302107 386831 315945
rect 421205 307819 421239 317373
rect 460213 307819 460247 317373
rect 470609 299523 470643 309077
rect 337209 292451 337243 298061
rect 325893 278783 325927 280177
rect 236285 251243 236319 260797
rect 239137 251243 239171 260797
rect 250085 259471 250119 269025
rect 266645 260831 266679 274601
rect 310897 263483 310931 278681
rect 330125 260899 330159 273921
rect 336933 270555 336967 280109
rect 337117 278783 337151 282897
rect 341165 280211 341199 289765
rect 358737 280279 358771 298061
rect 359105 288439 359139 298061
rect 372721 289867 372755 299421
rect 375665 289867 375699 299421
rect 386797 282795 386831 293029
rect 421205 288439 421239 298061
rect 460029 288439 460063 298061
rect 470609 280211 470643 289765
rect 372721 270555 372755 280109
rect 377137 270555 377171 280109
rect 341165 260899 341199 270453
rect 386797 263483 386831 278681
rect 460121 273139 460155 280109
rect 463801 270555 463835 275281
rect 460029 260967 460063 270453
rect 470609 260899 470643 270453
rect 250177 251107 250211 259301
rect 251465 251243 251499 260797
rect 259561 253759 259595 260797
rect 259561 244171 259595 251141
rect 265357 248251 265391 255901
rect 270693 240227 270727 260797
rect 272533 249747 272567 258009
rect 310897 251311 310931 256037
rect 284677 240159 284711 249713
rect 262597 226355 262631 235909
rect 270693 233835 270727 238697
rect 285965 234515 285999 244953
rect 288909 236011 288943 245565
rect 310713 241519 310747 251141
rect 299489 231863 299523 241417
rect 327181 240227 327215 253929
rect 336933 249815 336967 260797
rect 337117 241587 337151 254609
rect 358737 240159 358771 259369
rect 372721 251243 372755 260797
rect 377137 251243 377171 260797
rect 463709 251243 463743 260797
rect 367017 241519 367051 251141
rect 470609 241519 470643 251141
rect 323409 231795 323443 234685
rect 324605 231795 324639 240057
rect 272073 220779 272107 229041
rect 310805 222207 310839 231761
rect 327181 230571 327215 240057
rect 337117 230503 337151 234617
rect 290105 208403 290139 217957
rect 291669 204051 291703 214557
rect 299489 212551 299523 222105
rect 358737 220847 358771 230401
rect 341165 215271 341199 220745
rect 310805 202895 310839 212449
rect 250085 186303 250119 200073
rect 265173 195279 265207 200073
rect 272349 193171 272383 201433
rect 299489 193239 299523 202793
rect 336933 193239 336967 202793
rect 266645 186303 266679 191777
rect 259653 173995 259687 179537
rect 284677 171139 284711 180761
rect 288817 179435 288851 191777
rect 290013 179435 290047 188649
rect 294337 179435 294371 184229
rect 299857 183583 299891 188445
rect 306849 183583 306883 188445
rect 367017 183583 367051 193137
rect 285965 161483 285999 171037
rect 288817 167059 288851 176613
rect 294429 168419 294463 177973
rect 299857 171139 299891 180761
rect 301053 171139 301087 180761
rect 302617 171139 302651 180761
rect 337117 172567 337151 183481
rect 460121 176511 460155 183481
rect 330125 162979 330159 172465
rect 232329 133943 232363 143497
rect 259653 142171 259687 154173
rect 272165 148971 272199 157981
rect 232329 114563 232363 124117
rect 239137 115991 239171 125545
rect 249993 114563 250027 124117
rect 251465 115991 251499 125545
rect 259837 124219 259871 142001
rect 270693 139995 270727 144857
rect 272441 135235 272475 143497
rect 286057 140811 286091 158661
rect 294337 149107 294371 158661
rect 310805 147611 310839 153153
rect 330125 151827 330159 161381
rect 372813 157335 372847 164169
rect 421205 153255 421239 162809
rect 460121 161483 460155 166957
rect 341165 144891 341199 153153
rect 360209 144891 360243 147713
rect 265265 124219 265299 133841
rect 288633 131155 288667 140709
rect 289921 132447 289955 138057
rect 270693 120683 270727 125545
rect 272441 114563 272475 124117
rect 291485 122723 291519 131053
rect 294429 129795 294463 139349
rect 295533 131155 295567 140709
rect 323317 133943 323351 143497
rect 324605 132515 324639 143497
rect 330125 137955 330159 143497
rect 367017 135303 367051 144857
rect 372721 135303 372755 138125
rect 377137 135303 377171 140029
rect 296913 121499 296947 131053
rect 299857 114563 299891 124117
rect 306849 113271 306883 124117
rect 324697 113203 324731 122757
rect 337209 114563 337243 132413
rect 358737 125647 358771 135201
rect 421205 133943 421239 143497
rect 460121 142239 460155 151725
rect 463709 144959 463743 147713
rect 460121 132515 460155 142069
rect 339785 118643 339819 125545
rect 341165 118643 341199 125545
rect 247233 106335 247267 109021
rect 232329 95251 232363 104805
rect 251465 96679 251499 106233
rect 265265 103547 265299 113101
rect 232329 75939 232363 85493
rect 236285 77435 236319 86921
rect 247141 85595 247175 95149
rect 262781 92531 262815 102085
rect 266829 96475 266863 103445
rect 267933 93891 267967 103445
rect 270693 101371 270727 106233
rect 284677 103547 284711 113101
rect 291577 103615 291611 113101
rect 294337 102187 294371 109701
rect 296821 103547 296855 113101
rect 325985 104907 326019 106301
rect 327181 104907 327215 114461
rect 341165 106335 341199 115889
rect 367017 106335 367051 115889
rect 421205 114563 421239 124117
rect 470609 106335 470643 115889
rect 291669 92531 291703 102085
rect 295625 93891 295659 103445
rect 301145 93891 301179 103445
rect 306849 93891 306883 103445
rect 251465 77299 251499 86921
rect 262689 75939 262723 88961
rect 265173 84303 265207 88961
rect 310805 85595 310839 95149
rect 324605 93891 324639 103445
rect 291577 84235 291611 85561
rect 265357 74579 265391 84133
rect 239137 67643 239171 70465
rect 244473 67643 244507 70465
rect 270785 67643 270819 80733
rect 272257 74579 272291 84133
rect 232329 56627 232363 66181
rect 236285 56627 236319 66181
rect 239045 56627 239079 58021
rect 250085 57987 250119 67541
rect 272257 67099 272291 67677
rect 284677 66283 284711 84133
rect 285965 66283 285999 84133
rect 265173 57919 265207 62645
rect 270785 56627 270819 66181
rect 239137 48331 239171 53193
rect 236285 38675 236319 48229
rect 244565 48195 244599 56525
rect 273453 50983 273487 66181
rect 288725 64923 288759 82773
rect 299857 75939 299891 85493
rect 317705 75939 317739 88349
rect 324697 76007 324731 85493
rect 330125 77299 330159 102085
rect 339785 95251 339819 104737
rect 341165 95251 341199 104805
rect 386521 99331 386555 106233
rect 336933 75939 336967 86921
rect 337209 77299 337243 86921
rect 341073 77299 341107 90389
rect 360301 89675 360335 96577
rect 367017 87023 367051 96577
rect 421205 87023 421239 104805
rect 470609 87023 470643 96577
rect 358737 75939 358771 85493
rect 310805 66351 310839 75837
rect 324605 66351 324639 75837
rect 377137 67643 377171 70465
rect 386613 67643 386647 77197
rect 421205 75939 421239 85493
rect 470609 67643 470643 77197
rect 236285 31671 236319 38505
rect 239045 29019 239079 42041
rect 244565 37315 244599 46869
rect 236377 22763 236411 28917
rect 259745 27659 259779 37213
rect 262781 35955 262815 45509
rect 273545 38675 273579 48229
rect 294245 46971 294279 64821
rect 310805 60027 310839 66181
rect 299673 45611 299707 56525
rect 301053 46971 301087 56525
rect 323317 48331 323351 66181
rect 324605 61387 324639 66181
rect 330125 56627 330159 66181
rect 336933 56627 336967 66181
rect 324789 46971 324823 56525
rect 337301 47039 337335 56525
rect 339785 48331 339819 57885
rect 358645 56627 358679 66181
rect 357541 46971 357575 56457
rect 367017 48331 367051 66181
rect 375665 61999 375699 67541
rect 421205 56627 421239 66181
rect 460029 48331 460063 57885
rect 470609 48331 470643 57885
rect 267841 28611 267875 37213
rect 247141 18003 247175 27557
rect 249993 18003 250027 27557
rect 251373 19295 251407 27557
rect 265173 18003 265207 27557
rect 272257 26299 272291 35853
rect 284769 29019 284803 44693
rect 270509 17935 270543 22117
rect 284769 18003 284803 27557
rect 285965 18003 285999 27557
rect 294245 26299 294279 45509
rect 301145 26299 301179 35853
rect 303813 32419 303847 38573
rect 323317 37315 323351 46869
rect 327273 37315 327307 46869
rect 330125 37315 330159 46869
rect 336933 37315 336967 46869
rect 337209 37383 337243 46869
rect 341257 37315 341291 46869
rect 357633 37315 357667 46801
rect 358645 37315 358679 46869
rect 359013 37315 359047 46869
rect 367017 37315 367051 46869
rect 421205 37315 421239 46869
rect 460029 41395 460063 48161
rect 310897 26299 310931 35853
rect 341257 29087 341291 32249
rect 236285 8347 236319 17901
rect 244381 8347 244415 17901
rect 273453 10931 273487 17901
rect 310897 15215 310931 22117
rect 337117 18003 337151 18445
rect 295625 12223 295659 12461
rect 341257 9707 341291 27557
rect 357633 18003 357667 27557
rect 358553 9707 358587 27557
rect 366833 9707 366867 27557
rect 386245 16643 386279 26197
rect 421205 9707 421239 27557
rect 470609 9707 470643 19261
rect 227545 6987 227579 7633
rect 268393 5015 268427 5253
rect 224233 4811 224267 4913
rect 224141 4267 224175 4777
rect 249073 4267 249107 4981
rect 278053 5015 278087 5253
rect 287713 5015 287747 5457
rect 297097 5015 297131 5457
rect 257997 4267 258031 4981
rect 307033 4199 307067 4981
rect 317337 4743 317371 4845
rect 319453 4471 319487 4641
rect 322673 4607 322707 5049
rect 322765 4879 322799 5049
rect 325157 4811 325191 4981
rect 326169 4675 326203 4913
rect 327181 4811 327215 5049
rect 326629 4675 326663 4777
rect 326261 4641 326663 4675
rect 326261 4607 326295 4641
rect 337117 4471 337151 6069
rect 461225 4879 461259 5117
rect 466101 4947 466135 5253
rect 471345 4811 471379 5049
rect 471437 4811 471471 5525
rect 283113 4165 283331 4199
rect 355241 4165 355459 4199
rect 283113 4131 283147 4165
rect 269129 3927 269163 4097
rect 283205 3995 283239 4097
rect 283297 3995 283331 4165
rect 355241 4131 355275 4165
rect 332333 3927 332367 4097
rect 45477 3179 45511 3349
rect 82921 2975 82955 3145
rect 276305 3043 276339 3213
rect 282837 3043 282871 3349
rect 285873 3315 285907 3757
rect 292497 3315 292531 3689
rect 320833 3587 320867 3893
rect 320741 3519 320775 3553
rect 320925 3519 320959 3893
rect 326353 3723 326387 3893
rect 332241 3791 332275 3893
rect 332149 3587 332183 3757
rect 320741 3485 320959 3519
rect 335369 3587 335403 4097
rect 340797 4097 340889 4131
rect 335921 3723 335955 3893
rect 322765 3111 322799 3553
rect 335737 3043 335771 3553
rect 340647 3145 340739 3179
rect 335829 2975 335863 3145
rect 93869 2839 93903 2941
rect 335645 2839 335679 2941
rect 340705 2907 340739 3145
rect 340797 2839 340831 4097
rect 343925 2839 343959 3213
rect 344109 2907 344143 3213
rect 344385 2975 344419 3349
rect 345489 595 345523 3281
rect 345673 3179 345707 3349
rect 349169 3315 349203 4097
rect 347789 2771 347823 2941
rect 350089 2771 350123 2941
rect 352665 2907 352699 4097
rect 352849 2839 352883 3621
rect 352941 3383 352975 3621
rect 355333 3247 355367 4097
rect 355425 3655 355459 4165
rect 376769 3927 376803 4777
rect 361957 3451 361991 3689
rect 355425 3111 355459 3213
rect 362049 3179 362083 3689
rect 376861 3519 376895 4369
rect 376803 3485 376895 3519
rect 410993 3451 411027 3893
rect 417525 3723 417559 3961
rect 354873 3077 355459 3111
rect 354873 2907 354907 3077
rect 365729 2907 365763 3145
rect 375297 2907 375331 3077
rect 413201 2907 413235 3485
rect 418169 2839 418203 4097
rect 420101 3519 420135 3961
rect 422125 2839 422159 3689
rect 422953 3111 422987 3621
rect 423045 3519 423079 3689
rect 423137 3247 423171 3689
rect 426449 3179 426483 3689
rect 427737 3111 427771 4097
rect 437489 3995 437523 4233
rect 438259 4165 438409 4199
rect 430037 3451 430071 3689
rect 423045 2907 423079 3077
rect 430129 2771 430163 3689
rect 434579 3553 434637 3587
rect 432521 3111 432555 3417
rect 432613 2907 432647 3417
rect 435925 3247 435959 3961
rect 445861 3791 445895 4097
rect 441721 2839 441755 3689
rect 446781 3247 446815 4029
rect 451933 3859 451967 4097
rect 456809 3723 456843 3961
rect 449909 2975 449943 3621
rect 450277 2907 450311 3009
rect 451231 2805 451473 2839
rect 444849 595 444883 2805
rect 454693 2159 454727 3553
rect 456901 2907 456935 3689
rect 466377 2907 466411 3757
rect 456843 2873 456935 2907
rect 466193 2771 466227 2873
rect 466929 2839 466963 3757
rect 471529 595 471563 5593
rect 518173 3043 518207 3213
<< viali >>
rect 364533 685797 364567 685831
rect 364533 676209 364567 676243
rect 429577 684437 429611 684471
rect 559297 684437 559331 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 364533 618205 364567 618239
rect 364533 608617 364567 608651
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 364625 598893 364659 598927
rect 364625 589305 364659 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 247969 579309 248003 579343
rect 254225 579309 254259 579343
rect 292129 579309 292163 579343
rect 292129 579105 292163 579139
rect 415685 579309 415719 579343
rect 254225 578629 254259 578663
rect 247969 578561 248003 578595
rect 415685 578493 415719 578527
rect 428381 579309 428415 579343
rect 428381 578425 428415 578459
rect 441077 579309 441111 579343
rect 441077 578357 441111 578391
rect 453589 579309 453623 579343
rect 453589 578289 453623 578323
rect 455797 579309 455831 579343
rect 455797 578221 455831 578255
rect 346409 338657 346443 338691
rect 327089 338113 327123 338147
rect 315497 338045 315531 338079
rect 318901 338045 318935 338079
rect 319085 338045 319119 338079
rect 96077 337977 96111 338011
rect 96261 337977 96295 338011
rect 115397 337977 115431 338011
rect 115581 337977 115615 338011
rect 134717 337977 134751 338011
rect 134901 337977 134935 338011
rect 154037 337977 154071 338011
rect 154221 337977 154255 338011
rect 173357 337977 173391 338011
rect 173541 337977 173575 338011
rect 192677 337977 192711 338011
rect 192861 337977 192895 338011
rect 211997 337977 212031 338011
rect 212181 337977 212215 338011
rect 96261 337841 96295 337875
rect 96445 337841 96479 337875
rect 115581 337841 115615 337875
rect 115765 337841 115799 337875
rect 134901 337841 134935 337875
rect 135085 337841 135119 337875
rect 154221 337841 154255 337875
rect 154405 337841 154439 337875
rect 173541 337841 173575 337875
rect 173725 337841 173759 337875
rect 192861 337841 192895 337875
rect 193045 337841 193079 337875
rect 212181 337841 212215 337875
rect 212365 337841 212399 337875
rect 302157 337773 302191 337807
rect 96353 337569 96387 337603
rect 96537 337569 96571 337603
rect 115673 337569 115707 337603
rect 115857 337569 115891 337603
rect 134993 337569 135027 337603
rect 135177 337569 135211 337603
rect 154313 337569 154347 337603
rect 154497 337569 154531 337603
rect 173633 337569 173667 337603
rect 173817 337569 173851 337603
rect 192953 337569 192987 337603
rect 193137 337569 193171 337603
rect 212273 337569 212307 337603
rect 212457 337569 212491 337603
rect 241529 337705 241563 337739
rect 302249 337705 302283 337739
rect 303997 337773 304031 337807
rect 96261 337501 96295 337535
rect 96445 337501 96479 337535
rect 115581 337501 115615 337535
rect 115765 337501 115799 337535
rect 134901 337501 134935 337535
rect 135085 337501 135119 337535
rect 154221 337501 154255 337535
rect 154405 337501 154439 337535
rect 173541 337501 173575 337535
rect 173725 337501 173759 337535
rect 192861 337501 192895 337535
rect 193045 337501 193079 337535
rect 212181 337501 212215 337535
rect 212365 337501 212399 337535
rect 230489 337501 230523 337535
rect 230581 337637 230615 337671
rect 231225 337637 231259 337671
rect 234445 337637 234479 337671
rect 230581 337501 230615 337535
rect 241529 337501 241563 337535
rect 259745 337637 259779 337671
rect 96169 337433 96203 337467
rect 96353 337433 96387 337467
rect 115489 337433 115523 337467
rect 115673 337433 115707 337467
rect 134809 337433 134843 337467
rect 134993 337433 135027 337467
rect 154129 337433 154163 337467
rect 154313 337433 154347 337467
rect 173449 337433 173483 337467
rect 173633 337433 173667 337467
rect 192769 337433 192803 337467
rect 192953 337433 192987 337467
rect 212089 337433 212123 337467
rect 212273 337433 212307 337467
rect 234445 337433 234479 337467
rect 115397 337365 115431 337399
rect 115857 337365 115891 337399
rect 134717 337365 134751 337399
rect 135177 337365 135211 337399
rect 154037 337365 154071 337399
rect 154497 337365 154531 337399
rect 173357 337365 173391 337399
rect 173817 337365 173851 337399
rect 192677 337365 192711 337399
rect 193137 337365 193171 337399
rect 211997 337365 212031 337399
rect 212457 337365 212491 337399
rect 259745 337365 259779 337399
rect 318901 337909 318935 337943
rect 318993 337909 319027 337943
rect 318809 337773 318843 337807
rect 318993 337773 319027 337807
rect 336657 338113 336691 338147
rect 327089 337705 327123 337739
rect 335921 337841 335955 337875
rect 318901 337569 318935 337603
rect 318993 337569 319027 337603
rect 335829 337501 335863 337535
rect 318809 337433 318843 337467
rect 319085 337433 319119 337467
rect 334725 337365 334759 337399
rect 315497 337297 315531 337331
rect 326353 337297 326387 337331
rect 115581 337161 115615 337195
rect 115857 337161 115891 337195
rect 303997 337161 304031 337195
rect 326353 337161 326387 337195
rect 115489 337093 115523 337127
rect 115765 337093 115799 337127
rect 134809 337093 134843 337127
rect 135085 337093 135119 337127
rect 154129 337093 154163 337127
rect 154313 337093 154347 337127
rect 173449 337093 173483 337127
rect 173633 337093 173667 337127
rect 192769 337093 192803 337127
rect 192953 337093 192987 337127
rect 212089 337093 212123 337127
rect 212273 337093 212307 337127
rect 134717 337025 134751 337059
rect 134993 337025 135027 337059
rect 154037 337025 154071 337059
rect 154405 337025 154439 337059
rect 173357 337025 173391 337059
rect 173725 337025 173759 337059
rect 192677 337025 192711 337059
rect 193045 337025 193079 337059
rect 211997 337025 212031 337059
rect 212365 337025 212399 337059
rect 336013 337841 336047 337875
rect 336657 337705 336691 337739
rect 442365 338113 442399 338147
rect 372721 338045 372755 338079
rect 412465 338045 412499 338079
rect 372721 337773 372755 337807
rect 374653 337909 374687 337943
rect 346409 337705 346443 337739
rect 336013 337637 336047 337671
rect 344661 337637 344695 337671
rect 364993 337637 365027 337671
rect 341717 337501 341751 337535
rect 335921 337365 335955 337399
rect 336197 337365 336231 337399
rect 335829 337025 335863 337059
rect 340797 337365 340831 337399
rect 340797 337093 340831 337127
rect 340889 337365 340923 337399
rect 336197 336889 336231 336923
rect 340613 337025 340647 337059
rect 334725 336753 334759 336787
rect 341717 337229 341751 337263
rect 342821 337501 342855 337535
rect 344293 337501 344327 337535
rect 342821 337161 342855 337195
rect 345581 337365 345615 337399
rect 354045 337365 354079 337399
rect 345857 337161 345891 337195
rect 345857 336957 345891 336991
rect 365361 337569 365395 337603
rect 365085 337501 365119 337535
rect 365269 337501 365303 337535
rect 365361 337433 365395 337467
rect 374561 337433 374595 337467
rect 364993 337161 365027 337195
rect 369869 337365 369903 337399
rect 369869 337161 369903 337195
rect 374561 337161 374595 337195
rect 354045 336957 354079 336991
rect 432521 338045 432555 338079
rect 430037 337977 430071 338011
rect 412465 337705 412499 337739
rect 414121 337705 414155 337739
rect 430037 337705 430071 337739
rect 442273 338045 442307 338079
rect 434085 337977 434119 338011
rect 432521 337501 432555 337535
rect 432613 337773 432647 337807
rect 414121 337365 414155 337399
rect 432613 337365 432647 337399
rect 432705 337637 432739 337671
rect 374653 336957 374687 336991
rect 423045 337229 423079 337263
rect 431417 337161 431451 337195
rect 423045 336957 423079 336991
rect 429301 337093 429335 337127
rect 345581 336889 345615 336923
rect 340889 336821 340923 336855
rect 345489 336821 345523 336855
rect 345765 336821 345799 336855
rect 431417 337025 431451 337059
rect 434545 337909 434579 337943
rect 442273 337909 442307 337943
rect 483121 338045 483155 338079
rect 442365 337909 442399 337943
rect 444389 337977 444423 338011
rect 434269 337841 434303 337875
rect 434453 337841 434487 337875
rect 434545 337705 434579 337739
rect 437305 337637 437339 337671
rect 434085 337093 434119 337127
rect 436109 337433 436143 337467
rect 432705 336957 432739 336991
rect 432429 336889 432463 336923
rect 432613 336821 432647 336855
rect 436109 336821 436143 336855
rect 340797 336753 340831 336787
rect 340981 336753 341015 336787
rect 341165 336753 341199 336787
rect 429301 336753 429335 336787
rect 452025 337977 452059 338011
rect 449449 337841 449483 337875
rect 449449 337637 449483 337671
rect 451933 337773 451967 337807
rect 452025 337773 452059 337807
rect 455889 337977 455923 338011
rect 483213 337977 483247 338011
rect 461501 337909 461535 337943
rect 455889 337773 455923 337807
rect 456717 337841 456751 337875
rect 444389 337569 444423 337603
rect 437673 337501 437707 337535
rect 451933 337433 451967 337467
rect 445769 337365 445803 337399
rect 437489 337161 437523 337195
rect 437581 337161 437615 337195
rect 437489 336821 437523 336855
rect 445769 336821 445803 336855
rect 450369 337365 450403 337399
rect 450369 336821 450403 336855
rect 466377 337909 466411 337943
rect 461409 337637 461443 337671
rect 461501 337637 461535 337671
rect 463709 337841 463743 337875
rect 437397 336753 437431 336787
rect 456717 336753 456751 336787
rect 459017 337297 459051 337331
rect 461409 337297 461443 337331
rect 463709 337297 463743 337331
rect 466193 337297 466227 337331
rect 466377 337297 466411 337331
rect 469229 337909 469263 337943
rect 483121 337909 483155 337943
rect 483305 337909 483339 337943
rect 483121 337773 483155 337807
rect 483305 337773 483339 337807
rect 483121 337637 483155 337671
rect 483305 337637 483339 337671
rect 483029 337433 483063 337467
rect 483213 337433 483247 337467
rect 466285 337229 466319 337263
rect 469229 337229 469263 337263
rect 466193 336821 466227 336855
rect 466285 336889 466319 336923
rect 466377 336889 466411 336923
rect 284401 336685 284435 336719
rect 284401 335189 284435 335223
rect 288817 336685 288851 336719
rect 250177 334441 250211 334475
rect 250177 328457 250211 328491
rect 259837 328389 259871 328423
rect 259837 318801 259871 318835
rect 262689 322269 262723 322303
rect 266645 321589 266679 321623
rect 262689 317441 262723 317475
rect 265265 318869 265299 318903
rect 266645 318801 266679 318835
rect 267749 321589 267783 321623
rect 327273 336685 327307 336719
rect 302525 334713 302559 334747
rect 302525 328457 302559 328491
rect 327273 327097 327307 327131
rect 339785 336685 339819 336719
rect 288817 319073 288851 319107
rect 299857 327029 299891 327063
rect 267749 318801 267783 318835
rect 265265 317441 265299 317475
rect 421205 336685 421239 336719
rect 459017 336685 459051 336719
rect 339785 318801 339819 318835
rect 341349 328389 341383 328423
rect 341349 318801 341383 318835
rect 358737 328389 358771 328423
rect 469597 336753 469631 336787
rect 469413 336685 469447 336719
rect 466285 336617 466319 336651
rect 421205 327097 421239 327131
rect 470609 328389 470643 328423
rect 358737 318801 358771 318835
rect 359197 327029 359231 327063
rect 470609 318801 470643 318835
rect 359197 317713 359231 317747
rect 372721 318733 372755 318767
rect 299857 317441 299891 317475
rect 358737 317373 358771 317407
rect 262689 315945 262723 315979
rect 244473 311797 244507 311831
rect 244473 309145 244507 309179
rect 236285 309077 236319 309111
rect 259653 309077 259687 309111
rect 272165 314585 272199 314619
rect 262689 306357 262723 306391
rect 265265 309077 265299 309111
rect 259653 299557 259687 299591
rect 236285 299489 236319 299523
rect 265265 299489 265299 299523
rect 266645 298129 266679 298163
rect 266645 296701 266679 296735
rect 288725 311933 288759 311967
rect 284585 311865 284619 311899
rect 273453 309281 273487 309315
rect 285965 311865 285999 311899
rect 285965 306425 285999 306459
rect 284585 306357 284619 306391
rect 273453 301529 273487 301563
rect 272165 296701 272199 296735
rect 272165 295273 272199 295307
rect 251465 294661 251499 294695
rect 251465 289833 251499 289867
rect 310897 311933 310931 311967
rect 310897 307853 310931 307887
rect 339877 309077 339911 309111
rect 310713 307717 310747 307751
rect 337025 307717 337059 307751
rect 327273 302141 327307 302175
rect 310713 298129 310747 298163
rect 323317 299421 323351 299455
rect 288725 289969 288759 290003
rect 310897 293029 310931 293063
rect 295533 288473 295567 288507
rect 295533 287045 295567 287079
rect 272165 285685 272199 285719
rect 296821 286977 296855 287011
rect 266737 285617 266771 285651
rect 236285 280109 236319 280143
rect 236285 270521 236319 270555
rect 239137 280109 239171 280143
rect 239137 270521 239171 270555
rect 251465 280109 251499 280143
rect 259561 280109 259595 280143
rect 266737 276029 266771 276063
rect 324697 299421 324731 299455
rect 339877 299897 339911 299931
rect 341165 309077 341199 309111
rect 421205 317373 421239 317407
rect 372721 309145 372755 309179
rect 386797 315945 386831 315979
rect 358737 307785 358771 307819
rect 421205 307785 421239 307819
rect 460213 317373 460247 317407
rect 460213 307785 460247 307819
rect 470609 309077 470643 309111
rect 386797 302073 386831 302107
rect 341165 299489 341199 299523
rect 470609 299489 470643 299523
rect 337025 298197 337059 298231
rect 372721 299421 372755 299455
rect 327273 298129 327307 298163
rect 337209 298061 337243 298095
rect 337209 292417 337243 292451
rect 358737 298061 358771 298095
rect 324697 289833 324731 289867
rect 323317 288473 323351 288507
rect 341165 289765 341199 289799
rect 310897 282761 310931 282795
rect 337117 282897 337151 282931
rect 325893 280177 325927 280211
rect 325893 278749 325927 278783
rect 336933 280109 336967 280143
rect 296821 276029 296855 276063
rect 310897 278681 310931 278715
rect 259561 273037 259595 273071
rect 266645 274601 266679 274635
rect 251465 270521 251499 270555
rect 250085 269025 250119 269059
rect 236285 260797 236319 260831
rect 236285 251209 236319 251243
rect 239137 260797 239171 260831
rect 310897 263449 310931 263483
rect 330125 273921 330159 273955
rect 359105 298061 359139 298095
rect 372721 289833 372755 289867
rect 375665 299421 375699 299455
rect 421205 298061 421239 298095
rect 375665 289833 375699 289867
rect 386797 293029 386831 293063
rect 359105 288405 359139 288439
rect 421205 288405 421239 288439
rect 460029 298061 460063 298095
rect 460029 288405 460063 288439
rect 470609 289765 470643 289799
rect 386797 282761 386831 282795
rect 358737 280245 358771 280279
rect 341165 280177 341199 280211
rect 470609 280177 470643 280211
rect 337117 278749 337151 278783
rect 372721 280109 372755 280143
rect 336933 270521 336967 270555
rect 372721 270521 372755 270555
rect 377137 280109 377171 280143
rect 460121 280109 460155 280143
rect 377137 270521 377171 270555
rect 386797 278681 386831 278715
rect 330125 260865 330159 260899
rect 341165 270453 341199 270487
rect 460121 273105 460155 273139
rect 463801 275281 463835 275315
rect 463801 270521 463835 270555
rect 386797 263449 386831 263483
rect 460029 270453 460063 270487
rect 460029 260933 460063 260967
rect 470609 270453 470643 270487
rect 341165 260865 341199 260899
rect 470609 260865 470643 260899
rect 250085 259437 250119 259471
rect 251465 260797 251499 260831
rect 239137 251209 239171 251243
rect 250177 259301 250211 259335
rect 259561 260797 259595 260831
rect 266645 260797 266679 260831
rect 270693 260797 270727 260831
rect 259561 253725 259595 253759
rect 265357 255901 265391 255935
rect 251465 251209 251499 251243
rect 250177 251073 250211 251107
rect 259561 251141 259595 251175
rect 265357 248217 265391 248251
rect 259561 244137 259595 244171
rect 336933 260797 336967 260831
rect 272533 258009 272567 258043
rect 310897 256037 310931 256071
rect 310897 251277 310931 251311
rect 327181 253929 327215 253963
rect 310713 251141 310747 251175
rect 272533 249713 272567 249747
rect 284677 249713 284711 249747
rect 270693 240193 270727 240227
rect 288909 245565 288943 245599
rect 284677 240125 284711 240159
rect 285965 244953 285999 244987
rect 270693 238697 270727 238731
rect 262597 235909 262631 235943
rect 310713 241485 310747 241519
rect 288909 235977 288943 236011
rect 299489 241417 299523 241451
rect 285965 234481 285999 234515
rect 270693 233801 270727 233835
rect 372721 260797 372755 260831
rect 358737 259369 358771 259403
rect 336933 249781 336967 249815
rect 337117 254609 337151 254643
rect 337117 241553 337151 241587
rect 327181 240193 327215 240227
rect 372721 251209 372755 251243
rect 377137 260797 377171 260831
rect 377137 251209 377171 251243
rect 463709 260797 463743 260831
rect 463709 251209 463743 251243
rect 367017 251141 367051 251175
rect 367017 241485 367051 241519
rect 470609 251141 470643 251175
rect 470609 241485 470643 241519
rect 358737 240125 358771 240159
rect 324605 240057 324639 240091
rect 299489 231829 299523 231863
rect 323409 234685 323443 234719
rect 310805 231761 310839 231795
rect 323409 231761 323443 231795
rect 324605 231761 324639 231795
rect 327181 240057 327215 240091
rect 262597 226321 262631 226355
rect 272073 229041 272107 229075
rect 327181 230537 327215 230571
rect 337117 234617 337151 234651
rect 337117 230469 337151 230503
rect 310805 222173 310839 222207
rect 358737 230401 358771 230435
rect 272073 220745 272107 220779
rect 299489 222105 299523 222139
rect 290105 217957 290139 217991
rect 290105 208369 290139 208403
rect 291669 214557 291703 214591
rect 358737 220813 358771 220847
rect 341165 220745 341199 220779
rect 341165 215237 341199 215271
rect 299489 212517 299523 212551
rect 291669 204017 291703 204051
rect 310805 212449 310839 212483
rect 310805 202861 310839 202895
rect 299489 202793 299523 202827
rect 272349 201433 272383 201467
rect 250085 200073 250119 200107
rect 265173 200073 265207 200107
rect 265173 195245 265207 195279
rect 299489 193205 299523 193239
rect 336933 202793 336967 202827
rect 336933 193205 336967 193239
rect 272349 193137 272383 193171
rect 367017 193137 367051 193171
rect 250085 186269 250119 186303
rect 266645 191777 266679 191811
rect 266645 186269 266679 186303
rect 288817 191777 288851 191811
rect 284677 180761 284711 180795
rect 259653 179537 259687 179571
rect 259653 173961 259687 173995
rect 288817 179401 288851 179435
rect 290013 188649 290047 188683
rect 299857 188445 299891 188479
rect 290013 179401 290047 179435
rect 294337 184229 294371 184263
rect 299857 183549 299891 183583
rect 306849 188445 306883 188479
rect 306849 183549 306883 183583
rect 367017 183549 367051 183583
rect 337117 183481 337151 183515
rect 294337 179401 294371 179435
rect 299857 180761 299891 180795
rect 294429 177973 294463 178007
rect 284677 171105 284711 171139
rect 288817 176613 288851 176647
rect 285965 171037 285999 171071
rect 299857 171105 299891 171139
rect 301053 180761 301087 180795
rect 301053 171105 301087 171139
rect 302617 180761 302651 180795
rect 460121 183481 460155 183515
rect 460121 176477 460155 176511
rect 337117 172533 337151 172567
rect 302617 171105 302651 171139
rect 330125 172465 330159 172499
rect 294429 168385 294463 168419
rect 288817 167025 288851 167059
rect 460121 166957 460155 166991
rect 330125 162945 330159 162979
rect 372813 164169 372847 164203
rect 285965 161449 285999 161483
rect 330125 161381 330159 161415
rect 286057 158661 286091 158695
rect 272165 157981 272199 158015
rect 259653 154173 259687 154207
rect 232329 143497 232363 143531
rect 272165 148937 272199 148971
rect 259653 142137 259687 142171
rect 270693 144857 270727 144891
rect 232329 133909 232363 133943
rect 259837 142001 259871 142035
rect 239137 125545 239171 125579
rect 232329 124117 232363 124151
rect 251465 125545 251499 125579
rect 239137 115957 239171 115991
rect 249993 124117 250027 124151
rect 232329 114529 232363 114563
rect 270693 139961 270727 139995
rect 272441 143497 272475 143531
rect 294337 158661 294371 158695
rect 294337 149073 294371 149107
rect 310805 153153 310839 153187
rect 372813 157301 372847 157335
rect 421205 162809 421239 162843
rect 460121 161449 460155 161483
rect 421205 153221 421239 153255
rect 330125 151793 330159 151827
rect 341165 153153 341199 153187
rect 310805 147577 310839 147611
rect 460121 151725 460155 151759
rect 341165 144857 341199 144891
rect 360209 147713 360243 147747
rect 360209 144857 360243 144891
rect 367017 144857 367051 144891
rect 286057 140777 286091 140811
rect 323317 143497 323351 143531
rect 272441 135201 272475 135235
rect 288633 140709 288667 140743
rect 259837 124185 259871 124219
rect 265265 133841 265299 133875
rect 295533 140709 295567 140743
rect 294429 139349 294463 139383
rect 289921 138057 289955 138091
rect 289921 132413 289955 132447
rect 288633 131121 288667 131155
rect 291485 131053 291519 131087
rect 265265 124185 265299 124219
rect 270693 125545 270727 125579
rect 270693 120649 270727 120683
rect 272441 124117 272475 124151
rect 251465 115957 251499 115991
rect 249993 114529 250027 114563
rect 323317 133909 323351 133943
rect 324605 143497 324639 143531
rect 330125 143497 330159 143531
rect 330125 137921 330159 137955
rect 421205 143497 421239 143531
rect 377137 140029 377171 140063
rect 367017 135269 367051 135303
rect 372721 138125 372755 138159
rect 372721 135269 372755 135303
rect 377137 135269 377171 135303
rect 324605 132481 324639 132515
rect 358737 135201 358771 135235
rect 295533 131121 295567 131155
rect 337209 132413 337243 132447
rect 294429 129761 294463 129795
rect 296913 131053 296947 131087
rect 291485 122689 291519 122723
rect 296913 121465 296947 121499
rect 299857 124117 299891 124151
rect 272441 114529 272475 114563
rect 299857 114529 299891 114563
rect 306849 124117 306883 124151
rect 306849 113237 306883 113271
rect 324697 122757 324731 122791
rect 463709 147713 463743 147747
rect 463709 144925 463743 144959
rect 460121 142205 460155 142239
rect 421205 133909 421239 133943
rect 460121 142069 460155 142103
rect 460121 132481 460155 132515
rect 358737 125613 358771 125647
rect 339785 125545 339819 125579
rect 339785 118609 339819 118643
rect 341165 125545 341199 125579
rect 341165 118609 341199 118643
rect 421205 124117 421239 124151
rect 337209 114529 337243 114563
rect 341165 115889 341199 115923
rect 324697 113169 324731 113203
rect 327181 114461 327215 114495
rect 265265 113101 265299 113135
rect 247233 109021 247267 109055
rect 247233 106301 247267 106335
rect 251465 106233 251499 106267
rect 232329 104805 232363 104839
rect 284677 113101 284711 113135
rect 265265 103513 265299 103547
rect 270693 106233 270727 106267
rect 266829 103445 266863 103479
rect 251465 96645 251499 96679
rect 262781 102085 262815 102119
rect 232329 95217 232363 95251
rect 247141 95149 247175 95183
rect 236285 86921 236319 86955
rect 232329 85493 232363 85527
rect 266829 96441 266863 96475
rect 267933 103445 267967 103479
rect 291577 113101 291611 113135
rect 296821 113101 296855 113135
rect 291577 103581 291611 103615
rect 294337 109701 294371 109735
rect 284677 103513 284711 103547
rect 325985 106301 326019 106335
rect 325985 104873 326019 104907
rect 341165 106301 341199 106335
rect 367017 115889 367051 115923
rect 421205 114529 421239 114563
rect 470609 115889 470643 115923
rect 367017 106301 367051 106335
rect 470609 106301 470643 106335
rect 327181 104873 327215 104907
rect 386521 106233 386555 106267
rect 341165 104805 341199 104839
rect 296821 103513 296855 103547
rect 339785 104737 339819 104771
rect 294337 102153 294371 102187
rect 295625 103445 295659 103479
rect 270693 101337 270727 101371
rect 291669 102085 291703 102119
rect 267933 93857 267967 93891
rect 262781 92497 262815 92531
rect 295625 93857 295659 93891
rect 301145 103445 301179 103479
rect 301145 93857 301179 93891
rect 306849 103445 306883 103479
rect 324605 103445 324639 103479
rect 306849 93857 306883 93891
rect 310805 95149 310839 95183
rect 291669 92497 291703 92531
rect 262689 88961 262723 88995
rect 247141 85561 247175 85595
rect 251465 86921 251499 86955
rect 236285 77401 236319 77435
rect 251465 77265 251499 77299
rect 232329 75905 232363 75939
rect 265173 88961 265207 88995
rect 324605 93857 324639 93891
rect 330125 102085 330159 102119
rect 265173 84269 265207 84303
rect 291577 85561 291611 85595
rect 310805 85561 310839 85595
rect 317705 88349 317739 88383
rect 291577 84201 291611 84235
rect 299857 85493 299891 85527
rect 262689 75905 262723 75939
rect 265357 84133 265391 84167
rect 272257 84133 272291 84167
rect 265357 74545 265391 74579
rect 270785 80733 270819 80767
rect 239137 70465 239171 70499
rect 239137 67609 239171 67643
rect 244473 70465 244507 70499
rect 244473 67609 244507 67643
rect 272257 74545 272291 74579
rect 284677 84133 284711 84167
rect 270785 67609 270819 67643
rect 272257 67677 272291 67711
rect 250085 67541 250119 67575
rect 232329 66181 232363 66215
rect 232329 56593 232363 56627
rect 236285 66181 236319 66215
rect 236285 56593 236319 56627
rect 239045 58021 239079 58055
rect 272257 67065 272291 67099
rect 284677 66249 284711 66283
rect 285965 84133 285999 84167
rect 285965 66249 285999 66283
rect 288725 82773 288759 82807
rect 270785 66181 270819 66215
rect 250085 57953 250119 57987
rect 265173 62645 265207 62679
rect 265173 57885 265207 57919
rect 239045 56593 239079 56627
rect 270785 56593 270819 56627
rect 273453 66181 273487 66215
rect 244565 56525 244599 56559
rect 239137 53193 239171 53227
rect 239137 48297 239171 48331
rect 236285 48229 236319 48263
rect 299857 75905 299891 75939
rect 324697 85493 324731 85527
rect 339785 95217 339819 95251
rect 386521 99297 386555 99331
rect 421205 104805 421239 104839
rect 341165 95217 341199 95251
rect 360301 96577 360335 96611
rect 341073 90389 341107 90423
rect 330125 77265 330159 77299
rect 336933 86921 336967 86955
rect 324697 75973 324731 76007
rect 317705 75905 317739 75939
rect 337209 86921 337243 86955
rect 337209 77265 337243 77299
rect 360301 89641 360335 89675
rect 367017 96577 367051 96611
rect 367017 86989 367051 87023
rect 421205 86989 421239 87023
rect 470609 96577 470643 96611
rect 470609 86989 470643 87023
rect 341073 77265 341107 77299
rect 358737 85493 358771 85527
rect 336933 75905 336967 75939
rect 421205 85493 421239 85527
rect 358737 75905 358771 75939
rect 386613 77197 386647 77231
rect 310805 75837 310839 75871
rect 310805 66317 310839 66351
rect 324605 75837 324639 75871
rect 377137 70465 377171 70499
rect 377137 67609 377171 67643
rect 421205 75905 421239 75939
rect 470609 77197 470643 77231
rect 386613 67609 386647 67643
rect 470609 67609 470643 67643
rect 324605 66317 324639 66351
rect 375665 67541 375699 67575
rect 288725 64889 288759 64923
rect 310805 66181 310839 66215
rect 273453 50949 273487 50983
rect 294245 64821 294279 64855
rect 244565 48161 244599 48195
rect 273545 48229 273579 48263
rect 244565 46869 244599 46903
rect 236285 38641 236319 38675
rect 239045 42041 239079 42075
rect 236285 38505 236319 38539
rect 236285 31637 236319 31671
rect 244565 37281 244599 37315
rect 262781 45509 262815 45543
rect 239045 28985 239079 29019
rect 259745 37213 259779 37247
rect 236377 28917 236411 28951
rect 310805 59993 310839 60027
rect 323317 66181 323351 66215
rect 294245 46937 294279 46971
rect 299673 56525 299707 56559
rect 301053 56525 301087 56559
rect 324605 66181 324639 66215
rect 324605 61353 324639 61387
rect 330125 66181 330159 66215
rect 330125 56593 330159 56627
rect 336933 66181 336967 66215
rect 358645 66181 358679 66215
rect 336933 56593 336967 56627
rect 339785 57885 339819 57919
rect 323317 48297 323351 48331
rect 324789 56525 324823 56559
rect 301053 46937 301087 46971
rect 337301 56525 337335 56559
rect 358645 56593 358679 56627
rect 367017 66181 367051 66215
rect 339785 48297 339819 48331
rect 357541 56457 357575 56491
rect 337301 47005 337335 47039
rect 324789 46937 324823 46971
rect 375665 61965 375699 61999
rect 421205 66181 421239 66215
rect 421205 56593 421239 56627
rect 460029 57885 460063 57919
rect 367017 48297 367051 48331
rect 460029 48297 460063 48331
rect 470609 57885 470643 57919
rect 470609 48297 470643 48331
rect 357541 46937 357575 46971
rect 460029 48161 460063 48195
rect 299673 45577 299707 45611
rect 323317 46869 323351 46903
rect 294245 45509 294279 45543
rect 273545 38641 273579 38675
rect 284769 44693 284803 44727
rect 262781 35921 262815 35955
rect 267841 37213 267875 37247
rect 267841 28577 267875 28611
rect 272257 35853 272291 35887
rect 259745 27625 259779 27659
rect 236377 22729 236411 22763
rect 247141 27557 247175 27591
rect 247141 17969 247175 18003
rect 249993 27557 250027 27591
rect 251373 27557 251407 27591
rect 251373 19261 251407 19295
rect 265173 27557 265207 27591
rect 249993 17969 250027 18003
rect 284769 28985 284803 29019
rect 272257 26265 272291 26299
rect 284769 27557 284803 27591
rect 265173 17969 265207 18003
rect 270509 22117 270543 22151
rect 284769 17969 284803 18003
rect 285965 27557 285999 27591
rect 303813 38573 303847 38607
rect 294245 26265 294279 26299
rect 301145 35853 301179 35887
rect 323317 37281 323351 37315
rect 327273 46869 327307 46903
rect 327273 37281 327307 37315
rect 330125 46869 330159 46903
rect 330125 37281 330159 37315
rect 336933 46869 336967 46903
rect 337209 46869 337243 46903
rect 337209 37349 337243 37383
rect 341257 46869 341291 46903
rect 336933 37281 336967 37315
rect 358645 46869 358679 46903
rect 341257 37281 341291 37315
rect 357633 46801 357667 46835
rect 357633 37281 357667 37315
rect 358645 37281 358679 37315
rect 359013 46869 359047 46903
rect 359013 37281 359047 37315
rect 367017 46869 367051 46903
rect 367017 37281 367051 37315
rect 421205 46869 421239 46903
rect 460029 41361 460063 41395
rect 421205 37281 421239 37315
rect 303813 32385 303847 32419
rect 310897 35853 310931 35887
rect 301145 26265 301179 26299
rect 341257 32249 341291 32283
rect 341257 29053 341291 29087
rect 310897 26265 310931 26299
rect 341257 27557 341291 27591
rect 285965 17969 285999 18003
rect 310897 22117 310931 22151
rect 236285 17901 236319 17935
rect 236285 8313 236319 8347
rect 244381 17901 244415 17935
rect 270509 17901 270543 17935
rect 273453 17901 273487 17935
rect 337117 18445 337151 18479
rect 337117 17969 337151 18003
rect 310897 15181 310931 15215
rect 295625 12461 295659 12495
rect 295625 12189 295659 12223
rect 273453 10897 273487 10931
rect 357633 27557 357667 27591
rect 357633 17969 357667 18003
rect 358553 27557 358587 27591
rect 341257 9673 341291 9707
rect 358553 9673 358587 9707
rect 366833 27557 366867 27591
rect 421205 27557 421239 27591
rect 386245 26197 386279 26231
rect 386245 16609 386279 16643
rect 366833 9673 366867 9707
rect 421205 9673 421239 9707
rect 470609 19261 470643 19295
rect 470609 9673 470643 9707
rect 244381 8313 244415 8347
rect 227545 7633 227579 7667
rect 227545 6953 227579 6987
rect 337117 6069 337151 6103
rect 287713 5457 287747 5491
rect 268393 5253 268427 5287
rect 249073 4981 249107 5015
rect 224233 4913 224267 4947
rect 224141 4777 224175 4811
rect 224233 4777 224267 4811
rect 224141 4233 224175 4267
rect 249073 4233 249107 4267
rect 257997 4981 258031 5015
rect 268393 4981 268427 5015
rect 278053 5253 278087 5287
rect 278053 4981 278087 5015
rect 287713 4981 287747 5015
rect 297097 5457 297131 5491
rect 322673 5049 322707 5083
rect 297097 4981 297131 5015
rect 307033 4981 307067 5015
rect 257997 4233 258031 4267
rect 317337 4845 317371 4879
rect 317337 4709 317371 4743
rect 319453 4641 319487 4675
rect 322765 5049 322799 5083
rect 327181 5049 327215 5083
rect 322765 4845 322799 4879
rect 325157 4981 325191 5015
rect 325157 4777 325191 4811
rect 326169 4913 326203 4947
rect 326629 4777 326663 4811
rect 327181 4777 327215 4811
rect 326169 4641 326203 4675
rect 322673 4573 322707 4607
rect 326261 4573 326295 4607
rect 319453 4437 319487 4471
rect 471529 5593 471563 5627
rect 471437 5525 471471 5559
rect 466101 5253 466135 5287
rect 461225 5117 461259 5151
rect 466101 4913 466135 4947
rect 471345 5049 471379 5083
rect 461225 4845 461259 4879
rect 337117 4437 337151 4471
rect 376769 4777 376803 4811
rect 471345 4777 471379 4811
rect 471437 4777 471471 4811
rect 307033 4165 307067 4199
rect 269129 4097 269163 4131
rect 283113 4097 283147 4131
rect 283205 4097 283239 4131
rect 283205 3961 283239 3995
rect 283297 3961 283331 3995
rect 332333 4097 332367 4131
rect 269129 3893 269163 3927
rect 320833 3893 320867 3927
rect 285873 3757 285907 3791
rect 45477 3349 45511 3383
rect 282837 3349 282871 3383
rect 276305 3213 276339 3247
rect 45477 3145 45511 3179
rect 82921 3145 82955 3179
rect 276305 3009 276339 3043
rect 285873 3281 285907 3315
rect 292497 3689 292531 3723
rect 320741 3553 320775 3587
rect 320833 3553 320867 3587
rect 320925 3893 320959 3927
rect 326353 3893 326387 3927
rect 332241 3893 332275 3927
rect 332333 3893 332367 3927
rect 335369 4097 335403 4131
rect 326353 3689 326387 3723
rect 332149 3757 332183 3791
rect 332241 3757 332275 3791
rect 322765 3553 322799 3587
rect 332149 3553 332183 3587
rect 340889 4097 340923 4131
rect 349169 4097 349203 4131
rect 335921 3893 335955 3927
rect 335921 3689 335955 3723
rect 335369 3553 335403 3587
rect 335737 3553 335771 3587
rect 292497 3281 292531 3315
rect 322765 3077 322799 3111
rect 282837 3009 282871 3043
rect 335737 3009 335771 3043
rect 335829 3145 335863 3179
rect 340613 3145 340647 3179
rect 82921 2941 82955 2975
rect 93869 2941 93903 2975
rect 93869 2805 93903 2839
rect 335645 2941 335679 2975
rect 335829 2941 335863 2975
rect 340705 2873 340739 2907
rect 335645 2805 335679 2839
rect 344385 3349 344419 3383
rect 340797 2805 340831 2839
rect 343925 3213 343959 3247
rect 344109 3213 344143 3247
rect 345673 3349 345707 3383
rect 344385 2941 344419 2975
rect 345489 3281 345523 3315
rect 344109 2873 344143 2907
rect 343925 2805 343959 2839
rect 349169 3281 349203 3315
rect 352665 4097 352699 4131
rect 355241 4097 355275 4131
rect 355333 4097 355367 4131
rect 345673 3145 345707 3179
rect 347789 2941 347823 2975
rect 347789 2737 347823 2771
rect 350089 2941 350123 2975
rect 352665 2873 352699 2907
rect 352849 3621 352883 3655
rect 352941 3621 352975 3655
rect 352941 3349 352975 3383
rect 376769 3893 376803 3927
rect 376861 4369 376895 4403
rect 355425 3621 355459 3655
rect 361957 3689 361991 3723
rect 361957 3417 361991 3451
rect 362049 3689 362083 3723
rect 355333 3213 355367 3247
rect 355425 3213 355459 3247
rect 437489 4233 437523 4267
rect 418169 4097 418203 4131
rect 417525 3961 417559 3995
rect 376769 3485 376803 3519
rect 410993 3893 411027 3927
rect 417525 3689 417559 3723
rect 410993 3417 411027 3451
rect 413201 3485 413235 3519
rect 362049 3145 362083 3179
rect 365729 3145 365763 3179
rect 354873 2873 354907 2907
rect 365729 2873 365763 2907
rect 375297 3077 375331 3111
rect 375297 2873 375331 2907
rect 413201 2873 413235 2907
rect 352849 2805 352883 2839
rect 427737 4097 427771 4131
rect 420101 3961 420135 3995
rect 420101 3485 420135 3519
rect 422125 3689 422159 3723
rect 418169 2805 418203 2839
rect 423045 3689 423079 3723
rect 422953 3621 422987 3655
rect 423045 3485 423079 3519
rect 423137 3689 423171 3723
rect 423137 3213 423171 3247
rect 426449 3689 426483 3723
rect 426449 3145 426483 3179
rect 438225 4165 438259 4199
rect 438409 4165 438443 4199
rect 435925 3961 435959 3995
rect 437489 3961 437523 3995
rect 445861 4097 445895 4131
rect 430037 3689 430071 3723
rect 430037 3417 430071 3451
rect 430129 3689 430163 3723
rect 422953 3077 422987 3111
rect 423045 3077 423079 3111
rect 427737 3077 427771 3111
rect 423045 2873 423079 2907
rect 422125 2805 422159 2839
rect 350089 2737 350123 2771
rect 434545 3553 434579 3587
rect 434637 3553 434671 3587
rect 432521 3417 432555 3451
rect 432521 3077 432555 3111
rect 432613 3417 432647 3451
rect 451933 4097 451967 4131
rect 445861 3757 445895 3791
rect 446781 4029 446815 4063
rect 435925 3213 435959 3247
rect 441721 3689 441755 3723
rect 432613 2873 432647 2907
rect 451933 3825 451967 3859
rect 456809 3961 456843 3995
rect 466377 3757 466411 3791
rect 456809 3689 456843 3723
rect 456901 3689 456935 3723
rect 446781 3213 446815 3247
rect 449909 3621 449943 3655
rect 454693 3553 454727 3587
rect 449909 2941 449943 2975
rect 450277 3009 450311 3043
rect 450277 2873 450311 2907
rect 441721 2805 441755 2839
rect 444849 2805 444883 2839
rect 451197 2805 451231 2839
rect 451473 2805 451507 2839
rect 430129 2737 430163 2771
rect 345489 561 345523 595
rect 456809 2873 456843 2907
rect 466193 2873 466227 2907
rect 466377 2873 466411 2907
rect 466929 3757 466963 3791
rect 466929 2805 466963 2839
rect 466193 2737 466227 2771
rect 454693 2125 454727 2159
rect 444849 561 444883 595
rect 518173 3213 518207 3247
rect 518173 3009 518207 3043
rect 471529 561 471563 595
<< metal1 >>
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 358814 700992 358820 701004
rect 202840 700964 358820 700992
rect 202840 700952 202846 700964
rect 358814 700952 358820 700964
rect 358872 700952 358878 701004
rect 170306 700884 170312 700936
rect 170364 700924 170370 700936
rect 362954 700924 362960 700936
rect 170364 700896 362960 700924
rect 170364 700884 170370 700896
rect 362954 700884 362960 700896
rect 363012 700884 363018 700936
rect 328362 700816 328368 700868
rect 328420 700856 328426 700868
rect 527174 700856 527180 700868
rect 328420 700828 527180 700856
rect 328420 700816 328426 700828
rect 527174 700816 527180 700828
rect 527232 700816 527238 700868
rect 329742 700748 329748 700800
rect 329800 700788 329806 700800
rect 543458 700788 543464 700800
rect 329800 700760 543464 700788
rect 329800 700748 329806 700760
rect 543458 700748 543464 700760
rect 543516 700748 543522 700800
rect 154114 700680 154120 700732
rect 154172 700720 154178 700732
rect 367094 700720 367100 700732
rect 154172 700692 367100 700720
rect 154172 700680 154178 700692
rect 367094 700680 367100 700692
rect 367152 700680 367158 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 364334 700652 364340 700664
rect 137888 700624 364340 700652
rect 137888 700612 137894 700624
rect 364334 700612 364340 700624
rect 364392 700612 364398 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 368474 700584 368480 700596
rect 105504 700556 368480 700584
rect 105504 700544 105510 700556
rect 368474 700544 368480 700556
rect 368532 700544 368538 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 373994 700516 374000 700528
rect 89220 700488 374000 700516
rect 89220 700476 89226 700488
rect 373994 700476 374000 700488
rect 374052 700476 374058 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 371234 700448 371240 700460
rect 73028 700420 371240 700448
rect 73028 700408 73034 700420
rect 371234 700408 371240 700420
rect 371292 700408 371298 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 375374 700380 375380 700392
rect 40552 700352 375380 700380
rect 40552 700340 40558 700352
rect 375374 700340 375380 700352
rect 375432 700340 375438 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 379514 700312 379520 700324
rect 24360 700284 379520 700312
rect 24360 700272 24366 700284
rect 379514 700272 379520 700284
rect 379572 700272 379578 700324
rect 218974 700204 218980 700256
rect 219032 700244 219038 700256
rect 360194 700244 360200 700256
rect 219032 700216 360200 700244
rect 219032 700204 219038 700216
rect 360194 700204 360200 700216
rect 360252 700204 360258 700256
rect 336642 700136 336648 700188
rect 336700 700176 336706 700188
rect 478506 700176 478512 700188
rect 336700 700148 478512 700176
rect 336700 700136 336706 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 335262 700068 335268 700120
rect 335320 700108 335326 700120
rect 462314 700108 462320 700120
rect 335320 700080 462320 700108
rect 335320 700068 335326 700080
rect 462314 700068 462320 700080
rect 462372 700068 462378 700120
rect 235166 700000 235172 700052
rect 235224 700040 235230 700052
rect 356054 700040 356060 700052
rect 235224 700012 356060 700040
rect 235224 700000 235230 700012
rect 356054 700000 356060 700012
rect 356112 700000 356118 700052
rect 267642 699932 267648 699984
rect 267700 699972 267706 699984
rect 351914 699972 351920 699984
rect 267700 699944 351920 699972
rect 267700 699932 267706 699944
rect 351914 699932 351920 699944
rect 351972 699932 351978 699984
rect 283834 699864 283840 699916
rect 283892 699904 283898 699916
rect 354674 699904 354680 699916
rect 283892 699876 354680 699904
rect 283892 699864 283898 699876
rect 354674 699864 354680 699876
rect 354732 699864 354738 699916
rect 343542 699796 343548 699848
rect 343600 699836 343606 699848
rect 413646 699836 413652 699848
rect 343600 699808 413652 699836
rect 343600 699796 343606 699808
rect 413646 699796 413652 699808
rect 413704 699796 413710 699848
rect 340782 699728 340788 699780
rect 340840 699768 340846 699780
rect 397454 699768 397460 699780
rect 340840 699740 397460 699768
rect 340840 699728 340846 699740
rect 397454 699728 397460 699740
rect 397512 699728 397518 699780
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 332502 699660 332508 699712
rect 332560 699700 332566 699712
rect 346394 699700 346400 699712
rect 332560 699672 346400 699700
rect 332560 699660 332566 699672
rect 346394 699660 346400 699672
rect 346452 699660 346458 699712
rect 347774 699660 347780 699712
rect 347832 699700 347838 699712
rect 348786 699700 348792 699712
rect 347832 699672 348792 699700
rect 347832 699660 347838 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 321462 696940 321468 696992
rect 321520 696980 321526 696992
rect 580166 696980 580172 696992
rect 321520 696952 580172 696980
rect 321520 696940 321526 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 364610 687760 364616 687812
rect 364668 687800 364674 687812
rect 365162 687800 365168 687812
rect 364668 687772 365168 687800
rect 364668 687760 364674 687772
rect 365162 687760 365168 687772
rect 365220 687760 365226 687812
rect 429212 685936 429976 685964
rect 324222 685856 324228 685908
rect 324280 685896 324286 685908
rect 429212 685896 429240 685936
rect 324280 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 324280 685856 324286 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 364521 685831 364579 685837
rect 364521 685797 364533 685831
rect 364567 685828 364579 685831
rect 364610 685828 364616 685840
rect 364567 685800 364616 685828
rect 364567 685797 364579 685800
rect 364521 685791 364579 685797
rect 364610 685788 364616 685800
rect 364668 685788 364674 685840
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 382274 681748 382280 681760
rect 3568 681720 382280 681748
rect 3568 681708 3574 681720
rect 382274 681708 382280 681720
rect 382332 681708 382338 681760
rect 364518 676240 364524 676252
rect 364479 676212 364524 676240
rect 364518 676200 364524 676212
rect 364576 676200 364582 676252
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 320082 673480 320088 673532
rect 320140 673520 320146 673532
rect 580166 673520 580172 673532
rect 320140 673492 580172 673520
rect 320140 673480 320146 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 386414 667944 386420 667956
rect 3476 667916 386420 667944
rect 3476 667904 3482 667916
rect 386414 667904 386420 667916
rect 386472 667904 386478 667956
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 383654 652780 383660 652792
rect 3108 652752 383660 652780
rect 3108 652740 3114 652752
rect 383654 652740 383660 652752
rect 383712 652740 383718 652792
rect 315942 650020 315948 650072
rect 316000 650060 316006 650072
rect 580166 650060 580172 650072
rect 316000 650032 580172 650060
rect 316000 650020 316006 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 317322 638936 317328 638988
rect 317380 638976 317386 638988
rect 580166 638976 580172 638988
rect 317380 638948 580172 638976
rect 317380 638936 317386 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 313182 626560 313188 626612
rect 313240 626600 313246 626612
rect 580166 626600 580172 626612
rect 313240 626572 580172 626600
rect 313240 626560 313246 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 387794 623812 387800 623824
rect 3476 623784 387800 623812
rect 3476 623772 3482 623784
rect 387794 623772 387800 623784
rect 387852 623772 387858 623824
rect 364521 618239 364579 618245
rect 364521 618205 364533 618239
rect 364567 618236 364579 618239
rect 364610 618236 364616 618248
rect 364567 618208 364616 618236
rect 364567 618205 364579 618208
rect 364521 618199 364579 618205
rect 364610 618196 364616 618208
rect 364668 618196 364674 618248
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 391934 610008 391940 610020
rect 3476 609980 391940 610008
rect 3476 609968 3482 609980
rect 391934 609968 391940 609980
rect 391992 609968 391998 610020
rect 364518 608648 364524 608660
rect 364479 608620 364524 608648
rect 364518 608608 364524 608620
rect 364576 608608 364582 608660
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 309042 603100 309048 603152
rect 309100 603140 309106 603152
rect 580166 603140 580172 603152
rect 309100 603112 580172 603140
rect 309100 603100 309106 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 364610 598924 364616 598936
rect 364571 598896 364616 598924
rect 364610 598884 364616 598896
rect 364668 598884 364674 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 390554 594844 390560 594856
rect 3292 594816 390560 594844
rect 3292 594804 3298 594816
rect 390554 594804 390560 594816
rect 390612 594804 390618 594856
rect 311802 592016 311808 592068
rect 311860 592056 311866 592068
rect 580166 592056 580172 592068
rect 311860 592028 580172 592056
rect 311860 592016 311866 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 364613 589339 364671 589345
rect 364613 589305 364625 589339
rect 364659 589336 364671 589339
rect 364702 589336 364708 589348
rect 364659 589308 364708 589336
rect 364659 589305 364671 589308
rect 364613 589299 364671 589305
rect 364702 589296 364708 589308
rect 364760 589296 364766 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 344462 584672 344468 584724
rect 344520 584712 344526 584724
rect 364702 584712 364708 584724
rect 344520 584684 364708 584712
rect 344520 584672 344526 584684
rect 364702 584672 364708 584684
rect 364760 584672 364766 584724
rect 300762 584604 300768 584656
rect 300820 584644 300826 584656
rect 350810 584644 350816 584656
rect 300820 584616 350816 584644
rect 300820 584604 300826 584616
rect 350810 584604 350816 584616
rect 350868 584604 350874 584656
rect 338206 584536 338212 584588
rect 338264 584576 338270 584588
rect 429654 584576 429660 584588
rect 338264 584548 429660 584576
rect 338264 584536 338270 584548
rect 429654 584536 429660 584548
rect 429712 584536 429718 584588
rect 331858 584468 331864 584520
rect 331916 584508 331922 584520
rect 494238 584508 494244 584520
rect 331916 584480 494244 584508
rect 331916 584468 331922 584480
rect 494238 584468 494244 584480
rect 494296 584468 494302 584520
rect 325510 584400 325516 584452
rect 325568 584440 325574 584452
rect 559374 584440 559380 584452
rect 325568 584412 559380 584440
rect 325568 584400 325574 584412
rect 559374 584400 559380 584412
rect 559432 584400 559438 584452
rect 304534 583652 304540 583704
rect 304592 583692 304598 583704
rect 471422 583692 471428 583704
rect 304592 583664 471428 583692
rect 304592 583652 304598 583664
rect 471422 583652 471428 583664
rect 471480 583652 471486 583704
rect 298186 583584 298192 583636
rect 298244 583624 298250 583636
rect 471330 583624 471336 583636
rect 298244 583596 471336 583624
rect 298244 583584 298250 583596
rect 471330 583584 471336 583596
rect 471388 583584 471394 583636
rect 256050 583516 256056 583568
rect 256108 583556 256114 583568
rect 580626 583556 580632 583568
rect 256108 583528 580632 583556
rect 256108 583516 256114 583528
rect 580626 583516 580632 583528
rect 580684 583516 580690 583568
rect 245562 583448 245568 583500
rect 245620 583488 245626 583500
rect 580442 583488 580448 583500
rect 245620 583460 580448 583488
rect 245620 583448 245626 583460
rect 580442 583448 580448 583460
rect 580500 583448 580506 583500
rect 243446 583380 243452 583432
rect 243504 583420 243510 583432
rect 580258 583420 580264 583432
rect 243504 583392 580264 583420
rect 243504 583380 243510 583392
rect 580258 583380 580264 583392
rect 580316 583380 580322 583432
rect 4706 583312 4712 583364
rect 4764 583352 4770 583364
rect 399202 583352 399208 583364
rect 4764 583324 399208 583352
rect 4764 583312 4770 583324
rect 399202 583312 399208 583324
rect 399260 583312 399266 583364
rect 5442 583244 5448 583296
rect 5500 583284 5506 583296
rect 405550 583284 405556 583296
rect 5500 583256 405556 583284
rect 5500 583244 5506 583256
rect 405550 583244 405556 583256
rect 405608 583244 405614 583296
rect 10318 583176 10324 583228
rect 10376 583216 10382 583228
rect 411898 583216 411904 583228
rect 10376 583188 411904 583216
rect 10376 583176 10382 583188
rect 411898 583176 411904 583188
rect 411956 583176 411962 583228
rect 6270 583108 6276 583160
rect 6328 583148 6334 583160
rect 409782 583148 409788 583160
rect 6328 583120 409788 583148
rect 6328 583108 6334 583120
rect 409782 583108 409788 583120
rect 409840 583108 409846 583160
rect 3142 583040 3148 583092
rect 3200 583080 3206 583092
rect 407666 583080 407672 583092
rect 3200 583052 407672 583080
rect 3200 583040 3206 583052
rect 407666 583040 407672 583052
rect 407724 583040 407730 583092
rect 13078 582972 13084 583024
rect 13136 583012 13142 583024
rect 418154 583012 418160 583024
rect 13136 582984 418160 583012
rect 13136 582972 13142 582984
rect 418154 582972 418160 582984
rect 418212 582972 418218 583024
rect 14458 582904 14464 582956
rect 14516 582944 14522 582956
rect 424502 582944 424508 582956
rect 14516 582916 424508 582944
rect 14516 582904 14522 582916
rect 424502 582904 424508 582916
rect 424560 582904 424566 582956
rect 3234 582836 3240 582888
rect 3292 582876 3298 582888
rect 414014 582876 414020 582888
rect 3292 582848 414020 582876
rect 3292 582836 3298 582848
rect 414014 582836 414020 582848
rect 414072 582836 414078 582888
rect 5350 582768 5356 582820
rect 5408 582808 5414 582820
rect 422386 582808 422392 582820
rect 5408 582780 422392 582808
rect 5408 582768 5414 582780
rect 422386 582768 422392 582780
rect 422444 582768 422450 582820
rect 15838 582700 15844 582752
rect 15896 582740 15902 582752
rect 437106 582740 437112 582752
rect 15896 582712 437112 582740
rect 15896 582700 15902 582712
rect 437106 582700 437112 582712
rect 437164 582700 437170 582752
rect 4062 582632 4068 582684
rect 4120 582672 4126 582684
rect 430850 582672 430856 582684
rect 4120 582644 430856 582672
rect 4120 582632 4126 582644
rect 430850 582632 430856 582644
rect 430908 582632 430914 582684
rect 5258 582564 5264 582616
rect 5316 582604 5322 582616
rect 432966 582604 432972 582616
rect 5316 582576 432972 582604
rect 5316 582564 5322 582576
rect 432966 582564 432972 582576
rect 433024 582564 433030 582616
rect 3878 582496 3884 582548
rect 3936 582536 3942 582548
rect 434990 582536 434996 582548
rect 3936 582508 434996 582536
rect 3936 582496 3942 582508
rect 434990 582496 434996 582508
rect 435048 582496 435054 582548
rect 5166 582428 5172 582480
rect 5224 582468 5230 582480
rect 445570 582468 445576 582480
rect 5224 582440 445576 582468
rect 5224 582428 5230 582440
rect 445570 582428 445576 582440
rect 445628 582428 445634 582480
rect 3694 582360 3700 582412
rect 3752 582400 3758 582412
rect 443454 582400 443460 582412
rect 3752 582372 443460 582400
rect 3752 582360 3758 582372
rect 443454 582360 443460 582372
rect 443512 582360 443518 582412
rect 302418 581612 302424 581664
rect 302476 581652 302482 581664
rect 469582 581652 469588 581664
rect 302476 581624 469588 581652
rect 302476 581612 302482 581624
rect 469582 581612 469588 581624
rect 469640 581612 469646 581664
rect 296070 581544 296076 581596
rect 296128 581584 296134 581596
rect 469674 581584 469680 581596
rect 296128 581556 469680 581584
rect 296128 581544 296134 581556
rect 469674 581544 469680 581556
rect 469732 581544 469738 581596
rect 289722 581476 289728 581528
rect 289780 581516 289786 581528
rect 469766 581516 469772 581528
rect 289780 581488 469772 581516
rect 289780 581476 289786 581488
rect 469766 581476 469772 581488
rect 469824 581476 469830 581528
rect 287606 581408 287612 581460
rect 287664 581448 287670 581460
rect 470502 581448 470508 581460
rect 287664 581420 470508 581448
rect 287664 581408 287670 581420
rect 470502 581408 470508 581420
rect 470560 581408 470566 581460
rect 283466 581340 283472 581392
rect 283524 581380 283530 581392
rect 470410 581380 470416 581392
rect 283524 581352 470416 581380
rect 283524 581340 283530 581352
rect 470410 581340 470416 581352
rect 470468 581340 470474 581392
rect 281350 581272 281356 581324
rect 281408 581312 281414 581324
rect 470318 581312 470324 581324
rect 281408 581284 470324 581312
rect 281408 581272 281414 581284
rect 470318 581272 470324 581284
rect 470376 581272 470382 581324
rect 275002 581204 275008 581256
rect 275060 581244 275066 581256
rect 470226 581244 470232 581256
rect 275060 581216 470232 581244
rect 275060 581204 275066 581216
rect 470226 581204 470232 581216
rect 470284 581204 470290 581256
rect 268654 581136 268660 581188
rect 268712 581176 268718 581188
rect 470042 581176 470048 581188
rect 268712 581148 470048 581176
rect 268712 581136 268718 581148
rect 470042 581136 470048 581148
rect 470100 581136 470106 581188
rect 251818 581068 251824 581120
rect 251876 581108 251882 581120
rect 469858 581108 469864 581120
rect 251876 581080 469864 581108
rect 251876 581068 251882 581080
rect 469858 581068 469864 581080
rect 469916 581068 469922 581120
rect 264514 581000 264520 581052
rect 264572 581040 264578 581052
rect 580074 581040 580080 581052
rect 264572 581012 580080 581040
rect 264572 581000 264578 581012
rect 580074 581000 580080 581012
rect 580132 581000 580138 581052
rect 262398 580252 262404 580304
rect 262456 580292 262462 580304
rect 469950 580292 469956 580304
rect 262456 580264 469956 580292
rect 262456 580252 262462 580264
rect 469950 580252 469956 580264
rect 470008 580252 470014 580304
rect 306558 580184 306564 580236
rect 306616 580224 306622 580236
rect 580166 580224 580172 580236
rect 306616 580196 580172 580224
rect 306616 580184 306622 580196
rect 580166 580184 580172 580196
rect 580224 580184 580230 580236
rect 6638 580116 6644 580168
rect 6696 580156 6702 580168
rect 395062 580156 395068 580168
rect 6696 580128 395068 580156
rect 6696 580116 6702 580128
rect 395062 580116 395068 580128
rect 395120 580116 395126 580168
rect 6546 580048 6552 580100
rect 6604 580088 6610 580100
rect 397086 580088 397092 580100
rect 6604 580060 397092 580088
rect 6604 580048 6610 580060
rect 397086 580048 397092 580060
rect 397144 580048 397150 580100
rect 6454 579980 6460 580032
rect 6512 580020 6518 580032
rect 400950 580020 400956 580032
rect 6512 579992 400956 580020
rect 6512 579980 6518 579992
rect 400950 579980 400956 579992
rect 401008 579980 401014 580032
rect 6362 579912 6368 579964
rect 6420 579952 6426 579964
rect 403158 579952 403164 579964
rect 6420 579924 403164 579952
rect 6420 579912 6426 579924
rect 403158 579912 403164 579924
rect 403216 579912 403222 579964
rect 3786 579844 3792 579896
rect 3844 579884 3850 579896
rect 438854 579884 438860 579896
rect 3844 579856 438860 579884
rect 3844 579844 3850 579856
rect 438854 579844 438860 579856
rect 438912 579844 438918 579896
rect 4982 579776 4988 579828
rect 5040 579816 5046 579828
rect 451550 579816 451556 579828
rect 5040 579788 451556 579816
rect 5040 579776 5046 579788
rect 451550 579776 451556 579788
rect 451608 579776 451614 579828
rect 4890 579708 4896 579760
rect 4948 579748 4954 579760
rect 458266 579748 458272 579760
rect 4948 579720 458272 579748
rect 4948 579708 4954 579720
rect 458266 579708 458272 579720
rect 458324 579708 458330 579760
rect 6178 579640 6184 579692
rect 6236 579680 6242 579692
rect 464246 579680 464252 579692
rect 6236 579652 464252 579680
rect 6236 579640 6242 579652
rect 464246 579640 464252 579652
rect 464304 579640 464310 579692
rect 271138 579368 271144 579420
rect 271196 579408 271202 579420
rect 271196 579380 282224 579408
rect 271196 579368 271202 579380
rect 247954 579340 247960 579352
rect 247915 579312 247960 579340
rect 247954 579300 247960 579312
rect 248012 579300 248018 579352
rect 254210 579340 254216 579352
rect 254171 579312 254216 579340
rect 254210 579300 254216 579312
rect 254268 579300 254274 579352
rect 258442 579300 258448 579352
rect 258500 579300 258506 579352
rect 260650 579300 260656 579352
rect 260708 579300 260714 579352
rect 266906 579300 266912 579352
rect 266964 579300 266970 579352
rect 273162 579300 273168 579352
rect 273220 579300 273226 579352
rect 277302 579300 277308 579352
rect 277360 579300 277366 579352
rect 279602 579300 279608 579352
rect 279660 579300 279666 579352
rect 258460 578728 258488 579300
rect 260668 578796 260696 579300
rect 266924 578864 266952 579300
rect 273180 578932 273208 579300
rect 277320 579000 277348 579300
rect 279620 579068 279648 579300
rect 282196 579204 282224 579380
rect 285766 579300 285772 579352
rect 285824 579300 285830 579352
rect 292114 579340 292120 579352
rect 292075 579312 292120 579340
rect 292114 579300 292120 579312
rect 292172 579300 292178 579352
rect 415670 579340 415676 579352
rect 415631 579312 415676 579340
rect 415670 579300 415676 579312
rect 415728 579300 415734 579352
rect 428366 579340 428372 579352
rect 428327 579312 428372 579340
rect 428366 579300 428372 579312
rect 428424 579300 428430 579352
rect 441062 579340 441068 579352
rect 441023 579312 441068 579340
rect 441062 579300 441068 579312
rect 441120 579300 441126 579352
rect 453574 579340 453580 579352
rect 453535 579312 453580 579340
rect 453574 579300 453580 579312
rect 453632 579300 453638 579352
rect 455782 579340 455788 579352
rect 455743 579312 455788 579340
rect 455782 579300 455788 579312
rect 455840 579300 455846 579352
rect 285784 579272 285812 579300
rect 471238 579272 471244 579284
rect 285784 579244 471244 579272
rect 471238 579232 471244 579244
rect 471296 579232 471302 579284
rect 470134 579204 470140 579216
rect 282196 579176 470140 579204
rect 470134 579164 470140 579176
rect 470192 579164 470198 579216
rect 292117 579139 292175 579145
rect 292117 579105 292129 579139
rect 292163 579136 292175 579139
rect 579798 579136 579804 579148
rect 292163 579108 579804 579136
rect 292163 579105 292175 579108
rect 292117 579099 292175 579105
rect 579798 579096 579804 579108
rect 579856 579096 579862 579148
rect 579982 579068 579988 579080
rect 279620 579040 579988 579068
rect 579982 579028 579988 579040
rect 580040 579028 580046 579080
rect 579890 579000 579896 579012
rect 277320 578972 579896 579000
rect 579890 578960 579896 578972
rect 579948 578960 579954 579012
rect 580074 578932 580080 578944
rect 273180 578904 580080 578932
rect 580074 578892 580080 578904
rect 580132 578892 580138 578944
rect 580902 578864 580908 578876
rect 266924 578836 580908 578864
rect 580902 578824 580908 578836
rect 580960 578824 580966 578876
rect 580718 578796 580724 578808
rect 260668 578768 580724 578796
rect 580718 578756 580724 578768
rect 580776 578756 580782 578808
rect 580810 578728 580816 578740
rect 258460 578700 580816 578728
rect 580810 578688 580816 578700
rect 580868 578688 580874 578740
rect 254213 578663 254271 578669
rect 254213 578629 254225 578663
rect 254259 578660 254271 578663
rect 580534 578660 580540 578672
rect 254259 578632 580540 578660
rect 254259 578629 254271 578632
rect 254213 578623 254271 578629
rect 580534 578620 580540 578632
rect 580592 578620 580598 578672
rect 247957 578595 248015 578601
rect 247957 578561 247969 578595
rect 248003 578592 248015 578595
rect 580350 578592 580356 578604
rect 248003 578564 580356 578592
rect 248003 578561 248015 578564
rect 247957 578555 248015 578561
rect 580350 578552 580356 578564
rect 580408 578552 580414 578604
rect 3326 578484 3332 578536
rect 3384 578524 3390 578536
rect 415673 578527 415731 578533
rect 415673 578524 415685 578527
rect 3384 578496 415685 578524
rect 3384 578484 3390 578496
rect 415673 578493 415685 578496
rect 415719 578493 415731 578527
rect 415673 578487 415731 578493
rect 3970 578416 3976 578468
rect 4028 578456 4034 578468
rect 428369 578459 428427 578465
rect 428369 578456 428381 578459
rect 4028 578428 428381 578456
rect 4028 578416 4034 578428
rect 428369 578425 428381 578428
rect 428415 578425 428427 578459
rect 428369 578419 428427 578425
rect 3602 578348 3608 578400
rect 3660 578388 3666 578400
rect 441065 578391 441123 578397
rect 441065 578388 441077 578391
rect 3660 578360 441077 578388
rect 3660 578348 3666 578360
rect 441065 578357 441077 578360
rect 441111 578357 441123 578391
rect 441065 578351 441123 578357
rect 3418 578280 3424 578332
rect 3476 578320 3482 578332
rect 453577 578323 453635 578329
rect 453577 578320 453589 578323
rect 3476 578292 453589 578320
rect 3476 578280 3482 578292
rect 453577 578289 453589 578292
rect 453623 578289 453635 578323
rect 453577 578283 453635 578289
rect 3510 578212 3516 578264
rect 3568 578252 3574 578264
rect 455785 578255 455843 578261
rect 455785 578252 455797 578255
rect 3568 578224 455797 578252
rect 3568 578212 3574 578224
rect 455785 578221 455797 578224
rect 455831 578221 455843 578255
rect 455785 578215 455843 578221
rect 3050 567332 3056 567384
rect 3108 567372 3114 567384
rect 6638 567372 6644 567384
rect 3108 567344 6644 567372
rect 3108 567332 3114 567344
rect 6638 567332 6644 567344
rect 6696 567332 6702 567384
rect 469582 557472 469588 557524
rect 469640 557512 469646 557524
rect 579706 557512 579712 557524
rect 469640 557484 579712 557512
rect 469640 557472 469646 557484
rect 579706 557472 579712 557484
rect 579764 557472 579770 557524
rect 2774 553052 2780 553104
rect 2832 553092 2838 553104
rect 4706 553092 4712 553104
rect 2832 553064 4712 553092
rect 2832 553052 2838 553064
rect 4706 553052 4712 553064
rect 4764 553052 4770 553104
rect 471422 546388 471428 546440
rect 471480 546428 471486 546440
rect 579706 546428 579712 546440
rect 471480 546400 579712 546428
rect 471480 546388 471486 546400
rect 579706 546388 579712 546400
rect 579764 546388 579770 546440
rect 3050 538636 3056 538688
rect 3108 538676 3114 538688
rect 6546 538676 6552 538688
rect 3108 538648 6552 538676
rect 3108 538636 3114 538648
rect 6546 538636 6552 538648
rect 6604 538636 6610 538688
rect 469674 510552 469680 510604
rect 469732 510592 469738 510604
rect 579706 510592 579712 510604
rect 469732 510564 579712 510592
rect 469732 510552 469738 510564
rect 579706 510552 579712 510564
rect 579764 510552 579770 510604
rect 3050 510212 3056 510264
rect 3108 510252 3114 510264
rect 6454 510252 6460 510264
rect 3108 510224 6460 510252
rect 3108 510212 3114 510224
rect 6454 510212 6460 510224
rect 6512 510212 6518 510264
rect 471330 499468 471336 499520
rect 471388 499508 471394 499520
rect 579706 499508 579712 499520
rect 471388 499480 579712 499508
rect 471388 499468 471394 499480
rect 579706 499468 579712 499480
rect 579764 499468 579770 499520
rect 2774 496680 2780 496732
rect 2832 496720 2838 496732
rect 5442 496720 5448 496732
rect 2832 496692 5448 496720
rect 2832 496680 2838 496692
rect 5442 496680 5448 496692
rect 5500 496680 5506 496732
rect 2958 481108 2964 481160
rect 3016 481148 3022 481160
rect 6362 481148 6368 481160
rect 3016 481120 6368 481148
rect 3016 481108 3022 481120
rect 6362 481108 6368 481120
rect 6420 481108 6426 481160
rect 469766 463632 469772 463684
rect 469824 463672 469830 463684
rect 579706 463672 579712 463684
rect 469824 463644 579712 463672
rect 469824 463632 469830 463644
rect 579706 463632 579712 463644
rect 579764 463632 579770 463684
rect 470502 440172 470508 440224
rect 470560 440212 470566 440224
rect 579798 440212 579804 440224
rect 470560 440184 579804 440212
rect 470560 440172 470566 440184
rect 579798 440172 579804 440184
rect 579856 440172 579862 440224
rect 3142 438812 3148 438864
rect 3200 438852 3206 438864
rect 10318 438852 10324 438864
rect 3200 438824 10324 438852
rect 3200 438812 3206 438824
rect 10318 438812 10324 438824
rect 10376 438812 10382 438864
rect 3142 424056 3148 424108
rect 3200 424096 3206 424108
rect 6270 424096 6276 424108
rect 3200 424068 6276 424096
rect 3200 424056 3206 424068
rect 6270 424056 6276 424068
rect 6328 424056 6334 424108
rect 470410 416712 470416 416764
rect 470468 416752 470474 416764
rect 579798 416752 579804 416764
rect 470468 416724 579804 416752
rect 470468 416712 470474 416724
rect 579798 416712 579804 416724
rect 579856 416712 579862 416764
rect 471238 405628 471244 405680
rect 471296 405668 471302 405680
rect 579798 405668 579804 405680
rect 471296 405640 579804 405668
rect 471296 405628 471302 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 470318 393252 470324 393304
rect 470376 393292 470382 393304
rect 579798 393292 579804 393304
rect 470376 393264 579804 393292
rect 470376 393252 470382 393264
rect 579798 393252 579804 393264
rect 579856 393252 579862 393304
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 13078 380848 13084 380860
rect 3292 380820 13084 380848
rect 3292 380808 3298 380820
rect 13078 380808 13084 380820
rect 13136 380808 13142 380860
rect 470226 346332 470232 346384
rect 470284 346372 470290 346384
rect 579982 346372 579988 346384
rect 470284 346344 579988 346372
rect 470284 346332 470290 346344
rect 579982 346332 579988 346344
rect 580040 346332 580046 346384
rect 346397 338691 346455 338697
rect 346397 338657 346409 338691
rect 346443 338688 346455 338691
rect 348510 338688 348516 338700
rect 346443 338660 348516 338688
rect 346443 338657 346455 338660
rect 346397 338651 346455 338657
rect 348510 338648 348516 338660
rect 348568 338648 348574 338700
rect 316126 338104 316132 338156
rect 316184 338144 316190 338156
rect 316310 338144 316316 338156
rect 316184 338116 316316 338144
rect 316184 338104 316190 338116
rect 316310 338104 316316 338116
rect 316368 338104 316374 338156
rect 318794 338104 318800 338156
rect 318852 338144 318858 338156
rect 319806 338144 319812 338156
rect 318852 338116 319812 338144
rect 318852 338104 318858 338116
rect 319806 338104 319812 338116
rect 319864 338104 319870 338156
rect 327077 338147 327135 338153
rect 327077 338113 327089 338147
rect 327123 338144 327135 338147
rect 336645 338147 336703 338153
rect 336645 338144 336657 338147
rect 327123 338116 336657 338144
rect 327123 338113 327135 338116
rect 327077 338107 327135 338113
rect 336645 338113 336657 338116
rect 336691 338113 336703 338147
rect 336645 338107 336703 338113
rect 340322 338104 340328 338156
rect 340380 338144 340386 338156
rect 340690 338144 340696 338156
rect 340380 338116 340696 338144
rect 340380 338104 340386 338116
rect 340690 338104 340696 338116
rect 340748 338104 340754 338156
rect 442353 338147 442411 338153
rect 442353 338144 442365 338147
rect 442184 338116 442365 338144
rect 71038 338036 71044 338088
rect 71096 338076 71102 338088
rect 254946 338076 254952 338088
rect 71096 338048 254952 338076
rect 71096 338036 71102 338048
rect 254946 338036 254952 338048
rect 255004 338036 255010 338088
rect 314654 338036 314660 338088
rect 314712 338076 314718 338088
rect 315390 338076 315396 338088
rect 314712 338048 315396 338076
rect 314712 338036 314718 338048
rect 315390 338036 315396 338048
rect 315448 338036 315454 338088
rect 315485 338079 315543 338085
rect 315485 338045 315497 338079
rect 315531 338076 315543 338079
rect 318889 338079 318947 338085
rect 318889 338076 318901 338079
rect 315531 338048 318901 338076
rect 315531 338045 315543 338048
rect 315485 338039 315543 338045
rect 318889 338045 318901 338048
rect 318935 338045 318947 338079
rect 318889 338039 318947 338045
rect 319073 338079 319131 338085
rect 319073 338045 319085 338079
rect 319119 338076 319131 338079
rect 354398 338076 354404 338088
rect 319119 338048 354404 338076
rect 319119 338045 319131 338048
rect 319073 338039 319131 338045
rect 354398 338036 354404 338048
rect 354456 338036 354462 338088
rect 358078 338036 358084 338088
rect 358136 338076 358142 338088
rect 371510 338076 371516 338088
rect 358136 338048 371516 338076
rect 358136 338036 358142 338048
rect 371510 338036 371516 338048
rect 371568 338036 371574 338088
rect 372709 338079 372767 338085
rect 372709 338045 372721 338079
rect 372755 338076 372767 338079
rect 378870 338076 378876 338088
rect 372755 338048 378876 338076
rect 372755 338045 372767 338048
rect 372709 338039 372767 338045
rect 378870 338036 378876 338048
rect 378928 338036 378934 338088
rect 403342 338036 403348 338088
rect 403400 338076 403406 338088
rect 412453 338079 412511 338085
rect 412453 338076 412465 338079
rect 403400 338048 412465 338076
rect 403400 338036 403406 338048
rect 412453 338045 412465 338048
rect 412499 338045 412511 338079
rect 412453 338039 412511 338045
rect 414658 338036 414664 338088
rect 414716 338076 414722 338088
rect 429838 338076 429844 338088
rect 414716 338048 429844 338076
rect 414716 338036 414722 338048
rect 429838 338036 429844 338048
rect 429896 338036 429902 338088
rect 432509 338079 432567 338085
rect 432509 338045 432521 338079
rect 432555 338076 432567 338079
rect 442184 338076 442212 338116
rect 442353 338113 442365 338116
rect 442399 338113 442411 338147
rect 442353 338107 442411 338113
rect 432555 338048 442212 338076
rect 442261 338079 442319 338085
rect 432555 338045 432567 338048
rect 432509 338039 432567 338045
rect 442261 338045 442273 338079
rect 442307 338076 442319 338079
rect 483014 338076 483020 338088
rect 442307 338048 483020 338076
rect 442307 338045 442319 338048
rect 442261 338039 442319 338045
rect 483014 338036 483020 338048
rect 483072 338036 483078 338088
rect 483109 338079 483167 338085
rect 483109 338045 483121 338079
rect 483155 338045 483167 338079
rect 483109 338039 483167 338045
rect 66898 337968 66904 338020
rect 66956 338008 66962 338020
rect 96065 338011 96123 338017
rect 96065 338008 96077 338011
rect 66956 337980 96077 338008
rect 66956 337968 66962 337980
rect 96065 337977 96077 337980
rect 96111 337977 96123 338011
rect 96065 337971 96123 337977
rect 96249 338011 96307 338017
rect 96249 337977 96261 338011
rect 96295 338008 96307 338011
rect 115385 338011 115443 338017
rect 115385 338008 115397 338011
rect 96295 337980 115397 338008
rect 96295 337977 96307 337980
rect 96249 337971 96307 337977
rect 115385 337977 115397 337980
rect 115431 337977 115443 338011
rect 115385 337971 115443 337977
rect 115569 338011 115627 338017
rect 115569 337977 115581 338011
rect 115615 338008 115627 338011
rect 134705 338011 134763 338017
rect 134705 338008 134717 338011
rect 115615 337980 134717 338008
rect 115615 337977 115627 337980
rect 115569 337971 115627 337977
rect 134705 337977 134717 337980
rect 134751 337977 134763 338011
rect 134705 337971 134763 337977
rect 134889 338011 134947 338017
rect 134889 337977 134901 338011
rect 134935 338008 134947 338011
rect 154025 338011 154083 338017
rect 154025 338008 154037 338011
rect 134935 337980 154037 338008
rect 134935 337977 134947 337980
rect 134889 337971 134947 337977
rect 154025 337977 154037 337980
rect 154071 337977 154083 338011
rect 154025 337971 154083 337977
rect 154209 338011 154267 338017
rect 154209 337977 154221 338011
rect 154255 338008 154267 338011
rect 173345 338011 173403 338017
rect 173345 338008 173357 338011
rect 154255 337980 173357 338008
rect 154255 337977 154267 337980
rect 154209 337971 154267 337977
rect 173345 337977 173357 337980
rect 173391 337977 173403 338011
rect 173345 337971 173403 337977
rect 173529 338011 173587 338017
rect 173529 337977 173541 338011
rect 173575 338008 173587 338011
rect 192665 338011 192723 338017
rect 192665 338008 192677 338011
rect 173575 337980 192677 338008
rect 173575 337977 173587 337980
rect 173529 337971 173587 337977
rect 192665 337977 192677 337980
rect 192711 337977 192723 338011
rect 192665 337971 192723 337977
rect 192849 338011 192907 338017
rect 192849 337977 192861 338011
rect 192895 338008 192907 338011
rect 211985 338011 212043 338017
rect 211985 338008 211997 338011
rect 192895 337980 211997 338008
rect 192895 337977 192907 337980
rect 192849 337971 192907 337977
rect 211985 337977 211997 337980
rect 212031 337977 212043 338011
rect 211985 337971 212043 337977
rect 212169 338011 212227 338017
rect 212169 337977 212181 338011
rect 212215 338008 212227 338011
rect 252002 338008 252008 338020
rect 212215 337980 252008 338008
rect 212215 337977 212227 337980
rect 212169 337971 212227 337977
rect 252002 337968 252008 337980
rect 252060 337968 252066 338020
rect 306190 337968 306196 338020
rect 306248 338008 306254 338020
rect 355870 338008 355876 338020
rect 306248 337980 355876 338008
rect 306248 337968 306254 337980
rect 355870 337968 355876 337980
rect 355928 337968 355934 338020
rect 364242 337968 364248 338020
rect 364300 338008 364306 338020
rect 379330 338008 379336 338020
rect 364300 337980 379336 338008
rect 364300 337968 364306 337980
rect 379330 337968 379336 337980
rect 379388 337968 379394 338020
rect 397454 337968 397460 338020
rect 397512 338008 397518 338020
rect 403618 338008 403624 338020
rect 397512 337980 403624 338008
rect 397512 337968 397518 337980
rect 403618 337968 403624 337980
rect 403676 337968 403682 338020
rect 406286 337968 406292 338020
rect 406344 338008 406350 338020
rect 417418 338008 417424 338020
rect 406344 337980 417424 338008
rect 406344 337968 406350 337980
rect 417418 337968 417424 337980
rect 417476 337968 417482 338020
rect 424962 337968 424968 338020
rect 425020 338008 425026 338020
rect 430025 338011 430083 338017
rect 430025 338008 430037 338011
rect 425020 337980 430037 338008
rect 425020 337968 425026 337980
rect 430025 337977 430037 337980
rect 430071 337977 430083 338011
rect 430025 337971 430083 337977
rect 430114 337968 430120 338020
rect 430172 338008 430178 338020
rect 434073 338011 434131 338017
rect 434073 338008 434085 338011
rect 430172 337980 434085 338008
rect 430172 337968 430178 337980
rect 434073 337977 434085 337980
rect 434119 337977 434131 338011
rect 434073 337971 434131 337977
rect 444377 338011 444435 338017
rect 444377 337977 444389 338011
rect 444423 338008 444435 338011
rect 452013 338011 452071 338017
rect 452013 338008 452025 338011
rect 444423 337980 452025 338008
rect 444423 337977 444435 337980
rect 444377 337971 444435 337977
rect 452013 337977 452025 337980
rect 452059 337977 452071 338011
rect 452013 337971 452071 337977
rect 454770 337968 454776 338020
rect 454828 338008 454834 338020
rect 455877 338011 455935 338017
rect 455877 338008 455889 338011
rect 454828 337980 455889 338008
rect 454828 337968 454834 337980
rect 455877 337977 455889 337980
rect 455923 337977 455935 338011
rect 455877 337971 455935 337977
rect 459738 337968 459744 338020
rect 459796 338008 459802 338020
rect 460842 338008 460848 338020
rect 459796 337980 460848 338008
rect 459796 337968 459802 337980
rect 460842 337968 460848 337980
rect 460900 337968 460906 338020
rect 483124 338008 483152 338039
rect 483382 338036 483388 338088
rect 483440 338076 483446 338088
rect 499574 338076 499580 338088
rect 483440 338048 499580 338076
rect 483440 338036 483446 338048
rect 499574 338036 499580 338048
rect 499632 338036 499638 338088
rect 463528 337980 483152 338008
rect 483201 338011 483259 338017
rect 61378 337900 61384 337952
rect 61436 337940 61442 337952
rect 247586 337940 247592 337952
rect 61436 337912 247592 337940
rect 61436 337900 61442 337912
rect 247586 337900 247592 337912
rect 247644 337900 247650 337952
rect 258718 337900 258724 337952
rect 258776 337940 258782 337952
rect 272610 337940 272616 337952
rect 258776 337912 272616 337940
rect 258776 337900 258782 337912
rect 272610 337900 272616 337912
rect 272668 337900 272674 337952
rect 303154 337900 303160 337952
rect 303212 337940 303218 337952
rect 318889 337943 318947 337949
rect 318889 337940 318901 337943
rect 303212 337912 318901 337940
rect 303212 337900 303218 337912
rect 318889 337909 318901 337912
rect 318935 337909 318947 337943
rect 318889 337903 318947 337909
rect 318981 337943 319039 337949
rect 318981 337909 318993 337943
rect 319027 337940 319039 337943
rect 352926 337940 352932 337952
rect 319027 337912 352932 337940
rect 319027 337909 319039 337912
rect 318981 337903 319039 337909
rect 352926 337900 352932 337912
rect 352984 337900 352990 337952
rect 355318 337900 355324 337952
rect 355376 337940 355382 337952
rect 370038 337940 370044 337952
rect 355376 337912 370044 337940
rect 355376 337900 355382 337912
rect 370038 337900 370044 337912
rect 370096 337900 370102 337952
rect 374641 337943 374699 337949
rect 374641 337909 374653 337943
rect 374687 337940 374699 337943
rect 380342 337940 380348 337952
rect 374687 337912 380348 337940
rect 374687 337909 374699 337912
rect 374641 337903 374699 337909
rect 380342 337900 380348 337912
rect 380400 337900 380406 337952
rect 400398 337900 400404 337952
rect 400456 337940 400462 337952
rect 413278 337940 413284 337952
rect 400456 337912 413284 337940
rect 400456 337900 400462 337912
rect 413278 337900 413284 337912
rect 413336 337900 413342 337952
rect 413646 337900 413652 337952
rect 413704 337940 413710 337952
rect 420270 337940 420276 337952
rect 413704 337912 420276 337940
rect 413704 337900 413710 337912
rect 420270 337900 420276 337912
rect 420328 337900 420334 337952
rect 431310 337900 431316 337952
rect 431368 337940 431374 337952
rect 434533 337943 434591 337949
rect 434533 337940 434545 337943
rect 431368 337912 434545 337940
rect 431368 337900 431374 337912
rect 434533 337909 434545 337912
rect 434579 337909 434591 337943
rect 434533 337903 434591 337909
rect 435726 337900 435732 337952
rect 435784 337940 435790 337952
rect 442261 337943 442319 337949
rect 442261 337940 442273 337943
rect 435784 337912 442273 337940
rect 435784 337900 435790 337912
rect 442261 337909 442273 337912
rect 442307 337909 442319 337943
rect 442261 337903 442319 337909
rect 442353 337943 442411 337949
rect 442353 337909 442365 337943
rect 442399 337940 442411 337943
rect 442399 337912 451780 337940
rect 442399 337909 442411 337912
rect 442353 337903 442411 337909
rect 57238 337832 57244 337884
rect 57296 337872 57302 337884
rect 96249 337875 96307 337881
rect 96249 337872 96261 337875
rect 57296 337844 96261 337872
rect 57296 337832 57302 337844
rect 96249 337841 96261 337844
rect 96295 337841 96307 337875
rect 96249 337835 96307 337841
rect 96433 337875 96491 337881
rect 96433 337841 96445 337875
rect 96479 337872 96491 337875
rect 115569 337875 115627 337881
rect 115569 337872 115581 337875
rect 96479 337844 115581 337872
rect 96479 337841 96491 337844
rect 96433 337835 96491 337841
rect 115569 337841 115581 337844
rect 115615 337841 115627 337875
rect 115569 337835 115627 337841
rect 115753 337875 115811 337881
rect 115753 337841 115765 337875
rect 115799 337872 115811 337875
rect 134889 337875 134947 337881
rect 134889 337872 134901 337875
rect 115799 337844 134901 337872
rect 115799 337841 115811 337844
rect 115753 337835 115811 337841
rect 134889 337841 134901 337844
rect 134935 337841 134947 337875
rect 134889 337835 134947 337841
rect 135073 337875 135131 337881
rect 135073 337841 135085 337875
rect 135119 337872 135131 337875
rect 154209 337875 154267 337881
rect 154209 337872 154221 337875
rect 135119 337844 154221 337872
rect 135119 337841 135131 337844
rect 135073 337835 135131 337841
rect 154209 337841 154221 337844
rect 154255 337841 154267 337875
rect 154209 337835 154267 337841
rect 154393 337875 154451 337881
rect 154393 337841 154405 337875
rect 154439 337872 154451 337875
rect 173529 337875 173587 337881
rect 173529 337872 173541 337875
rect 154439 337844 173541 337872
rect 154439 337841 154451 337844
rect 154393 337835 154451 337841
rect 173529 337841 173541 337844
rect 173575 337841 173587 337875
rect 173529 337835 173587 337841
rect 173713 337875 173771 337881
rect 173713 337841 173725 337875
rect 173759 337872 173771 337875
rect 192849 337875 192907 337881
rect 192849 337872 192861 337875
rect 173759 337844 192861 337872
rect 173759 337841 173771 337844
rect 173713 337835 173771 337841
rect 192849 337841 192861 337844
rect 192895 337841 192907 337875
rect 192849 337835 192907 337841
rect 193033 337875 193091 337881
rect 193033 337841 193045 337875
rect 193079 337872 193091 337875
rect 212169 337875 212227 337881
rect 212169 337872 212181 337875
rect 193079 337844 212181 337872
rect 193079 337841 193091 337844
rect 193033 337835 193091 337841
rect 212169 337841 212181 337844
rect 212215 337841 212227 337875
rect 212169 337835 212227 337841
rect 212353 337875 212411 337881
rect 212353 337841 212365 337875
rect 212399 337872 212411 337875
rect 247126 337872 247132 337884
rect 212399 337844 247132 337872
rect 212399 337841 212411 337844
rect 212353 337835 212411 337841
rect 247126 337832 247132 337844
rect 247184 337832 247190 337884
rect 290458 337832 290464 337884
rect 290516 337872 290522 337884
rect 335909 337875 335967 337881
rect 335909 337872 335921 337875
rect 290516 337844 335921 337872
rect 290516 337832 290522 337844
rect 335909 337841 335921 337844
rect 335955 337841 335967 337875
rect 335909 337835 335967 337841
rect 336001 337875 336059 337881
rect 336001 337841 336013 337875
rect 336047 337872 336059 337875
rect 347038 337872 347044 337884
rect 336047 337844 347044 337872
rect 336047 337841 336059 337844
rect 336001 337835 336059 337841
rect 347038 337832 347044 337844
rect 347096 337832 347102 337884
rect 348418 337832 348424 337884
rect 348476 337872 348482 337884
rect 365622 337872 365628 337884
rect 348476 337844 365628 337872
rect 348476 337832 348482 337844
rect 365622 337832 365628 337844
rect 365680 337832 365686 337884
rect 411714 337832 411720 337884
rect 411772 337872 411778 337884
rect 412542 337872 412548 337884
rect 411772 337844 412548 337872
rect 411772 337832 411778 337844
rect 412542 337832 412548 337844
rect 412600 337832 412606 337884
rect 416056 337844 416820 337872
rect 50338 337764 50344 337816
rect 50396 337804 50402 337816
rect 244182 337804 244188 337816
rect 50396 337776 244188 337804
rect 50396 337764 50402 337776
rect 244182 337764 244188 337776
rect 244240 337764 244246 337816
rect 259638 337764 259644 337816
rect 259696 337804 259702 337816
rect 260098 337804 260104 337816
rect 259696 337776 260104 337804
rect 259696 337764 259702 337776
rect 260098 337764 260104 337776
rect 260156 337764 260162 337816
rect 288250 337764 288256 337816
rect 288308 337804 288314 337816
rect 302145 337807 302203 337813
rect 302145 337804 302157 337807
rect 288308 337776 302157 337804
rect 288308 337764 288314 337776
rect 302145 337773 302157 337776
rect 302191 337773 302203 337807
rect 302145 337767 302203 337773
rect 303985 337807 304043 337813
rect 303985 337773 303997 337807
rect 304031 337804 304043 337807
rect 318797 337807 318855 337813
rect 318797 337804 318809 337807
rect 304031 337776 318809 337804
rect 304031 337773 304043 337776
rect 303985 337767 304043 337773
rect 318797 337773 318809 337776
rect 318843 337773 318855 337807
rect 318797 337767 318855 337773
rect 318981 337807 319039 337813
rect 318981 337773 318993 337807
rect 319027 337804 319039 337807
rect 351914 337804 351920 337816
rect 319027 337776 351920 337804
rect 319027 337773 319039 337776
rect 318981 337767 319039 337773
rect 351914 337764 351920 337776
rect 351972 337764 351978 337816
rect 362862 337764 362868 337816
rect 362920 337804 362926 337816
rect 372709 337807 372767 337813
rect 372709 337804 372721 337807
rect 362920 337776 372721 337804
rect 362920 337764 362926 337776
rect 372709 337773 372721 337776
rect 372755 337773 372767 337807
rect 377398 337804 377404 337816
rect 372709 337767 372767 337773
rect 372816 337776 377404 337804
rect 39298 337696 39304 337748
rect 39356 337736 39362 337748
rect 57974 337736 57980 337748
rect 39356 337708 57980 337736
rect 39356 337696 39362 337708
rect 57974 337696 57980 337708
rect 58032 337696 58038 337748
rect 67542 337696 67548 337748
rect 67600 337736 67606 337748
rect 241517 337739 241575 337745
rect 241517 337736 241529 337739
rect 67600 337708 241529 337736
rect 67600 337696 67606 337708
rect 241517 337705 241529 337708
rect 241563 337705 241575 337739
rect 241517 337699 241575 337705
rect 249058 337696 249064 337748
rect 249116 337736 249122 337748
rect 250530 337736 250536 337748
rect 249116 337708 250536 337736
rect 249116 337696 249122 337708
rect 250530 337696 250536 337708
rect 250588 337696 250594 337748
rect 251450 337696 251456 337748
rect 251508 337736 251514 337748
rect 252462 337736 252468 337748
rect 251508 337708 252468 337736
rect 251508 337696 251514 337708
rect 252462 337696 252468 337708
rect 252520 337696 252526 337748
rect 254578 337696 254584 337748
rect 254636 337736 254642 337748
rect 262306 337736 262312 337748
rect 254636 337708 262312 337736
rect 254636 337696 254642 337708
rect 262306 337696 262312 337708
rect 262364 337696 262370 337748
rect 302237 337739 302295 337745
rect 302237 337705 302249 337739
rect 302283 337736 302295 337739
rect 307754 337736 307760 337748
rect 302283 337708 307760 337736
rect 302283 337705 302295 337708
rect 302237 337699 302295 337705
rect 307754 337696 307760 337708
rect 307812 337696 307818 337748
rect 317322 337696 317328 337748
rect 317380 337736 317386 337748
rect 327077 337739 327135 337745
rect 327077 337736 327089 337739
rect 317380 337708 327089 337736
rect 317380 337696 317386 337708
rect 327077 337705 327089 337708
rect 327123 337705 327135 337739
rect 327077 337699 327135 337705
rect 336645 337739 336703 337745
rect 336645 337705 336657 337739
rect 336691 337736 336703 337739
rect 346397 337739 346455 337745
rect 346397 337736 346409 337739
rect 336691 337708 346409 337736
rect 336691 337705 336703 337708
rect 336645 337699 336703 337705
rect 346397 337705 346409 337708
rect 346443 337705 346455 337739
rect 346397 337699 346455 337705
rect 356698 337696 356704 337748
rect 356756 337736 356762 337748
rect 360746 337736 360752 337748
rect 356756 337708 360752 337736
rect 356756 337696 356762 337708
rect 360746 337696 360752 337708
rect 360804 337696 360810 337748
rect 372816 337736 372844 337776
rect 377398 337764 377404 337776
rect 377456 337764 377462 337816
rect 388438 337764 388444 337816
rect 388496 337804 388502 337816
rect 389174 337804 389180 337816
rect 388496 337776 389180 337804
rect 388496 337764 388502 337776
rect 389174 337764 389180 337776
rect 389232 337764 389238 337816
rect 396074 337764 396080 337816
rect 396132 337804 396138 337816
rect 398190 337804 398196 337816
rect 396132 337776 398196 337804
rect 396132 337764 396138 337776
rect 398190 337764 398196 337776
rect 398248 337764 398254 337816
rect 404354 337764 404360 337816
rect 404412 337804 404418 337816
rect 416056 337804 416084 337844
rect 404412 337776 416084 337804
rect 404412 337764 404418 337776
rect 416130 337764 416136 337816
rect 416188 337804 416194 337816
rect 416682 337804 416688 337816
rect 416188 337776 416688 337804
rect 416188 337764 416194 337776
rect 416682 337764 416688 337776
rect 416740 337764 416746 337816
rect 416792 337804 416820 337844
rect 417602 337832 417608 337884
rect 417660 337872 417666 337884
rect 434257 337875 434315 337881
rect 434257 337872 434269 337875
rect 417660 337844 434269 337872
rect 417660 337832 417666 337844
rect 434257 337841 434269 337844
rect 434303 337841 434315 337875
rect 434257 337835 434315 337841
rect 434441 337875 434499 337881
rect 434441 337841 434453 337875
rect 434487 337872 434499 337875
rect 449437 337875 449495 337881
rect 449437 337872 449449 337875
rect 434487 337844 449449 337872
rect 434487 337841 434499 337844
rect 434441 337835 434499 337841
rect 449437 337841 449449 337844
rect 449483 337841 449495 337875
rect 451752 337872 451780 337912
rect 451826 337900 451832 337952
rect 451884 337940 451890 337952
rect 461489 337943 461547 337949
rect 461489 337940 461501 337943
rect 451884 337912 461501 337940
rect 451884 337900 451890 337912
rect 461489 337909 461501 337912
rect 461535 337909 461547 337943
rect 461489 337903 461547 337909
rect 456705 337875 456763 337881
rect 456705 337872 456717 337875
rect 451752 337844 456717 337872
rect 449437 337835 449495 337841
rect 456705 337841 456717 337844
rect 456751 337841 456763 337875
rect 456705 337835 456763 337841
rect 460658 337832 460664 337884
rect 460716 337872 460722 337884
rect 463528 337872 463556 337980
rect 483201 337977 483213 338011
rect 483247 338008 483259 338011
rect 525058 338008 525064 338020
rect 483247 337980 525064 338008
rect 483247 337977 483259 337980
rect 483201 337971 483259 337977
rect 525058 337968 525064 337980
rect 525116 337968 525122 338020
rect 463602 337900 463608 337952
rect 463660 337940 463666 337952
rect 466365 337943 466423 337949
rect 466365 337940 466377 337943
rect 463660 337912 466377 337940
rect 463660 337900 463666 337912
rect 466365 337909 466377 337912
rect 466411 337909 466423 337943
rect 466365 337903 466423 337909
rect 467098 337900 467104 337952
rect 467156 337940 467162 337952
rect 467742 337940 467748 337952
rect 467156 337912 467748 337940
rect 467156 337900 467162 337912
rect 467742 337900 467748 337912
rect 467800 337900 467806 337952
rect 468018 337900 468024 337952
rect 468076 337940 468082 337952
rect 469122 337940 469128 337952
rect 468076 337912 469128 337940
rect 468076 337900 468082 337912
rect 469122 337900 469128 337912
rect 469180 337900 469186 337952
rect 469217 337943 469275 337949
rect 469217 337909 469229 337943
rect 469263 337940 469275 337943
rect 483109 337943 483167 337949
rect 483109 337940 483121 337943
rect 469263 337912 483121 337940
rect 469263 337909 469275 337912
rect 469217 337903 469275 337909
rect 483109 337909 483121 337912
rect 483155 337909 483167 337943
rect 483109 337903 483167 337909
rect 483293 337943 483351 337949
rect 483293 337909 483305 337943
rect 483339 337940 483351 337943
rect 527818 337940 527824 337952
rect 483339 337912 527824 337940
rect 483339 337909 483351 337912
rect 483293 337903 483351 337909
rect 527818 337900 527824 337912
rect 527876 337900 527882 337952
rect 460716 337844 463556 337872
rect 463697 337875 463755 337881
rect 460716 337832 460722 337844
rect 463697 337841 463709 337875
rect 463743 337872 463755 337875
rect 483014 337872 483020 337884
rect 463743 337844 483020 337872
rect 463743 337841 463755 337844
rect 463697 337835 463755 337841
rect 483014 337832 483020 337844
rect 483072 337832 483078 337884
rect 483382 337832 483388 337884
rect 483440 337872 483446 337884
rect 523678 337872 523684 337884
rect 483440 337844 523684 337872
rect 483440 337832 483446 337844
rect 523678 337832 523684 337844
rect 523736 337832 523742 337884
rect 420178 337804 420184 337816
rect 416792 337776 420184 337804
rect 420178 337764 420184 337776
rect 420236 337764 420242 337816
rect 422018 337764 422024 337816
rect 422076 337804 422082 337816
rect 432601 337807 432659 337813
rect 432601 337804 432613 337807
rect 422076 337776 432613 337804
rect 422076 337764 422082 337776
rect 432601 337773 432613 337776
rect 432647 337773 432659 337807
rect 432601 337767 432659 337773
rect 438670 337764 438676 337816
rect 438728 337804 438734 337816
rect 438728 337776 442948 337804
rect 438728 337764 438734 337776
rect 375926 337736 375932 337748
rect 361592 337708 372844 337736
rect 372908 337708 375932 337736
rect 32398 337628 32404 337680
rect 32456 337668 32462 337680
rect 230569 337671 230627 337677
rect 230569 337668 230581 337671
rect 32456 337640 230581 337668
rect 32456 337628 32462 337640
rect 230569 337637 230581 337640
rect 230615 337637 230627 337671
rect 230569 337631 230627 337637
rect 230658 337628 230664 337680
rect 230716 337668 230722 337680
rect 231118 337668 231124 337680
rect 230716 337640 231124 337668
rect 230716 337628 230722 337640
rect 231118 337628 231124 337640
rect 231176 337628 231182 337680
rect 231213 337671 231271 337677
rect 231213 337637 231225 337671
rect 231259 337668 231271 337671
rect 234433 337671 234491 337677
rect 234433 337668 234445 337671
rect 231259 337640 234445 337668
rect 231259 337637 231271 337640
rect 231213 337631 231271 337637
rect 234433 337637 234445 337640
rect 234479 337637 234491 337671
rect 234433 337631 234491 337637
rect 255958 337628 255964 337680
rect 256016 337668 256022 337680
rect 259733 337671 259791 337677
rect 259733 337668 259745 337671
rect 256016 337640 259745 337668
rect 256016 337628 256022 337640
rect 259733 337637 259745 337640
rect 259779 337637 259791 337671
rect 259733 337631 259791 337637
rect 260098 337628 260104 337680
rect 260156 337668 260162 337680
rect 277026 337668 277032 337680
rect 260156 337640 277032 337668
rect 260156 337628 260162 337640
rect 277026 337628 277032 337640
rect 277084 337628 277090 337680
rect 285582 337628 285588 337680
rect 285640 337668 285646 337680
rect 336001 337671 336059 337677
rect 336001 337668 336013 337671
rect 285640 337640 336013 337668
rect 285640 337628 285646 337640
rect 336001 337637 336013 337640
rect 336047 337637 336059 337671
rect 336001 337631 336059 337637
rect 336090 337628 336096 337680
rect 336148 337668 336154 337680
rect 344554 337668 344560 337680
rect 336148 337640 344560 337668
rect 336148 337628 336154 337640
rect 344554 337628 344560 337640
rect 344612 337628 344618 337680
rect 344649 337671 344707 337677
rect 344649 337637 344661 337671
rect 344695 337668 344707 337671
rect 349982 337668 349988 337680
rect 344695 337640 349988 337668
rect 344695 337637 344707 337640
rect 344649 337631 344707 337637
rect 349982 337628 349988 337640
rect 350040 337628 350046 337680
rect 354858 337668 354864 337680
rect 350276 337640 354864 337668
rect 35158 337560 35164 337612
rect 35216 337600 35222 337612
rect 96341 337603 96399 337609
rect 96341 337600 96353 337603
rect 35216 337572 96353 337600
rect 35216 337560 35222 337572
rect 96341 337569 96353 337572
rect 96387 337569 96399 337603
rect 96341 337563 96399 337569
rect 96525 337603 96583 337609
rect 96525 337569 96537 337603
rect 96571 337600 96583 337603
rect 115661 337603 115719 337609
rect 115661 337600 115673 337603
rect 96571 337572 115673 337600
rect 96571 337569 96583 337572
rect 96525 337563 96583 337569
rect 115661 337569 115673 337572
rect 115707 337569 115719 337603
rect 115661 337563 115719 337569
rect 115845 337603 115903 337609
rect 115845 337569 115857 337603
rect 115891 337600 115903 337603
rect 134981 337603 135039 337609
rect 134981 337600 134993 337603
rect 115891 337572 134993 337600
rect 115891 337569 115903 337572
rect 115845 337563 115903 337569
rect 134981 337569 134993 337572
rect 135027 337569 135039 337603
rect 134981 337563 135039 337569
rect 135165 337603 135223 337609
rect 135165 337569 135177 337603
rect 135211 337600 135223 337603
rect 154301 337603 154359 337609
rect 154301 337600 154313 337603
rect 135211 337572 154313 337600
rect 135211 337569 135223 337572
rect 135165 337563 135223 337569
rect 154301 337569 154313 337572
rect 154347 337569 154359 337603
rect 154301 337563 154359 337569
rect 154485 337603 154543 337609
rect 154485 337569 154497 337603
rect 154531 337600 154543 337603
rect 173621 337603 173679 337609
rect 173621 337600 173633 337603
rect 154531 337572 173633 337600
rect 154531 337569 154543 337572
rect 154485 337563 154543 337569
rect 173621 337569 173633 337572
rect 173667 337569 173679 337603
rect 173621 337563 173679 337569
rect 173805 337603 173863 337609
rect 173805 337569 173817 337603
rect 173851 337600 173863 337603
rect 192941 337603 192999 337609
rect 192941 337600 192953 337603
rect 173851 337572 192953 337600
rect 173851 337569 173863 337572
rect 173805 337563 173863 337569
rect 192941 337569 192953 337572
rect 192987 337569 192999 337603
rect 192941 337563 192999 337569
rect 193125 337603 193183 337609
rect 193125 337569 193137 337603
rect 193171 337600 193183 337603
rect 212261 337603 212319 337609
rect 212261 337600 212273 337603
rect 193171 337572 212273 337600
rect 193171 337569 193183 337572
rect 193125 337563 193183 337569
rect 212261 337569 212273 337572
rect 212307 337569 212319 337603
rect 212261 337563 212319 337569
rect 212445 337603 212503 337609
rect 212445 337569 212457 337603
rect 212491 337600 212503 337603
rect 241698 337600 241704 337612
rect 212491 337572 241704 337600
rect 212491 337569 212503 337572
rect 212445 337563 212503 337569
rect 241698 337560 241704 337572
rect 241756 337560 241762 337612
rect 261386 337560 261392 337612
rect 261444 337600 261450 337612
rect 279970 337600 279976 337612
rect 261444 337572 279976 337600
rect 261444 337560 261450 337572
rect 279970 337560 279976 337572
rect 280028 337560 280034 337612
rect 281442 337560 281448 337612
rect 281500 337600 281506 337612
rect 318889 337603 318947 337609
rect 318889 337600 318901 337603
rect 281500 337572 318901 337600
rect 281500 337560 281506 337572
rect 318889 337569 318901 337572
rect 318935 337569 318947 337603
rect 318889 337563 318947 337569
rect 318981 337603 319039 337609
rect 318981 337569 318993 337603
rect 319027 337600 319039 337603
rect 345566 337600 345572 337612
rect 319027 337572 345572 337600
rect 319027 337569 319039 337572
rect 318981 337563 319039 337569
rect 345566 337560 345572 337572
rect 345624 337560 345630 337612
rect 345750 337560 345756 337612
rect 345808 337600 345814 337612
rect 350166 337600 350172 337612
rect 345808 337572 350172 337600
rect 345808 337560 345814 337572
rect 350166 337560 350172 337572
rect 350224 337560 350230 337612
rect 28258 337492 28264 337544
rect 28316 337532 28322 337544
rect 96249 337535 96307 337541
rect 96249 337532 96261 337535
rect 28316 337504 96261 337532
rect 28316 337492 28322 337504
rect 96249 337501 96261 337504
rect 96295 337501 96307 337535
rect 96249 337495 96307 337501
rect 96433 337535 96491 337541
rect 96433 337501 96445 337535
rect 96479 337532 96491 337535
rect 115569 337535 115627 337541
rect 115569 337532 115581 337535
rect 96479 337504 115581 337532
rect 96479 337501 96491 337504
rect 96433 337495 96491 337501
rect 115569 337501 115581 337504
rect 115615 337501 115627 337535
rect 115569 337495 115627 337501
rect 115753 337535 115811 337541
rect 115753 337501 115765 337535
rect 115799 337532 115811 337535
rect 134889 337535 134947 337541
rect 134889 337532 134901 337535
rect 115799 337504 134901 337532
rect 115799 337501 115811 337504
rect 115753 337495 115811 337501
rect 134889 337501 134901 337504
rect 134935 337501 134947 337535
rect 134889 337495 134947 337501
rect 135073 337535 135131 337541
rect 135073 337501 135085 337535
rect 135119 337532 135131 337535
rect 154209 337535 154267 337541
rect 154209 337532 154221 337535
rect 135119 337504 154221 337532
rect 135119 337501 135131 337504
rect 135073 337495 135131 337501
rect 154209 337501 154221 337504
rect 154255 337501 154267 337535
rect 154209 337495 154267 337501
rect 154393 337535 154451 337541
rect 154393 337501 154405 337535
rect 154439 337532 154451 337535
rect 173529 337535 173587 337541
rect 173529 337532 173541 337535
rect 154439 337504 173541 337532
rect 154439 337501 154451 337504
rect 154393 337495 154451 337501
rect 173529 337501 173541 337504
rect 173575 337501 173587 337535
rect 173529 337495 173587 337501
rect 173713 337535 173771 337541
rect 173713 337501 173725 337535
rect 173759 337532 173771 337535
rect 192849 337535 192907 337541
rect 192849 337532 192861 337535
rect 173759 337504 192861 337532
rect 173759 337501 173771 337504
rect 173713 337495 173771 337501
rect 192849 337501 192861 337504
rect 192895 337501 192907 337535
rect 192849 337495 192907 337501
rect 193033 337535 193091 337541
rect 193033 337501 193045 337535
rect 193079 337532 193091 337535
rect 212169 337535 212227 337541
rect 212169 337532 212181 337535
rect 193079 337504 212181 337532
rect 193079 337501 193091 337504
rect 193033 337495 193091 337501
rect 212169 337501 212181 337504
rect 212215 337501 212227 337535
rect 212169 337495 212227 337501
rect 212353 337535 212411 337541
rect 212353 337501 212365 337535
rect 212399 337532 212411 337535
rect 230477 337535 230535 337541
rect 230477 337532 230489 337535
rect 212399 337504 230489 337532
rect 212399 337501 212411 337504
rect 212353 337495 212411 337501
rect 230477 337501 230489 337504
rect 230523 337501 230535 337535
rect 230477 337495 230535 337501
rect 230569 337535 230627 337541
rect 230569 337501 230581 337535
rect 230615 337532 230627 337535
rect 237834 337532 237840 337544
rect 230615 337504 237840 337532
rect 230615 337501 230627 337504
rect 230569 337495 230627 337501
rect 237834 337492 237840 337504
rect 237892 337492 237898 337544
rect 241517 337535 241575 337541
rect 241517 337501 241529 337535
rect 241563 337532 241575 337535
rect 244642 337532 244648 337544
rect 241563 337504 244648 337532
rect 241563 337501 241575 337504
rect 241517 337495 241575 337501
rect 244642 337492 244648 337504
rect 244700 337492 244706 337544
rect 253198 337492 253204 337544
rect 253256 337532 253262 337544
rect 259362 337532 259368 337544
rect 253256 337504 259368 337532
rect 253256 337492 253262 337504
rect 259362 337492 259368 337504
rect 259420 337492 259426 337544
rect 275554 337532 275560 337544
rect 259472 337504 275560 337532
rect 19978 337424 19984 337476
rect 20036 337464 20042 337476
rect 96157 337467 96215 337473
rect 96157 337464 96169 337467
rect 20036 337436 96169 337464
rect 20036 337424 20042 337436
rect 96157 337433 96169 337436
rect 96203 337433 96215 337467
rect 96157 337427 96215 337433
rect 96341 337467 96399 337473
rect 96341 337433 96353 337467
rect 96387 337464 96399 337467
rect 115477 337467 115535 337473
rect 115477 337464 115489 337467
rect 96387 337436 115489 337464
rect 96387 337433 96399 337436
rect 96341 337427 96399 337433
rect 115477 337433 115489 337436
rect 115523 337433 115535 337467
rect 115477 337427 115535 337433
rect 115661 337467 115719 337473
rect 115661 337433 115673 337467
rect 115707 337464 115719 337467
rect 134797 337467 134855 337473
rect 134797 337464 134809 337467
rect 115707 337436 134809 337464
rect 115707 337433 115719 337436
rect 115661 337427 115719 337433
rect 134797 337433 134809 337436
rect 134843 337433 134855 337467
rect 134797 337427 134855 337433
rect 134981 337467 135039 337473
rect 134981 337433 134993 337467
rect 135027 337464 135039 337467
rect 154117 337467 154175 337473
rect 154117 337464 154129 337467
rect 135027 337436 154129 337464
rect 135027 337433 135039 337436
rect 134981 337427 135039 337433
rect 154117 337433 154129 337436
rect 154163 337433 154175 337467
rect 154117 337427 154175 337433
rect 154301 337467 154359 337473
rect 154301 337433 154313 337467
rect 154347 337464 154359 337467
rect 173437 337467 173495 337473
rect 173437 337464 173449 337467
rect 154347 337436 173449 337464
rect 154347 337433 154359 337436
rect 154301 337427 154359 337433
rect 173437 337433 173449 337436
rect 173483 337433 173495 337467
rect 173437 337427 173495 337433
rect 173621 337467 173679 337473
rect 173621 337433 173633 337467
rect 173667 337464 173679 337467
rect 192757 337467 192815 337473
rect 192757 337464 192769 337467
rect 173667 337436 192769 337464
rect 173667 337433 173679 337436
rect 173621 337427 173679 337433
rect 192757 337433 192769 337436
rect 192803 337433 192815 337467
rect 192757 337427 192815 337433
rect 192941 337467 192999 337473
rect 192941 337433 192953 337467
rect 192987 337464 192999 337467
rect 212077 337467 212135 337473
rect 212077 337464 212089 337467
rect 192987 337436 212089 337464
rect 192987 337433 192999 337436
rect 192941 337427 192999 337433
rect 212077 337433 212089 337436
rect 212123 337433 212135 337467
rect 212077 337427 212135 337433
rect 212261 337467 212319 337473
rect 212261 337433 212273 337467
rect 212307 337464 212319 337467
rect 234338 337464 234344 337476
rect 212307 337436 234344 337464
rect 212307 337433 212319 337436
rect 212261 337427 212319 337433
rect 234338 337424 234344 337436
rect 234396 337424 234402 337476
rect 234433 337467 234491 337473
rect 234433 337433 234445 337467
rect 234479 337464 234491 337467
rect 238294 337464 238300 337476
rect 234479 337436 238300 337464
rect 234479 337433 234491 337436
rect 234433 337427 234491 337433
rect 238294 337424 238300 337436
rect 238352 337424 238358 337476
rect 258810 337424 258816 337476
rect 258868 337464 258874 337476
rect 259472 337464 259500 337504
rect 275554 337492 275560 337504
rect 275612 337492 275618 337544
rect 275922 337492 275928 337544
rect 275980 337532 275986 337544
rect 335817 337535 335875 337541
rect 335817 337532 335829 337535
rect 275980 337504 335829 337532
rect 275980 337492 275986 337504
rect 335817 337501 335829 337504
rect 335863 337501 335875 337535
rect 341610 337532 341616 337544
rect 335817 337495 335875 337501
rect 336016 337504 341616 337532
rect 269666 337464 269672 337476
rect 258868 337436 259500 337464
rect 259656 337436 269672 337464
rect 258868 337424 258874 337436
rect 13078 337356 13084 337408
rect 13136 337396 13142 337408
rect 115385 337399 115443 337405
rect 115385 337396 115397 337399
rect 13136 337368 115397 337396
rect 13136 337356 13142 337368
rect 115385 337365 115397 337368
rect 115431 337365 115443 337399
rect 115385 337359 115443 337365
rect 115845 337399 115903 337405
rect 115845 337365 115857 337399
rect 115891 337396 115903 337399
rect 134705 337399 134763 337405
rect 134705 337396 134717 337399
rect 115891 337368 134717 337396
rect 115891 337365 115903 337368
rect 115845 337359 115903 337365
rect 134705 337365 134717 337368
rect 134751 337365 134763 337399
rect 134705 337359 134763 337365
rect 135165 337399 135223 337405
rect 135165 337365 135177 337399
rect 135211 337396 135223 337399
rect 154025 337399 154083 337405
rect 154025 337396 154037 337399
rect 135211 337368 154037 337396
rect 135211 337365 135223 337368
rect 135165 337359 135223 337365
rect 154025 337365 154037 337368
rect 154071 337365 154083 337399
rect 154025 337359 154083 337365
rect 154485 337399 154543 337405
rect 154485 337365 154497 337399
rect 154531 337396 154543 337399
rect 173345 337399 173403 337405
rect 173345 337396 173357 337399
rect 154531 337368 173357 337396
rect 154531 337365 154543 337368
rect 154485 337359 154543 337365
rect 173345 337365 173357 337368
rect 173391 337365 173403 337399
rect 173345 337359 173403 337365
rect 173805 337399 173863 337405
rect 173805 337365 173817 337399
rect 173851 337396 173863 337399
rect 192665 337399 192723 337405
rect 192665 337396 192677 337399
rect 173851 337368 192677 337396
rect 173851 337365 173863 337368
rect 173805 337359 173863 337365
rect 192665 337365 192677 337368
rect 192711 337365 192723 337399
rect 192665 337359 192723 337365
rect 193125 337399 193183 337405
rect 193125 337365 193137 337399
rect 193171 337396 193183 337399
rect 211985 337399 212043 337405
rect 211985 337396 211997 337399
rect 193171 337368 211997 337396
rect 193171 337365 193183 337368
rect 193125 337359 193183 337365
rect 211985 337365 211997 337368
rect 212031 337365 212043 337399
rect 211985 337359 212043 337365
rect 212445 337399 212503 337405
rect 212445 337365 212457 337399
rect 212491 337396 212503 337399
rect 233510 337396 233516 337408
rect 212491 337368 233516 337396
rect 212491 337365 212503 337368
rect 212445 337359 212503 337365
rect 233510 337356 233516 337368
rect 233568 337356 233574 337408
rect 233878 337356 233884 337408
rect 233936 337396 233942 337408
rect 241238 337396 241244 337408
rect 233936 337368 241244 337396
rect 233936 337356 233942 337368
rect 241238 337356 241244 337368
rect 241296 337356 241302 337408
rect 250438 337356 250444 337408
rect 250496 337396 250502 337408
rect 253474 337396 253480 337408
rect 250496 337368 253480 337396
rect 250496 337356 250502 337368
rect 253474 337356 253480 337368
rect 253532 337356 253538 337408
rect 257338 337356 257344 337408
rect 257396 337396 257402 337408
rect 259656 337396 259684 337436
rect 269666 337424 269672 337436
rect 269724 337424 269730 337476
rect 271782 337424 271788 337476
rect 271840 337464 271846 337476
rect 318797 337467 318855 337473
rect 318797 337464 318809 337467
rect 271840 337436 318809 337464
rect 271840 337424 271846 337436
rect 318797 337433 318809 337436
rect 318843 337433 318855 337467
rect 318797 337427 318855 337433
rect 319073 337467 319131 337473
rect 319073 337433 319085 337467
rect 319119 337464 319131 337467
rect 336016 337464 336044 337504
rect 341610 337492 341616 337504
rect 341668 337492 341674 337544
rect 341705 337535 341763 337541
rect 341705 337501 341717 337535
rect 341751 337532 341763 337535
rect 342714 337532 342720 337544
rect 341751 337504 342720 337532
rect 341751 337501 341763 337504
rect 341705 337495 341763 337501
rect 342714 337492 342720 337504
rect 342772 337492 342778 337544
rect 342809 337535 342867 337541
rect 342809 337501 342821 337535
rect 342855 337532 342867 337535
rect 344281 337535 344339 337541
rect 344281 337532 344293 337535
rect 342855 337504 344293 337532
rect 342855 337501 342867 337504
rect 342809 337495 342867 337501
rect 344281 337501 344293 337504
rect 344327 337501 344339 337535
rect 344281 337495 344339 337501
rect 344370 337492 344376 337544
rect 344428 337532 344434 337544
rect 350276 337532 350304 337640
rect 354858 337628 354864 337640
rect 354916 337628 354922 337680
rect 358722 337628 358728 337680
rect 358780 337668 358786 337680
rect 361592 337668 361620 337708
rect 358780 337640 361620 337668
rect 364981 337671 365039 337677
rect 358780 337628 358786 337640
rect 364981 337637 364993 337671
rect 365027 337668 365039 337671
rect 372908 337668 372936 337708
rect 375926 337696 375932 337708
rect 375984 337696 375990 337748
rect 392578 337696 392584 337748
rect 392636 337736 392642 337748
rect 393222 337736 393228 337748
rect 392636 337708 393228 337736
rect 392636 337696 392642 337708
rect 393222 337696 393228 337708
rect 393280 337696 393286 337748
rect 394050 337696 394056 337748
rect 394108 337736 394114 337748
rect 394602 337736 394608 337748
rect 394108 337708 394608 337736
rect 394108 337696 394114 337708
rect 394602 337696 394608 337708
rect 394660 337696 394666 337748
rect 396534 337696 396540 337748
rect 396592 337736 396598 337748
rect 398098 337736 398104 337748
rect 396592 337708 398104 337736
rect 396592 337696 396598 337708
rect 398098 337696 398104 337708
rect 398156 337696 398162 337748
rect 410242 337696 410248 337748
rect 410300 337736 410306 337748
rect 411162 337736 411168 337748
rect 410300 337708 411168 337736
rect 410300 337696 410306 337708
rect 411162 337696 411168 337708
rect 411220 337696 411226 337748
rect 411254 337696 411260 337748
rect 411312 337736 411318 337748
rect 412358 337736 412364 337748
rect 411312 337708 412364 337736
rect 411312 337696 411318 337708
rect 412358 337696 412364 337708
rect 412416 337696 412422 337748
rect 412453 337739 412511 337745
rect 412453 337705 412465 337739
rect 412499 337736 412511 337739
rect 414109 337739 414167 337745
rect 414109 337736 414121 337739
rect 412499 337708 414121 337736
rect 412499 337705 412511 337708
rect 412453 337699 412511 337705
rect 414109 337705 414121 337708
rect 414155 337705 414167 337739
rect 414109 337699 414167 337705
rect 414198 337696 414204 337748
rect 414256 337736 414262 337748
rect 415302 337736 415308 337748
rect 414256 337708 415308 337736
rect 414256 337696 414262 337708
rect 415302 337696 415308 337708
rect 415360 337696 415366 337748
rect 415578 337696 415584 337748
rect 415636 337736 415642 337748
rect 416498 337736 416504 337748
rect 415636 337708 416504 337736
rect 415636 337696 415642 337708
rect 416498 337696 416504 337708
rect 416556 337696 416562 337748
rect 417050 337696 417056 337748
rect 417108 337736 417114 337748
rect 417970 337736 417976 337748
rect 417108 337708 417976 337736
rect 417108 337696 417114 337708
rect 417970 337696 417976 337708
rect 418028 337696 418034 337748
rect 425422 337696 425428 337748
rect 425480 337736 425486 337748
rect 428458 337736 428464 337748
rect 425480 337708 428464 337736
rect 425480 337696 425486 337708
rect 428458 337696 428464 337708
rect 428516 337696 428522 337748
rect 430025 337739 430083 337745
rect 430025 337705 430037 337739
rect 430071 337736 430083 337739
rect 434533 337739 434591 337745
rect 430071 337708 432828 337736
rect 430071 337705 430083 337708
rect 430025 337699 430083 337705
rect 365027 337640 372936 337668
rect 365027 337637 365039 337640
rect 364981 337631 365039 337637
rect 373902 337628 373908 337680
rect 373960 337668 373966 337680
rect 383286 337668 383292 337680
rect 373960 337640 383292 337668
rect 373960 337628 373966 337640
rect 383286 337628 383292 337640
rect 383344 337628 383350 337680
rect 393590 337628 393596 337680
rect 393648 337668 393654 337680
rect 397454 337668 397460 337680
rect 393648 337640 397460 337668
rect 393648 337628 393654 337640
rect 397454 337628 397460 337640
rect 397512 337628 397518 337680
rect 398006 337628 398012 337680
rect 398064 337668 398070 337680
rect 399478 337668 399484 337680
rect 398064 337640 399484 337668
rect 398064 337628 398070 337640
rect 399478 337628 399484 337640
rect 399536 337628 399542 337680
rect 404814 337628 404820 337680
rect 404872 337668 404878 337680
rect 424318 337668 424324 337680
rect 404872 337640 424324 337668
rect 404872 337628 404878 337640
rect 424318 337628 424324 337640
rect 424376 337628 424382 337680
rect 426434 337628 426440 337680
rect 426492 337668 426498 337680
rect 432693 337671 432751 337677
rect 432693 337668 432705 337671
rect 426492 337640 432705 337668
rect 426492 337628 426498 337640
rect 432693 337637 432705 337640
rect 432739 337637 432751 337671
rect 432800 337668 432828 337708
rect 434533 337705 434545 337739
rect 434579 337736 434591 337739
rect 434579 337708 437428 337736
rect 434579 337705 434591 337708
rect 434533 337699 434591 337705
rect 437293 337671 437351 337677
rect 437293 337668 437305 337671
rect 432800 337640 437305 337668
rect 432693 337631 432751 337637
rect 437293 337637 437305 337640
rect 437339 337637 437351 337671
rect 437400 337668 437428 337708
rect 437474 337696 437480 337748
rect 437532 337736 437538 337748
rect 442350 337736 442356 337748
rect 437532 337708 442356 337736
rect 437532 337696 437538 337708
rect 442350 337696 442356 337708
rect 442408 337696 442414 337748
rect 442920 337736 442948 337776
rect 446030 337764 446036 337816
rect 446088 337804 446094 337816
rect 451921 337807 451979 337813
rect 451921 337804 451933 337807
rect 446088 337776 451933 337804
rect 446088 337764 446094 337776
rect 451921 337773 451933 337776
rect 451967 337773 451979 337807
rect 451921 337767 451979 337773
rect 452013 337807 452071 337813
rect 452013 337773 452025 337807
rect 452059 337804 452071 337807
rect 455690 337804 455696 337816
rect 452059 337776 455696 337804
rect 452059 337773 452071 337776
rect 452013 337767 452071 337773
rect 455690 337764 455696 337776
rect 455748 337764 455754 337816
rect 455877 337807 455935 337813
rect 455877 337773 455889 337807
rect 455923 337804 455935 337807
rect 483109 337807 483167 337813
rect 483109 337804 483121 337807
rect 455923 337776 483121 337804
rect 455923 337773 455935 337776
rect 455877 337767 455935 337773
rect 483109 337773 483121 337776
rect 483155 337773 483167 337807
rect 483109 337767 483167 337773
rect 483293 337807 483351 337813
rect 483293 337773 483305 337807
rect 483339 337804 483351 337807
rect 520918 337804 520924 337816
rect 483339 337776 520924 337804
rect 483339 337773 483351 337776
rect 483293 337767 483351 337773
rect 520918 337764 520924 337776
rect 520976 337764 520982 337816
rect 483014 337736 483020 337748
rect 442920 337708 483020 337736
rect 483014 337696 483020 337708
rect 483072 337696 483078 337748
rect 483382 337696 483388 337748
rect 483440 337736 483446 337748
rect 506474 337736 506480 337748
rect 483440 337708 506480 337736
rect 483440 337696 483446 337708
rect 506474 337696 506480 337708
rect 506532 337696 506538 337748
rect 449437 337671 449495 337677
rect 437400 337640 442488 337668
rect 437293 337631 437351 337637
rect 351178 337560 351184 337612
rect 351236 337600 351242 337612
rect 365349 337603 365407 337609
rect 365349 337600 365361 337603
rect 351236 337572 365361 337600
rect 351236 337560 351242 337572
rect 365349 337569 365361 337572
rect 365395 337569 365407 337603
rect 365349 337563 365407 337569
rect 371142 337560 371148 337612
rect 371200 337600 371206 337612
rect 382274 337600 382280 337612
rect 371200 337572 382280 337600
rect 371200 337560 371206 337572
rect 382274 337560 382280 337572
rect 382332 337560 382338 337612
rect 398926 337560 398932 337612
rect 398984 337600 398990 337612
rect 406378 337600 406384 337612
rect 398984 337572 406384 337600
rect 398984 337560 398990 337572
rect 406378 337560 406384 337572
rect 406436 337560 406442 337612
rect 407298 337560 407304 337612
rect 407356 337600 407362 337612
rect 427078 337600 427084 337612
rect 407356 337572 427084 337600
rect 407356 337560 407362 337572
rect 427078 337560 427084 337572
rect 427136 337560 427142 337612
rect 427906 337560 427912 337612
rect 427964 337600 427970 337612
rect 427964 337572 432736 337600
rect 427964 337560 427970 337572
rect 344428 337504 350304 337532
rect 344428 337492 344434 337504
rect 351822 337492 351828 337544
rect 351880 337532 351886 337544
rect 365073 337535 365131 337541
rect 365073 337532 365085 337535
rect 351880 337504 365085 337532
rect 351880 337492 351886 337504
rect 365073 337501 365085 337504
rect 365119 337501 365131 337535
rect 365073 337495 365131 337501
rect 365257 337535 365315 337541
rect 365257 337501 365269 337535
rect 365303 337532 365315 337535
rect 374454 337532 374460 337544
rect 365303 337504 374460 337532
rect 365303 337501 365315 337504
rect 365257 337495 365315 337501
rect 374454 337492 374460 337504
rect 374512 337492 374518 337544
rect 375282 337492 375288 337544
rect 375340 337532 375346 337544
rect 383746 337532 383752 337544
rect 375340 337504 383752 337532
rect 375340 337492 375346 337504
rect 383746 337492 383752 337504
rect 383804 337492 383810 337544
rect 395062 337492 395068 337544
rect 395120 337532 395126 337544
rect 395890 337532 395896 337544
rect 395120 337504 395896 337532
rect 395120 337492 395126 337504
rect 395890 337492 395896 337504
rect 395948 337492 395954 337544
rect 405826 337492 405832 337544
rect 405884 337532 405890 337544
rect 426434 337532 426440 337544
rect 405884 337504 426440 337532
rect 405884 337492 405890 337504
rect 426434 337492 426440 337504
rect 426492 337492 426498 337544
rect 432509 337535 432567 337541
rect 432509 337532 432521 337535
rect 426544 337504 432521 337532
rect 344094 337464 344100 337476
rect 319119 337436 336044 337464
rect 336108 337436 344100 337464
rect 319119 337433 319131 337436
rect 319073 337427 319131 337433
rect 257396 337368 259684 337396
rect 259733 337399 259791 337405
rect 257396 337356 257402 337368
rect 259733 337365 259745 337399
rect 259779 337396 259791 337399
rect 266722 337396 266728 337408
rect 259779 337368 266728 337396
rect 259779 337365 259791 337368
rect 259733 337359 259791 337365
rect 266722 337356 266728 337368
rect 266780 337356 266786 337408
rect 269022 337356 269028 337408
rect 269080 337396 269086 337408
rect 334713 337399 334771 337405
rect 334713 337396 334725 337399
rect 269080 337368 334725 337396
rect 269080 337356 269086 337368
rect 334713 337365 334725 337368
rect 334759 337365 334771 337399
rect 334713 337359 334771 337365
rect 335909 337399 335967 337405
rect 335909 337365 335921 337399
rect 335955 337396 335967 337399
rect 336108 337396 336136 337436
rect 344094 337424 344100 337436
rect 344152 337424 344158 337476
rect 347498 337464 347504 337476
rect 344204 337436 347504 337464
rect 335955 337368 336136 337396
rect 336185 337399 336243 337405
rect 335955 337365 335967 337368
rect 335909 337359 335967 337365
rect 336185 337365 336197 337399
rect 336231 337396 336243 337399
rect 340785 337399 340843 337405
rect 340785 337396 340797 337399
rect 336231 337368 340797 337396
rect 336231 337365 336243 337368
rect 336185 337359 336243 337365
rect 340785 337365 340797 337368
rect 340831 337365 340843 337399
rect 340785 337359 340843 337365
rect 340877 337399 340935 337405
rect 340877 337365 340889 337399
rect 340923 337396 340935 337399
rect 344204 337396 344232 337436
rect 347498 337424 347504 337436
rect 347556 337424 347562 337476
rect 349062 337424 349068 337476
rect 349120 337464 349126 337476
rect 365349 337467 365407 337473
rect 349120 337436 365024 337464
rect 349120 337424 349126 337436
rect 340923 337368 344232 337396
rect 345569 337399 345627 337405
rect 340923 337365 340935 337368
rect 340877 337359 340935 337365
rect 345569 337365 345581 337399
rect 345615 337396 345627 337399
rect 354033 337399 354091 337405
rect 354033 337396 354045 337399
rect 345615 337368 354045 337396
rect 345615 337365 345627 337368
rect 345569 337359 345627 337365
rect 354033 337365 354045 337368
rect 354079 337365 354091 337399
rect 354033 337359 354091 337365
rect 79318 337288 79324 337340
rect 79376 337328 79382 337340
rect 260834 337328 260840 337340
rect 79376 337300 260840 337328
rect 79376 337288 79382 337300
rect 260834 337288 260840 337300
rect 260892 337288 260898 337340
rect 272794 337288 272800 337340
rect 272852 337328 272858 337340
rect 272852 337300 306236 337328
rect 272852 337288 272858 337300
rect 84838 337220 84844 337272
rect 84896 337260 84902 337272
rect 263778 337260 263784 337272
rect 84896 337232 263784 337260
rect 84896 337220 84902 337232
rect 263778 337220 263784 337232
rect 263836 337220 263842 337272
rect 271322 337220 271328 337272
rect 271380 337260 271386 337272
rect 271380 337232 306144 337260
rect 271380 337220 271386 337232
rect 77938 337152 77944 337204
rect 77996 337192 78002 337204
rect 115569 337195 115627 337201
rect 115569 337192 115581 337195
rect 77996 337164 115581 337192
rect 77996 337152 78002 337164
rect 115569 337161 115581 337164
rect 115615 337161 115627 337195
rect 115569 337155 115627 337161
rect 115845 337195 115903 337201
rect 115845 337161 115857 337195
rect 115891 337192 115903 337195
rect 257890 337192 257896 337204
rect 115891 337164 257896 337192
rect 115891 337161 115903 337164
rect 115845 337155 115903 337161
rect 257890 337152 257896 337164
rect 257948 337152 257954 337204
rect 297910 337152 297916 337204
rect 297968 337192 297974 337204
rect 303985 337195 304043 337201
rect 303985 337192 303997 337195
rect 297968 337164 303997 337192
rect 297968 337152 297974 337164
rect 303985 337161 303997 337164
rect 304031 337161 304043 337195
rect 303985 337155 304043 337161
rect 100662 337084 100668 337136
rect 100720 337124 100726 337136
rect 115477 337127 115535 337133
rect 115477 337124 115489 337127
rect 100720 337096 115489 337124
rect 100720 337084 100726 337096
rect 115477 337093 115489 337096
rect 115523 337093 115535 337127
rect 115477 337087 115535 337093
rect 115753 337127 115811 337133
rect 115753 337093 115765 337127
rect 115799 337124 115811 337127
rect 134797 337127 134855 337133
rect 134797 337124 134809 337127
rect 115799 337096 134809 337124
rect 115799 337093 115811 337096
rect 115753 337087 115811 337093
rect 134797 337093 134809 337096
rect 134843 337093 134855 337127
rect 134797 337087 134855 337093
rect 135073 337127 135131 337133
rect 135073 337093 135085 337127
rect 135119 337124 135131 337127
rect 154117 337127 154175 337133
rect 154117 337124 154129 337127
rect 135119 337096 154129 337124
rect 135119 337093 135131 337096
rect 135073 337087 135131 337093
rect 154117 337093 154129 337096
rect 154163 337093 154175 337127
rect 154117 337087 154175 337093
rect 154301 337127 154359 337133
rect 154301 337093 154313 337127
rect 154347 337124 154359 337127
rect 173437 337127 173495 337133
rect 173437 337124 173449 337127
rect 154347 337096 173449 337124
rect 154347 337093 154359 337096
rect 154301 337087 154359 337093
rect 173437 337093 173449 337096
rect 173483 337093 173495 337127
rect 173437 337087 173495 337093
rect 173621 337127 173679 337133
rect 173621 337093 173633 337127
rect 173667 337124 173679 337127
rect 192757 337127 192815 337133
rect 192757 337124 192769 337127
rect 173667 337096 192769 337124
rect 173667 337093 173679 337096
rect 173621 337087 173679 337093
rect 192757 337093 192769 337096
rect 192803 337093 192815 337127
rect 192757 337087 192815 337093
rect 192941 337127 192999 337133
rect 192941 337093 192953 337127
rect 192987 337124 192999 337127
rect 212077 337127 212135 337133
rect 212077 337124 212089 337127
rect 192987 337096 212089 337124
rect 192987 337093 192999 337096
rect 192941 337087 192999 337093
rect 212077 337093 212089 337096
rect 212123 337093 212135 337127
rect 212077 337087 212135 337093
rect 212261 337127 212319 337133
rect 212261 337093 212273 337127
rect 212307 337124 212319 337127
rect 271138 337124 271144 337136
rect 212307 337096 271144 337124
rect 212307 337093 212319 337096
rect 212261 337087 212319 337093
rect 271138 337084 271144 337096
rect 271196 337084 271202 337136
rect 306116 337124 306144 337232
rect 306208 337192 306236 337300
rect 309778 337288 309784 337340
rect 309836 337328 309842 337340
rect 315485 337331 315543 337337
rect 315485 337328 315497 337331
rect 309836 337300 315497 337328
rect 309836 337288 309842 337300
rect 315485 337297 315497 337300
rect 315531 337297 315543 337331
rect 315485 337291 315543 337297
rect 316034 337288 316040 337340
rect 316092 337328 316098 337340
rect 316862 337328 316868 337340
rect 316092 337300 316868 337328
rect 316092 337288 316098 337300
rect 316862 337288 316868 337300
rect 316920 337288 316926 337340
rect 317414 337288 317420 337340
rect 317472 337328 317478 337340
rect 318334 337328 318340 337340
rect 317472 337300 318340 337328
rect 317472 337288 317478 337300
rect 318334 337288 318340 337300
rect 318392 337288 318398 337340
rect 318886 337288 318892 337340
rect 318944 337328 318950 337340
rect 319254 337328 319260 337340
rect 318944 337300 319260 337328
rect 318944 337288 318950 337300
rect 319254 337288 319260 337300
rect 319312 337288 319318 337340
rect 320174 337288 320180 337340
rect 320232 337328 320238 337340
rect 320726 337328 320732 337340
rect 320232 337300 320732 337328
rect 320232 337288 320238 337300
rect 320726 337288 320732 337300
rect 320784 337288 320790 337340
rect 326341 337331 326399 337337
rect 326341 337297 326353 337331
rect 326387 337328 326399 337331
rect 361758 337328 361764 337340
rect 326387 337300 361764 337328
rect 326387 337297 326399 337300
rect 326341 337291 326399 337297
rect 361758 337288 361764 337300
rect 361816 337288 361822 337340
rect 312538 337220 312544 337272
rect 312596 337260 312602 337272
rect 341705 337263 341763 337269
rect 341705 337260 341717 337263
rect 312596 337232 341717 337260
rect 312596 337220 312602 337232
rect 341705 337229 341717 337232
rect 341751 337229 341763 337263
rect 341705 337223 341763 337229
rect 341794 337220 341800 337272
rect 341852 337260 341858 337272
rect 348970 337260 348976 337272
rect 341852 337232 348976 337260
rect 341852 337220 341858 337232
rect 348970 337220 348976 337232
rect 349028 337220 349034 337272
rect 359458 337220 359464 337272
rect 359516 337260 359522 337272
rect 363690 337260 363696 337272
rect 359516 337232 363696 337260
rect 359516 337220 359522 337232
rect 363690 337220 363696 337232
rect 363748 337220 363754 337272
rect 364996 337260 365024 337436
rect 365349 337433 365361 337467
rect 365395 337464 365407 337467
rect 372062 337464 372068 337476
rect 365395 337436 372068 337464
rect 365395 337433 365407 337436
rect 365349 337427 365407 337433
rect 372062 337424 372068 337436
rect 372120 337424 372126 337476
rect 374549 337467 374607 337473
rect 374549 337433 374561 337467
rect 374595 337464 374607 337467
rect 381814 337464 381820 337476
rect 374595 337436 381820 337464
rect 374595 337433 374607 337436
rect 374549 337427 374607 337433
rect 381814 337424 381820 337436
rect 381872 337424 381878 337476
rect 396994 337424 397000 337476
rect 397052 337464 397058 337476
rect 405918 337464 405924 337476
rect 397052 337436 405924 337464
rect 397052 337424 397058 337436
rect 405918 337424 405924 337436
rect 405976 337424 405982 337476
rect 420546 337424 420552 337476
rect 420604 337464 420610 337476
rect 426544 337464 426572 337504
rect 432509 337501 432521 337504
rect 432555 337501 432567 337535
rect 432708 337532 432736 337572
rect 436646 337560 436652 337612
rect 436704 337600 436710 337612
rect 437382 337600 437388 337612
rect 436704 337572 437388 337600
rect 436704 337560 436710 337572
rect 437382 337560 437388 337572
rect 437440 337560 437446 337612
rect 437661 337535 437719 337541
rect 432708 337504 437612 337532
rect 432509 337495 432567 337501
rect 420604 337436 426572 337464
rect 420604 337424 420610 337436
rect 432782 337424 432788 337476
rect 432840 337464 432846 337476
rect 436097 337467 436155 337473
rect 436097 337464 436109 337467
rect 432840 337436 436109 337464
rect 432840 337424 432846 337436
rect 436097 337433 436109 337436
rect 436143 337433 436155 337467
rect 436097 337427 436155 337433
rect 437198 337424 437204 337476
rect 437256 337464 437262 337476
rect 437474 337464 437480 337476
rect 437256 337436 437480 337464
rect 437256 337424 437262 337436
rect 437474 337424 437480 337436
rect 437532 337424 437538 337476
rect 437584 337464 437612 337504
rect 437661 337501 437673 337535
rect 437707 337532 437719 337535
rect 439590 337532 439596 337544
rect 437707 337504 439596 337532
rect 437707 337501 437719 337504
rect 437661 337495 437719 337501
rect 439590 337492 439596 337504
rect 439648 337492 439654 337544
rect 442258 337464 442264 337476
rect 437584 337436 442264 337464
rect 442258 337424 442264 337436
rect 442316 337424 442322 337476
rect 442460 337464 442488 337640
rect 449437 337637 449449 337671
rect 449483 337668 449495 337671
rect 455598 337668 455604 337680
rect 449483 337640 455604 337668
rect 449483 337637 449495 337640
rect 449437 337631 449495 337637
rect 455598 337628 455604 337640
rect 455656 337628 455662 337680
rect 457714 337628 457720 337680
rect 457772 337668 457778 337680
rect 461397 337671 461455 337677
rect 461397 337668 461409 337671
rect 457772 337640 461409 337668
rect 457772 337628 457778 337640
rect 461397 337637 461409 337640
rect 461443 337637 461455 337671
rect 461397 337631 461455 337637
rect 461489 337671 461547 337677
rect 461489 337637 461501 337671
rect 461535 337668 461547 337671
rect 483109 337671 483167 337677
rect 483109 337668 483121 337671
rect 461535 337640 483121 337668
rect 461535 337637 461547 337640
rect 461489 337631 461547 337637
rect 483109 337637 483121 337640
rect 483155 337637 483167 337671
rect 483109 337631 483167 337637
rect 483293 337671 483351 337677
rect 483293 337637 483305 337671
rect 483339 337668 483351 337671
rect 521010 337668 521016 337680
rect 483339 337640 521016 337668
rect 483339 337637 483351 337640
rect 483293 337631 483351 337637
rect 521010 337628 521016 337640
rect 521068 337628 521074 337680
rect 443086 337560 443092 337612
rect 443144 337600 443150 337612
rect 444377 337603 444435 337609
rect 444377 337600 444389 337603
rect 443144 337572 444389 337600
rect 443144 337560 443150 337572
rect 444377 337569 444389 337572
rect 444423 337569 444435 337603
rect 444377 337563 444435 337569
rect 448974 337560 448980 337612
rect 449032 337600 449038 337612
rect 483014 337600 483020 337612
rect 449032 337572 483020 337600
rect 449032 337560 449038 337572
rect 483014 337560 483020 337572
rect 483072 337560 483078 337612
rect 483474 337560 483480 337612
rect 483532 337600 483538 337612
rect 518158 337600 518164 337612
rect 483532 337572 518164 337600
rect 483532 337560 483538 337572
rect 518158 337560 518164 337572
rect 518216 337560 518222 337612
rect 463602 337492 463608 337544
rect 463660 337532 463666 337544
rect 483106 337532 483112 337544
rect 463660 337504 483112 337532
rect 463660 337492 463666 337504
rect 483106 337492 483112 337504
rect 483164 337492 483170 337544
rect 483290 337492 483296 337544
rect 483348 337532 483354 337544
rect 514018 337532 514024 337544
rect 483348 337504 514024 337532
rect 483348 337492 483354 337504
rect 514018 337492 514024 337504
rect 514076 337492 514082 337544
rect 449158 337464 449164 337476
rect 442460 337436 449164 337464
rect 449158 337424 449164 337436
rect 449216 337424 449222 337476
rect 451921 337467 451979 337473
rect 451921 337433 451933 337467
rect 451967 337464 451979 337467
rect 483017 337467 483075 337473
rect 483017 337464 483029 337467
rect 451967 337436 483029 337464
rect 451967 337433 451979 337436
rect 451921 337427 451979 337433
rect 483017 337433 483029 337436
rect 483063 337433 483075 337467
rect 483017 337427 483075 337433
rect 483201 337467 483259 337473
rect 483201 337433 483213 337467
rect 483247 337464 483259 337467
rect 516778 337464 516784 337476
rect 483247 337436 516784 337464
rect 483247 337433 483259 337436
rect 483201 337427 483259 337433
rect 516778 337424 516784 337436
rect 516836 337424 516842 337476
rect 369762 337356 369768 337408
rect 369820 337396 369826 337408
rect 369857 337399 369915 337405
rect 369857 337396 369869 337399
rect 369820 337368 369869 337396
rect 369820 337356 369826 337368
rect 369857 337365 369869 337368
rect 369903 337365 369915 337399
rect 369857 337359 369915 337365
rect 400950 337356 400956 337408
rect 401008 337396 401014 337408
rect 402238 337396 402244 337408
rect 401008 337368 402244 337396
rect 401008 337356 401014 337368
rect 402238 337356 402244 337368
rect 402296 337356 402302 337408
rect 408770 337396 408776 337408
rect 402808 337368 408776 337396
rect 367002 337288 367008 337340
rect 367060 337328 367066 337340
rect 380802 337328 380808 337340
rect 367060 337300 380808 337328
rect 367060 337288 367066 337300
rect 380802 337288 380808 337300
rect 380860 337288 380866 337340
rect 398466 337288 398472 337340
rect 398524 337328 398530 337340
rect 402808 337328 402836 337368
rect 408770 337356 408776 337368
rect 408828 337356 408834 337408
rect 409138 337356 409144 337408
rect 409196 337396 409202 337408
rect 409196 337368 412680 337396
rect 409196 337356 409202 337368
rect 398524 337300 402836 337328
rect 398524 337288 398530 337300
rect 372982 337260 372988 337272
rect 364996 337232 372988 337260
rect 372982 337220 372988 337232
rect 373040 337220 373046 337272
rect 412652 337260 412680 337368
rect 412726 337356 412732 337408
rect 412784 337396 412790 337408
rect 413830 337396 413836 337408
rect 412784 337368 413836 337396
rect 412784 337356 412790 337368
rect 413830 337356 413836 337368
rect 413888 337356 413894 337408
rect 414109 337399 414167 337405
rect 414109 337365 414121 337399
rect 414155 337396 414167 337399
rect 421190 337396 421196 337408
rect 414155 337368 421196 337396
rect 414155 337365 414167 337368
rect 414109 337359 414167 337365
rect 421190 337356 421196 337368
rect 421248 337356 421254 337408
rect 432601 337399 432659 337405
rect 432601 337365 432613 337399
rect 432647 337396 432659 337399
rect 438118 337396 438124 337408
rect 432647 337368 438124 337396
rect 432647 337365 432659 337368
rect 432601 337359 432659 337365
rect 438118 337356 438124 337368
rect 438176 337356 438182 337408
rect 440142 337356 440148 337408
rect 440200 337396 440206 337408
rect 445757 337399 445815 337405
rect 445757 337396 445769 337399
rect 440200 337368 445769 337396
rect 440200 337356 440206 337368
rect 445757 337365 445769 337368
rect 445803 337365 445815 337399
rect 445757 337359 445815 337365
rect 450357 337399 450415 337405
rect 450357 337365 450369 337399
rect 450403 337396 450415 337399
rect 510614 337396 510620 337408
rect 450403 337368 510620 337396
rect 450403 337365 450415 337368
rect 450357 337359 450415 337365
rect 510614 337356 510620 337368
rect 510672 337356 510678 337408
rect 421006 337288 421012 337340
rect 421064 337328 421070 337340
rect 459005 337331 459063 337337
rect 459005 337328 459017 337331
rect 421064 337300 459017 337328
rect 421064 337288 421070 337300
rect 459005 337297 459017 337300
rect 459051 337297 459063 337331
rect 461397 337331 461455 337337
rect 459005 337291 459063 337297
rect 459112 337300 460428 337328
rect 423033 337263 423091 337269
rect 423033 337260 423045 337263
rect 412652 337232 423045 337260
rect 423033 337229 423045 337232
rect 423079 337229 423091 337263
rect 423033 337223 423091 337229
rect 423490 337220 423496 337272
rect 423548 337260 423554 337272
rect 459112 337260 459140 337300
rect 423548 337232 459140 337260
rect 423548 337220 423554 337232
rect 459186 337220 459192 337272
rect 459244 337260 459250 337272
rect 460290 337260 460296 337272
rect 459244 337232 460296 337260
rect 459244 337220 459250 337232
rect 460290 337220 460296 337232
rect 460348 337220 460354 337272
rect 460400 337260 460428 337300
rect 461397 337297 461409 337331
rect 461443 337328 461455 337331
rect 463697 337331 463755 337337
rect 463697 337328 463709 337331
rect 461443 337300 463709 337328
rect 461443 337297 461455 337300
rect 461397 337291 461455 337297
rect 463697 337297 463709 337300
rect 463743 337297 463755 337331
rect 463697 337291 463755 337297
rect 464614 337288 464620 337340
rect 464672 337328 464678 337340
rect 466181 337331 466239 337337
rect 466181 337328 466193 337331
rect 464672 337300 466193 337328
rect 464672 337288 464678 337300
rect 466181 337297 466193 337300
rect 466227 337297 466239 337331
rect 466181 337291 466239 337297
rect 466365 337331 466423 337337
rect 466365 337297 466377 337331
rect 466411 337297 466423 337331
rect 466365 337291 466423 337297
rect 466273 337263 466331 337269
rect 466273 337260 466285 337263
rect 460400 337232 466285 337260
rect 466273 337229 466285 337232
rect 466319 337229 466331 337263
rect 466380 337260 466408 337291
rect 466546 337288 466552 337340
rect 466604 337328 466610 337340
rect 529198 337328 529204 337340
rect 466604 337300 529204 337328
rect 466604 337288 466610 337300
rect 529198 337288 529204 337300
rect 529256 337288 529262 337340
rect 469217 337263 469275 337269
rect 469217 337260 469229 337263
rect 466380 337232 469229 337260
rect 466273 337223 466331 337229
rect 469217 337229 469229 337232
rect 469263 337229 469275 337263
rect 469217 337223 469275 337229
rect 469490 337220 469496 337272
rect 469548 337260 469554 337272
rect 530578 337260 530584 337272
rect 469548 337232 530584 337260
rect 469548 337220 469554 337232
rect 530578 337220 530584 337232
rect 530636 337220 530642 337272
rect 314194 337192 314200 337204
rect 306208 337164 314200 337192
rect 314194 337152 314200 337164
rect 314252 337152 314258 337204
rect 321462 337152 321468 337204
rect 321520 337192 321526 337204
rect 326341 337195 326399 337201
rect 326341 337192 326353 337195
rect 321520 337164 326353 337192
rect 321520 337152 321526 337164
rect 326341 337161 326353 337164
rect 326387 337161 326399 337195
rect 342809 337195 342867 337201
rect 342809 337192 342821 337195
rect 326341 337155 326399 337161
rect 326448 337164 342821 337192
rect 312722 337124 312728 337136
rect 306116 337096 312728 337124
rect 312722 337084 312728 337096
rect 312780 337084 312786 337136
rect 316678 337084 316684 337136
rect 316736 337124 316742 337136
rect 326448 337124 326476 337164
rect 342809 337161 342821 337164
rect 342855 337161 342867 337195
rect 342809 337155 342867 337161
rect 342898 337152 342904 337204
rect 342956 337192 342962 337204
rect 345845 337195 345903 337201
rect 345845 337192 345857 337195
rect 342956 337164 345857 337192
rect 342956 337152 342962 337164
rect 345845 337161 345857 337164
rect 345891 337161 345903 337195
rect 345845 337155 345903 337161
rect 355962 337152 355968 337204
rect 356020 337192 356026 337204
rect 364981 337195 365039 337201
rect 364981 337192 364993 337195
rect 356020 337164 364993 337192
rect 356020 337152 356026 337164
rect 364981 337161 364993 337164
rect 365027 337161 365039 337195
rect 364981 337155 365039 337161
rect 369857 337195 369915 337201
rect 369857 337161 369869 337195
rect 369903 337192 369915 337195
rect 374549 337195 374607 337201
rect 374549 337192 374561 337195
rect 369903 337164 374561 337192
rect 369903 337161 369915 337164
rect 369857 337155 369915 337161
rect 374549 337161 374561 337164
rect 374595 337161 374607 337195
rect 385218 337192 385224 337204
rect 374549 337155 374607 337161
rect 380728 337164 385224 337192
rect 316736 337096 326476 337124
rect 316736 337084 316742 337096
rect 335262 337084 335268 337136
rect 335320 337124 335326 337136
rect 340785 337127 340843 337133
rect 335320 337096 340736 337124
rect 335320 337084 335326 337096
rect 95878 337016 95884 337068
rect 95936 337056 95942 337068
rect 134705 337059 134763 337065
rect 134705 337056 134717 337059
rect 95936 337028 134717 337056
rect 95936 337016 95942 337028
rect 134705 337025 134717 337028
rect 134751 337025 134763 337059
rect 134705 337019 134763 337025
rect 134981 337059 135039 337065
rect 134981 337025 134993 337059
rect 135027 337056 135039 337059
rect 154025 337059 154083 337065
rect 154025 337056 154037 337059
rect 135027 337028 154037 337056
rect 135027 337025 135039 337028
rect 134981 337019 135039 337025
rect 154025 337025 154037 337028
rect 154071 337025 154083 337059
rect 154025 337019 154083 337025
rect 154393 337059 154451 337065
rect 154393 337025 154405 337059
rect 154439 337056 154451 337059
rect 173345 337059 173403 337065
rect 173345 337056 173357 337059
rect 154439 337028 173357 337056
rect 154439 337025 154451 337028
rect 154393 337019 154451 337025
rect 173345 337025 173357 337028
rect 173391 337025 173403 337059
rect 173345 337019 173403 337025
rect 173713 337059 173771 337065
rect 173713 337025 173725 337059
rect 173759 337056 173771 337059
rect 192665 337059 192723 337065
rect 192665 337056 192677 337059
rect 173759 337028 192677 337056
rect 173759 337025 173771 337028
rect 173713 337019 173771 337025
rect 192665 337025 192677 337028
rect 192711 337025 192723 337059
rect 192665 337019 192723 337025
rect 193033 337059 193091 337065
rect 193033 337025 193045 337059
rect 193079 337056 193091 337059
rect 211985 337059 212043 337065
rect 211985 337056 211997 337059
rect 193079 337028 211997 337056
rect 193079 337025 193091 337028
rect 193033 337019 193091 337025
rect 211985 337025 211997 337028
rect 212031 337025 212043 337059
rect 211985 337019 212043 337025
rect 212353 337059 212411 337065
rect 212353 337025 212365 337059
rect 212399 337056 212411 337059
rect 265250 337056 265256 337068
rect 212399 337028 265256 337056
rect 212399 337025 212411 337028
rect 212353 337019 212411 337025
rect 265250 337016 265256 337028
rect 265308 337016 265314 337068
rect 335817 337059 335875 337065
rect 335817 337025 335829 337059
rect 335863 337056 335875 337059
rect 340601 337059 340659 337065
rect 340601 337056 340613 337059
rect 335863 337028 340613 337056
rect 335863 337025 335875 337028
rect 335817 337019 335875 337025
rect 340601 337025 340613 337028
rect 340647 337025 340659 337059
rect 340708 337056 340736 337096
rect 340785 337093 340797 337127
rect 340831 337124 340843 337127
rect 366634 337124 366640 337136
rect 340831 337096 366640 337124
rect 340831 337093 340843 337096
rect 340785 337087 340843 337093
rect 366634 337084 366640 337096
rect 366692 337084 366698 337136
rect 369118 337084 369124 337136
rect 369176 337124 369182 337136
rect 371050 337124 371056 337136
rect 369176 337096 371056 337124
rect 369176 337084 369182 337096
rect 371050 337084 371056 337096
rect 371108 337084 371114 337136
rect 367646 337056 367652 337068
rect 340708 337028 367652 337056
rect 340601 337019 340659 337025
rect 367646 337016 367652 337028
rect 367704 337016 367710 337068
rect 107562 336948 107568 337000
rect 107620 336988 107626 337000
rect 274082 336988 274088 337000
rect 107620 336960 274088 336988
rect 107620 336948 107626 336960
rect 274082 336948 274088 336960
rect 274140 336948 274146 337000
rect 319438 336948 319444 337000
rect 319496 336988 319502 337000
rect 345845 336991 345903 336997
rect 319496 336960 345704 336988
rect 319496 336948 319502 336960
rect 102778 336880 102784 336932
rect 102836 336920 102842 336932
rect 268194 336920 268200 336932
rect 102836 336892 268200 336920
rect 102836 336880 102842 336892
rect 268194 336880 268200 336892
rect 268252 336880 268258 336932
rect 333238 336880 333244 336932
rect 333296 336920 333302 336932
rect 336185 336923 336243 336929
rect 336185 336920 336197 336923
rect 333296 336892 336197 336920
rect 333296 336880 333302 336892
rect 336185 336889 336197 336892
rect 336231 336889 336243 336923
rect 336185 336883 336243 336889
rect 338758 336880 338764 336932
rect 338816 336920 338822 336932
rect 338816 336892 340736 336920
rect 338816 336880 338822 336892
rect 118602 336812 118608 336864
rect 118660 336852 118666 336864
rect 278498 336852 278504 336864
rect 118660 336824 278504 336852
rect 118660 336812 118666 336824
rect 278498 336812 278504 336824
rect 278556 336812 278562 336864
rect 327718 336812 327724 336864
rect 327776 336852 327782 336864
rect 340708 336852 340736 336892
rect 340782 336880 340788 336932
rect 340840 336920 340846 336932
rect 345569 336923 345627 336929
rect 345569 336920 345581 336923
rect 340840 336892 345581 336920
rect 340840 336880 340846 336892
rect 345569 336889 345581 336892
rect 345615 336889 345627 336923
rect 345569 336883 345627 336889
rect 340877 336855 340935 336861
rect 340877 336852 340889 336855
rect 327776 336824 340552 336852
rect 340708 336824 340889 336852
rect 327776 336812 327782 336824
rect 125502 336744 125508 336796
rect 125560 336784 125566 336796
rect 281166 336784 281172 336796
rect 125560 336756 281172 336784
rect 125560 336744 125566 336756
rect 281166 336744 281172 336756
rect 281224 336744 281230 336796
rect 334713 336787 334771 336793
rect 334713 336753 334725 336787
rect 334759 336784 334771 336787
rect 340230 336784 340236 336796
rect 334759 336756 340236 336784
rect 334759 336753 334771 336756
rect 334713 336747 334771 336753
rect 340230 336744 340236 336756
rect 340288 336744 340294 336796
rect 251818 336676 251824 336728
rect 251876 336716 251882 336728
rect 256418 336716 256424 336728
rect 251876 336688 256424 336716
rect 251876 336676 251882 336688
rect 256418 336676 256424 336688
rect 256476 336676 256482 336728
rect 262858 336676 262864 336728
rect 262916 336716 262922 336728
rect 263042 336716 263048 336728
rect 262916 336688 263048 336716
rect 262916 336676 262922 336688
rect 263042 336676 263048 336688
rect 263100 336676 263106 336728
rect 284386 336716 284392 336728
rect 284347 336688 284392 336716
rect 284386 336676 284392 336688
rect 284444 336676 284450 336728
rect 288805 336719 288863 336725
rect 288805 336685 288817 336719
rect 288851 336716 288863 336719
rect 288986 336716 288992 336728
rect 288851 336688 288992 336716
rect 288851 336685 288863 336688
rect 288805 336679 288863 336685
rect 288986 336676 288992 336688
rect 289044 336676 289050 336728
rect 327261 336719 327319 336725
rect 327261 336685 327273 336719
rect 327307 336716 327319 336719
rect 327626 336716 327632 336728
rect 327307 336688 327632 336716
rect 327307 336685 327319 336688
rect 327261 336679 327319 336685
rect 327626 336676 327632 336688
rect 327684 336676 327690 336728
rect 339773 336719 339831 336725
rect 339773 336685 339785 336719
rect 339819 336716 339831 336719
rect 340322 336716 340328 336728
rect 339819 336688 340328 336716
rect 339819 336685 339831 336688
rect 339773 336679 339831 336685
rect 340322 336676 340328 336688
rect 340380 336676 340386 336728
rect 340524 336580 340552 336824
rect 340877 336821 340889 336824
rect 340923 336821 340935 336855
rect 340877 336815 340935 336821
rect 341076 336824 343220 336852
rect 340785 336787 340843 336793
rect 340785 336753 340797 336787
rect 340831 336784 340843 336787
rect 340969 336787 341027 336793
rect 340969 336784 340981 336787
rect 340831 336756 340981 336784
rect 340831 336753 340843 336756
rect 340785 336747 340843 336753
rect 340969 336753 340981 336756
rect 341015 336753 341027 336787
rect 340969 336747 341027 336753
rect 341076 336580 341104 336824
rect 341153 336787 341211 336793
rect 341153 336753 341165 336787
rect 341199 336784 341211 336787
rect 343082 336784 343088 336796
rect 341199 336756 343088 336784
rect 341199 336753 341211 336756
rect 341153 336747 341211 336753
rect 343082 336744 343088 336756
rect 343140 336744 343146 336796
rect 343192 336784 343220 336824
rect 344278 336812 344284 336864
rect 344336 336852 344342 336864
rect 345477 336855 345535 336861
rect 345477 336852 345489 336855
rect 344336 336824 345489 336852
rect 344336 336812 344342 336824
rect 345477 336821 345489 336824
rect 345523 336821 345535 336855
rect 345477 336815 345535 336821
rect 345566 336784 345572 336796
rect 343192 336756 345572 336784
rect 345566 336744 345572 336756
rect 345624 336744 345630 336796
rect 345676 336784 345704 336960
rect 345845 336957 345857 336991
rect 345891 336988 345903 336991
rect 353386 336988 353392 337000
rect 345891 336960 353392 336988
rect 345891 336957 345903 336960
rect 345845 336951 345903 336957
rect 353386 336948 353392 336960
rect 353444 336948 353450 337000
rect 354033 336991 354091 336997
rect 354033 336957 354045 336991
rect 354079 336988 354091 336991
rect 354079 336960 364932 336988
rect 354079 336957 354091 336960
rect 354033 336951 354091 336957
rect 345934 336880 345940 336932
rect 345992 336920 345998 336932
rect 360286 336920 360292 336932
rect 345992 336892 360292 336920
rect 345992 336880 345998 336892
rect 360286 336880 360292 336892
rect 360344 336880 360350 336932
rect 364904 336920 364932 336960
rect 366910 336948 366916 337000
rect 366968 336988 366974 337000
rect 374641 336991 374699 336997
rect 374641 336988 374653 336991
rect 366968 336960 374653 336988
rect 366968 336948 366974 336960
rect 374641 336957 374653 336960
rect 374687 336957 374699 336991
rect 374641 336951 374699 336957
rect 378042 336948 378048 337000
rect 378100 336988 378106 337000
rect 380728 336988 380756 337164
rect 385218 337152 385224 337164
rect 385276 337152 385282 337204
rect 401870 337152 401876 337204
rect 401928 337192 401934 337204
rect 416958 337192 416964 337204
rect 401928 337164 416964 337192
rect 401928 337152 401934 337164
rect 416958 337152 416964 337164
rect 417016 337152 417022 337204
rect 431218 337192 431224 337204
rect 422404 337164 431224 337192
rect 380802 337084 380808 337136
rect 380860 337124 380866 337136
rect 386230 337124 386236 337136
rect 380860 337096 386236 337124
rect 380860 337084 380866 337096
rect 386230 337084 386236 337096
rect 386288 337084 386294 337136
rect 415118 337084 415124 337136
rect 415176 337124 415182 337136
rect 421558 337124 421564 337136
rect 415176 337096 421564 337124
rect 415176 337084 415182 337096
rect 421558 337084 421564 337096
rect 421616 337084 421622 337136
rect 407758 337016 407764 337068
rect 407816 337056 407822 337068
rect 409138 337056 409144 337068
rect 407816 337028 409144 337056
rect 407816 337016 407822 337028
rect 409138 337016 409144 337028
rect 409196 337016 409202 337068
rect 419074 337016 419080 337068
rect 419132 337056 419138 337068
rect 422404 337056 422432 337164
rect 431218 337152 431224 337164
rect 431276 337152 431282 337204
rect 431405 337195 431463 337201
rect 431405 337161 431417 337195
rect 431451 337192 431463 337195
rect 433518 337192 433524 337204
rect 431451 337164 433524 337192
rect 431451 337161 431463 337164
rect 431405 337155 431463 337161
rect 433518 337152 433524 337164
rect 433576 337152 433582 337204
rect 434254 337152 434260 337204
rect 434312 337192 434318 337204
rect 437477 337195 437535 337201
rect 437477 337192 437489 337195
rect 434312 337164 437489 337192
rect 434312 337152 434318 337164
rect 437477 337161 437489 337164
rect 437523 337161 437535 337195
rect 437477 337155 437535 337161
rect 437569 337195 437627 337201
rect 437569 337161 437581 337195
rect 437615 337192 437627 337195
rect 492674 337192 492680 337204
rect 437615 337164 492680 337192
rect 437615 337161 437627 337164
rect 437569 337155 437627 337161
rect 492674 337152 492680 337164
rect 492732 337152 492738 337204
rect 429289 337127 429347 337133
rect 429289 337093 429301 337127
rect 429335 337124 429347 337127
rect 433978 337124 433984 337136
rect 429335 337096 433984 337124
rect 429335 337093 429347 337096
rect 429289 337087 429347 337093
rect 433978 337084 433984 337096
rect 434036 337084 434042 337136
rect 434073 337127 434131 337133
rect 434073 337093 434085 337127
rect 434119 337124 434131 337127
rect 485774 337124 485780 337136
rect 434119 337096 485780 337124
rect 434119 337093 434131 337096
rect 434073 337087 434131 337093
rect 485774 337084 485780 337096
rect 485832 337084 485838 337136
rect 419132 337028 422432 337056
rect 419132 337016 419138 337028
rect 422478 337016 422484 337068
rect 422536 337056 422542 337068
rect 424410 337056 424416 337068
rect 422536 337028 424416 337056
rect 422536 337016 422542 337028
rect 424410 337016 424416 337028
rect 424468 337016 424474 337068
rect 431405 337059 431463 337065
rect 431405 337056 431417 337059
rect 427832 337028 431417 337056
rect 378100 336960 380756 336988
rect 378100 336948 378106 336960
rect 382182 336948 382188 337000
rect 382240 336988 382246 337000
rect 386690 336988 386696 337000
rect 382240 336960 386696 336988
rect 382240 336948 382246 336960
rect 386690 336948 386696 336960
rect 386748 336948 386754 337000
rect 401410 336948 401416 337000
rect 401468 336988 401474 337000
rect 404998 336988 405004 337000
rect 401468 336960 405004 336988
rect 401468 336948 401474 336960
rect 404998 336948 405004 336960
rect 405056 336948 405062 337000
rect 409230 336948 409236 337000
rect 409288 336988 409294 337000
rect 423033 336991 423091 336997
rect 409288 336960 422984 336988
rect 409288 336948 409294 336960
rect 369578 336920 369584 336932
rect 364904 336892 369584 336920
rect 369578 336880 369584 336892
rect 369636 336880 369642 336932
rect 384298 336880 384304 336932
rect 384356 336920 384362 336932
rect 387702 336920 387708 336932
rect 384356 336892 387708 336920
rect 384356 336880 384362 336892
rect 387702 336880 387708 336892
rect 387760 336880 387766 336932
rect 345753 336855 345811 336861
rect 345753 336821 345765 336855
rect 345799 336852 345811 336855
rect 357342 336852 357348 336864
rect 345799 336824 357348 336852
rect 345799 336821 345811 336824
rect 345753 336815 345811 336821
rect 357342 336812 357348 336824
rect 357400 336812 357406 336864
rect 362218 336812 362224 336864
rect 362276 336852 362282 336864
rect 365162 336852 365168 336864
rect 362276 336824 365168 336852
rect 362276 336812 362282 336824
rect 365162 336812 365168 336824
rect 365220 336812 365226 336864
rect 381630 336812 381636 336864
rect 381688 336852 381694 336864
rect 384758 336852 384764 336864
rect 381688 336824 384764 336852
rect 381688 336812 381694 336824
rect 384758 336812 384764 336824
rect 384816 336812 384822 336864
rect 384942 336812 384948 336864
rect 385000 336852 385006 336864
rect 388162 336852 388168 336864
rect 385000 336824 388168 336852
rect 385000 336812 385006 336824
rect 388162 336812 388168 336824
rect 388220 336812 388226 336864
rect 419994 336812 420000 336864
rect 420052 336852 420058 336864
rect 420730 336852 420736 336864
rect 420052 336824 420736 336852
rect 420052 336812 420058 336824
rect 420730 336812 420736 336824
rect 420788 336812 420794 336864
rect 351454 336784 351460 336796
rect 345676 336756 351460 336784
rect 351454 336744 351460 336756
rect 351512 336744 351518 336796
rect 352558 336744 352564 336796
rect 352616 336784 352622 336796
rect 357802 336784 357808 336796
rect 352616 336756 357808 336784
rect 352616 336744 352622 336756
rect 357802 336744 357808 336756
rect 357860 336744 357866 336796
rect 363598 336744 363604 336796
rect 363656 336784 363662 336796
rect 364702 336784 364708 336796
rect 363656 336756 364708 336784
rect 363656 336744 363662 336756
rect 364702 336744 364708 336756
rect 364760 336744 364766 336796
rect 370498 336744 370504 336796
rect 370556 336784 370562 336796
rect 372522 336784 372528 336796
rect 370556 336756 372528 336784
rect 370556 336744 370562 336756
rect 372522 336744 372528 336756
rect 372580 336744 372586 336796
rect 376018 336744 376024 336796
rect 376076 336784 376082 336796
rect 376938 336784 376944 336796
rect 376076 336756 376944 336784
rect 376076 336744 376082 336756
rect 376938 336744 376944 336756
rect 376996 336744 377002 336796
rect 377674 336744 377680 336796
rect 377732 336784 377738 336796
rect 378410 336784 378416 336796
rect 377732 336756 378416 336784
rect 377732 336744 377738 336756
rect 378410 336744 378416 336756
rect 378468 336744 378474 336796
rect 380158 336744 380164 336796
rect 380216 336784 380222 336796
rect 381354 336784 381360 336796
rect 380216 336756 381360 336784
rect 380216 336744 380222 336756
rect 381354 336744 381360 336756
rect 381412 336744 381418 336796
rect 381538 336744 381544 336796
rect 381596 336784 381602 336796
rect 382826 336784 382832 336796
rect 381596 336756 382832 336784
rect 381596 336744 381602 336756
rect 382826 336744 382832 336756
rect 382884 336744 382890 336796
rect 387058 336744 387064 336796
rect 387116 336784 387122 336796
rect 388714 336784 388720 336796
rect 387116 336756 388720 336784
rect 387116 336744 387122 336756
rect 388714 336744 388720 336756
rect 388772 336744 388778 336796
rect 392394 336744 392400 336796
rect 392452 336784 392458 336796
rect 393590 336784 393596 336796
rect 392452 336756 393596 336784
rect 392452 336744 392458 336756
rect 393590 336744 393596 336756
rect 393648 336744 393654 336796
rect 418522 336744 418528 336796
rect 418580 336784 418586 336796
rect 419442 336784 419448 336796
rect 418580 336756 419448 336784
rect 418580 336744 418586 336756
rect 419442 336744 419448 336756
rect 419500 336744 419506 336796
rect 419534 336744 419540 336796
rect 419592 336784 419598 336796
rect 420822 336784 420828 336796
rect 419592 336756 420828 336784
rect 419592 336744 419598 336756
rect 420822 336744 420828 336756
rect 420880 336744 420886 336796
rect 421466 336744 421472 336796
rect 421524 336784 421530 336796
rect 422202 336784 422208 336796
rect 421524 336756 422208 336784
rect 421524 336744 421530 336756
rect 422202 336744 422208 336756
rect 422260 336744 422266 336796
rect 422956 336784 422984 336960
rect 423033 336957 423045 336991
rect 423079 336988 423091 336991
rect 427832 336988 427860 337028
rect 431405 337025 431417 337028
rect 431451 337025 431463 337059
rect 477586 337056 477592 337068
rect 431405 337019 431463 337025
rect 432524 337028 477592 337056
rect 423079 336960 427860 336988
rect 423079 336957 423091 336960
rect 423033 336951 423091 336957
rect 428366 336948 428372 337000
rect 428424 336988 428430 337000
rect 431310 336988 431316 337000
rect 428424 336960 431316 336988
rect 428424 336948 428430 336960
rect 431310 336948 431316 336960
rect 431368 336948 431374 337000
rect 423950 336880 423956 336932
rect 424008 336920 424014 336932
rect 432417 336923 432475 336929
rect 432417 336920 432429 336923
rect 424008 336892 432429 336920
rect 424008 336880 424014 336892
rect 432417 336889 432429 336892
rect 432463 336889 432475 336923
rect 432417 336883 432475 336889
rect 426894 336812 426900 336864
rect 426952 336852 426958 336864
rect 432524 336852 432552 337028
rect 477586 337016 477592 337028
rect 477644 337016 477650 337068
rect 432693 336991 432751 336997
rect 432693 336957 432705 336991
rect 432739 336988 432751 336991
rect 475378 336988 475384 337000
rect 432739 336960 475384 336988
rect 432739 336957 432751 336960
rect 432693 336951 432751 336957
rect 475378 336948 475384 336960
rect 475436 336948 475442 337000
rect 466273 336923 466331 336929
rect 466273 336920 466285 336923
rect 432708 336892 466285 336920
rect 426952 336824 432552 336852
rect 432601 336855 432659 336861
rect 426952 336812 426958 336824
rect 432601 336821 432613 336855
rect 432647 336852 432659 336855
rect 432708 336852 432736 336892
rect 466273 336889 466285 336892
rect 466319 336889 466331 336923
rect 466273 336883 466331 336889
rect 466365 336923 466423 336929
rect 466365 336889 466377 336923
rect 466411 336920 466423 336923
rect 469214 336920 469220 336932
rect 466411 336892 469220 336920
rect 466411 336889 466423 336892
rect 466365 336883 466423 336889
rect 469214 336880 469220 336892
rect 469272 336880 469278 336932
rect 469324 336892 470732 336920
rect 432647 336824 432736 336852
rect 432647 336821 432659 336824
rect 432601 336815 432659 336821
rect 434714 336812 434720 336864
rect 434772 336852 434778 336864
rect 436002 336852 436008 336864
rect 434772 336824 436008 336852
rect 434772 336812 434778 336824
rect 436002 336812 436008 336824
rect 436060 336812 436066 336864
rect 436097 336855 436155 336861
rect 436097 336821 436109 336855
rect 436143 336852 436155 336855
rect 437477 336855 437535 336861
rect 437477 336852 437489 336855
rect 436143 336824 437489 336852
rect 436143 336821 436155 336824
rect 436097 336815 436155 336821
rect 437477 336821 437489 336824
rect 437523 336821 437535 336855
rect 439498 336852 439504 336864
rect 437477 336815 437535 336821
rect 437584 336824 439504 336852
rect 429289 336787 429347 336793
rect 429289 336784 429301 336787
rect 422956 336756 429301 336784
rect 429289 336753 429301 336756
rect 429335 336753 429347 336787
rect 429289 336747 429347 336753
rect 429378 336744 429384 336796
rect 429436 336784 429442 336796
rect 430482 336784 430488 336796
rect 429436 336756 430488 336784
rect 429436 336744 429442 336756
rect 430482 336744 430488 336756
rect 430540 336744 430546 336796
rect 430850 336744 430856 336796
rect 430908 336784 430914 336796
rect 431862 336784 431868 336796
rect 430908 336756 431868 336784
rect 430908 336744 430914 336756
rect 431862 336744 431868 336756
rect 431920 336744 431926 336796
rect 432322 336744 432328 336796
rect 432380 336784 432386 336796
rect 433150 336784 433156 336796
rect 432380 336756 433156 336784
rect 432380 336744 432386 336756
rect 433150 336744 433156 336756
rect 433208 336744 433214 336796
rect 433702 336744 433708 336796
rect 433760 336784 433766 336796
rect 434622 336784 434628 336796
rect 433760 336756 434628 336784
rect 433760 336744 433766 336756
rect 434622 336744 434628 336756
rect 434680 336744 434686 336796
rect 435174 336744 435180 336796
rect 435232 336784 435238 336796
rect 435910 336784 435916 336796
rect 435232 336756 435916 336784
rect 435232 336744 435238 336756
rect 435910 336744 435916 336756
rect 435968 336744 435974 336796
rect 436186 336744 436192 336796
rect 436244 336784 436250 336796
rect 437290 336784 437296 336796
rect 436244 336756 437296 336784
rect 436244 336744 436250 336756
rect 437290 336744 437296 336756
rect 437348 336744 437354 336796
rect 437385 336787 437443 336793
rect 437385 336753 437397 336787
rect 437431 336784 437443 336787
rect 437584 336784 437612 336824
rect 439498 336812 439504 336824
rect 439556 336812 439562 336864
rect 441614 336812 441620 336864
rect 441672 336852 441678 336864
rect 443638 336852 443644 336864
rect 441672 336824 443644 336852
rect 441672 336812 441678 336824
rect 443638 336812 443644 336824
rect 443696 336812 443702 336864
rect 444558 336812 444564 336864
rect 444616 336852 444622 336864
rect 445662 336852 445668 336864
rect 444616 336824 445668 336852
rect 444616 336812 444622 336824
rect 445662 336812 445668 336824
rect 445720 336812 445726 336864
rect 445757 336855 445815 336861
rect 445757 336821 445769 336855
rect 445803 336852 445815 336855
rect 450357 336855 450415 336861
rect 450357 336852 450369 336855
rect 445803 336824 450369 336852
rect 445803 336821 445815 336824
rect 445757 336815 445815 336821
rect 450357 336821 450369 336824
rect 450403 336821 450415 336855
rect 450357 336815 450415 336821
rect 450446 336812 450452 336864
rect 450504 336852 450510 336864
rect 451182 336852 451188 336864
rect 450504 336824 451188 336852
rect 450504 336812 450510 336824
rect 451182 336812 451188 336824
rect 451240 336812 451246 336864
rect 453298 336812 453304 336864
rect 453356 336852 453362 336864
rect 453942 336852 453948 336864
rect 453356 336824 453948 336852
rect 453356 336812 453362 336824
rect 453942 336812 453948 336824
rect 454000 336812 454006 336864
rect 456794 336812 456800 336864
rect 456852 336852 456858 336864
rect 458082 336852 458088 336864
rect 456852 336824 458088 336852
rect 456852 336812 456858 336824
rect 458082 336812 458088 336824
rect 458140 336812 458146 336864
rect 459646 336852 459652 336864
rect 458192 336824 459652 336852
rect 437431 336756 437612 336784
rect 437431 336753 437443 336756
rect 437385 336747 437443 336753
rect 439130 336744 439136 336796
rect 439188 336784 439194 336796
rect 440142 336784 440148 336796
rect 439188 336756 440148 336784
rect 439188 336744 439194 336756
rect 440142 336744 440148 336756
rect 440200 336744 440206 336796
rect 440602 336744 440608 336796
rect 440660 336784 440666 336796
rect 441522 336784 441528 336796
rect 440660 336756 441528 336784
rect 440660 336744 440666 336756
rect 441522 336744 441528 336756
rect 441580 336744 441586 336796
rect 442074 336744 442080 336796
rect 442132 336784 442138 336796
rect 442902 336784 442908 336796
rect 442132 336756 442908 336784
rect 442132 336744 442138 336756
rect 442902 336744 442908 336756
rect 442960 336744 442966 336796
rect 443546 336744 443552 336796
rect 443604 336784 443610 336796
rect 444282 336784 444288 336796
rect 443604 336756 444288 336784
rect 443604 336744 443610 336756
rect 444282 336744 444288 336756
rect 444340 336744 444346 336796
rect 445018 336744 445024 336796
rect 445076 336784 445082 336796
rect 445570 336784 445576 336796
rect 445076 336756 445576 336784
rect 445076 336744 445082 336756
rect 445570 336744 445576 336756
rect 445628 336744 445634 336796
rect 446490 336744 446496 336796
rect 446548 336784 446554 336796
rect 447042 336784 447048 336796
rect 446548 336756 447048 336784
rect 446548 336744 446554 336756
rect 447042 336744 447048 336756
rect 447100 336744 447106 336796
rect 447502 336744 447508 336796
rect 447560 336784 447566 336796
rect 447560 336756 448192 336784
rect 447560 336744 447566 336756
rect 421190 336716 421196 336728
rect 421151 336688 421196 336716
rect 421190 336676 421196 336688
rect 421248 336676 421254 336728
rect 448164 336648 448192 336756
rect 448238 336744 448244 336796
rect 448296 336784 448302 336796
rect 448422 336784 448428 336796
rect 448296 336756 448428 336784
rect 448296 336744 448302 336756
rect 448422 336744 448428 336756
rect 448480 336744 448486 336796
rect 449894 336744 449900 336796
rect 449952 336784 449958 336796
rect 450998 336784 451004 336796
rect 449952 336756 451004 336784
rect 449952 336744 449958 336756
rect 450998 336744 451004 336756
rect 451056 336744 451062 336796
rect 451366 336744 451372 336796
rect 451424 336784 451430 336796
rect 452470 336784 452476 336796
rect 451424 336756 452476 336784
rect 451424 336744 451430 336756
rect 452470 336744 452476 336756
rect 452528 336744 452534 336796
rect 452838 336744 452844 336796
rect 452896 336784 452902 336796
rect 453758 336784 453764 336796
rect 452896 336756 453764 336784
rect 452896 336744 452902 336756
rect 453758 336744 453764 336756
rect 453816 336744 453822 336796
rect 454310 336744 454316 336796
rect 454368 336784 454374 336796
rect 455230 336784 455236 336796
rect 454368 336756 455236 336784
rect 454368 336744 454374 336756
rect 455230 336744 455236 336756
rect 455288 336744 455294 336796
rect 455782 336744 455788 336796
rect 455840 336784 455846 336796
rect 456610 336784 456616 336796
rect 455840 336756 456616 336784
rect 455840 336744 455846 336756
rect 456610 336744 456616 336756
rect 456668 336744 456674 336796
rect 456705 336787 456763 336793
rect 456705 336753 456717 336787
rect 456751 336784 456763 336787
rect 456751 336756 457208 336784
rect 456751 336753 456763 336756
rect 456705 336747 456763 336753
rect 457180 336716 457208 336756
rect 457254 336744 457260 336796
rect 457312 336784 457318 336796
rect 457990 336784 457996 336796
rect 457312 336756 457996 336784
rect 457312 336744 457318 336756
rect 457990 336744 457996 336756
rect 458048 336744 458054 336796
rect 458192 336784 458220 336824
rect 459646 336812 459652 336824
rect 459704 336812 459710 336864
rect 463786 336852 463792 336864
rect 459756 336824 463792 336852
rect 458100 336756 458220 336784
rect 458100 336716 458128 336756
rect 458266 336744 458272 336796
rect 458324 336784 458330 336796
rect 459462 336784 459468 336796
rect 458324 336756 459468 336784
rect 458324 336744 458330 336756
rect 459462 336744 459468 336756
rect 459520 336744 459526 336796
rect 457180 336688 458128 336716
rect 459005 336719 459063 336725
rect 459005 336685 459017 336719
rect 459051 336716 459063 336719
rect 459756 336716 459784 336824
rect 463786 336812 463792 336824
rect 463844 336812 463850 336864
rect 466181 336855 466239 336861
rect 466181 336821 466193 336855
rect 466227 336821 466239 336855
rect 466181 336815 466239 336821
rect 461210 336744 461216 336796
rect 461268 336784 461274 336796
rect 462130 336784 462136 336796
rect 461268 336756 462136 336784
rect 461268 336744 461274 336756
rect 462130 336744 462136 336756
rect 462188 336744 462194 336796
rect 462682 336744 462688 336796
rect 462740 336784 462746 336796
rect 463510 336784 463516 336796
rect 462740 336756 463516 336784
rect 462740 336744 462746 336756
rect 463510 336744 463516 336756
rect 463568 336744 463574 336796
rect 464154 336744 464160 336796
rect 464212 336784 464218 336796
rect 464982 336784 464988 336796
rect 464212 336756 464988 336784
rect 464212 336744 464218 336756
rect 464982 336744 464988 336756
rect 465040 336744 465046 336796
rect 466196 336784 466224 336815
rect 469324 336784 469352 336892
rect 470594 336852 470600 336864
rect 465092 336756 466132 336784
rect 466196 336756 469352 336784
rect 469508 336824 470600 336852
rect 459051 336688 459784 336716
rect 459051 336685 459063 336688
rect 459005 336679 459063 336685
rect 461946 336676 461952 336728
rect 462004 336716 462010 336728
rect 465092 336716 465120 336756
rect 462004 336688 465120 336716
rect 466104 336716 466132 336756
rect 469401 336719 469459 336725
rect 469401 336716 469413 336719
rect 466104 336688 469413 336716
rect 462004 336676 462010 336688
rect 469401 336685 469413 336688
rect 469447 336685 469459 336719
rect 469401 336679 469459 336685
rect 448422 336648 448428 336660
rect 448164 336620 448428 336648
rect 448422 336608 448428 336620
rect 448480 336608 448486 336660
rect 466273 336651 466331 336657
rect 466273 336617 466285 336651
rect 466319 336648 466331 336651
rect 469508 336648 469536 336824
rect 470594 336812 470600 336824
rect 470652 336812 470658 336864
rect 470704 336852 470732 336892
rect 509878 336852 509884 336864
rect 470704 336824 509884 336852
rect 509878 336812 509884 336824
rect 509936 336812 509942 336864
rect 469585 336787 469643 336793
rect 469585 336753 469597 336787
rect 469631 336784 469643 336787
rect 505738 336784 505744 336796
rect 469631 336756 505744 336784
rect 469631 336753 469643 336756
rect 469585 336747 469643 336753
rect 505738 336744 505744 336756
rect 505796 336744 505802 336796
rect 466319 336620 469536 336648
rect 466319 336617 466331 336620
rect 466273 336611 466331 336617
rect 340524 336552 341104 336580
rect 247678 336472 247684 336524
rect 247736 336512 247742 336524
rect 248598 336512 248604 336524
rect 247736 336484 248604 336512
rect 247736 336472 247742 336484
rect 248598 336472 248604 336484
rect 248656 336472 248662 336524
rect 248506 336064 248512 336116
rect 248564 336104 248570 336116
rect 249518 336104 249524 336116
rect 248564 336076 249524 336104
rect 248564 336064 248570 336076
rect 249518 336064 249524 336076
rect 249576 336064 249582 336116
rect 236178 335656 236184 335708
rect 236236 335696 236242 335708
rect 237006 335696 237012 335708
rect 236236 335668 237012 335696
rect 236236 335656 236242 335668
rect 237006 335656 237012 335668
rect 237064 335656 237070 335708
rect 302234 335656 302240 335708
rect 302292 335696 302298 335708
rect 302694 335696 302700 335708
rect 302292 335668 302700 335696
rect 302292 335656 302298 335668
rect 302694 335656 302700 335668
rect 302752 335656 302758 335708
rect 332686 335656 332692 335708
rect 332744 335696 332750 335708
rect 333422 335696 333428 335708
rect 332744 335668 333428 335696
rect 332744 335656 332750 335668
rect 333422 335656 333428 335668
rect 333480 335656 333486 335708
rect 334066 335656 334072 335708
rect 334124 335696 334130 335708
rect 334894 335696 334900 335708
rect 334124 335668 334900 335696
rect 334124 335656 334130 335668
rect 334894 335656 334900 335668
rect 334952 335656 334958 335708
rect 236086 335588 236092 335640
rect 236144 335628 236150 335640
rect 236546 335628 236552 335640
rect 236144 335600 236552 335628
rect 236144 335588 236150 335600
rect 236546 335588 236552 335600
rect 236604 335588 236610 335640
rect 241606 335588 241612 335640
rect 241664 335628 241670 335640
rect 242342 335628 242348 335640
rect 241664 335600 242348 335628
rect 241664 335588 241670 335600
rect 242342 335588 242348 335600
rect 242400 335588 242406 335640
rect 260926 335588 260932 335640
rect 260984 335628 260990 335640
rect 261478 335628 261484 335640
rect 260984 335600 261484 335628
rect 260984 335588 260990 335600
rect 261478 335588 261484 335600
rect 261536 335588 261542 335640
rect 263686 335588 263692 335640
rect 263744 335628 263750 335640
rect 264422 335628 264428 335640
rect 263744 335600 264428 335628
rect 263744 335588 263750 335600
rect 264422 335588 264428 335600
rect 264480 335588 264486 335640
rect 265066 335588 265072 335640
rect 265124 335628 265130 335640
rect 265894 335628 265900 335640
rect 265124 335600 265900 335628
rect 265124 335588 265130 335600
rect 265894 335588 265900 335600
rect 265952 335588 265958 335640
rect 266446 335588 266452 335640
rect 266504 335628 266510 335640
rect 267366 335628 267372 335640
rect 266504 335600 267372 335628
rect 266504 335588 266510 335600
rect 267366 335588 267372 335600
rect 267424 335588 267430 335640
rect 280246 335588 280252 335640
rect 280304 335628 280310 335640
rect 280614 335628 280620 335640
rect 280304 335600 280620 335628
rect 280304 335588 280310 335600
rect 280614 335588 280620 335600
rect 280672 335588 280678 335640
rect 281534 335588 281540 335640
rect 281592 335628 281598 335640
rect 282086 335628 282092 335640
rect 281592 335600 282092 335628
rect 281592 335588 281598 335600
rect 282086 335588 282092 335600
rect 282144 335588 282150 335640
rect 283006 335588 283012 335640
rect 283064 335628 283070 335640
rect 283558 335628 283564 335640
rect 283064 335600 283564 335628
rect 283064 335588 283070 335600
rect 283558 335588 283564 335600
rect 283616 335588 283622 335640
rect 285674 335588 285680 335640
rect 285732 335628 285738 335640
rect 285950 335628 285956 335640
rect 285732 335600 285956 335628
rect 285732 335588 285738 335600
rect 285950 335588 285956 335600
rect 286008 335588 286014 335640
rect 286042 335588 286048 335640
rect 286100 335628 286106 335640
rect 286594 335628 286600 335640
rect 286100 335600 286600 335628
rect 286100 335588 286106 335600
rect 286594 335588 286600 335600
rect 286652 335588 286658 335640
rect 287054 335588 287060 335640
rect 287112 335628 287118 335640
rect 287974 335628 287980 335640
rect 287112 335600 287980 335628
rect 287112 335588 287118 335600
rect 287974 335588 287980 335600
rect 288032 335588 288038 335640
rect 288434 335588 288440 335640
rect 288492 335628 288498 335640
rect 289446 335628 289452 335640
rect 288492 335600 289452 335628
rect 288492 335588 288498 335600
rect 289446 335588 289452 335600
rect 289504 335588 289510 335640
rect 292758 335588 292764 335640
rect 292816 335628 292822 335640
rect 293310 335628 293316 335640
rect 292816 335600 293316 335628
rect 292816 335588 292822 335600
rect 293310 335588 293316 335600
rect 293368 335588 293374 335640
rect 298278 335588 298284 335640
rect 298336 335628 298342 335640
rect 298646 335628 298652 335640
rect 298336 335600 298652 335628
rect 298336 335588 298342 335600
rect 298646 335588 298652 335600
rect 298704 335588 298710 335640
rect 300854 335588 300860 335640
rect 300912 335628 300918 335640
rect 301222 335628 301228 335640
rect 300912 335600 301228 335628
rect 300912 335588 300918 335600
rect 301222 335588 301228 335600
rect 301280 335588 301286 335640
rect 303614 335588 303620 335640
rect 303672 335628 303678 335640
rect 304166 335628 304172 335640
rect 303672 335600 304172 335628
rect 303672 335588 303678 335600
rect 304166 335588 304172 335600
rect 304224 335588 304230 335640
rect 304994 335588 305000 335640
rect 305052 335628 305058 335640
rect 305638 335628 305644 335640
rect 305052 335600 305644 335628
rect 305052 335588 305058 335600
rect 305638 335588 305644 335600
rect 305696 335588 305702 335640
rect 307754 335588 307760 335640
rect 307812 335628 307818 335640
rect 308582 335628 308588 335640
rect 307812 335600 308588 335628
rect 307812 335588 307818 335600
rect 308582 335588 308588 335600
rect 308640 335588 308646 335640
rect 309134 335588 309140 335640
rect 309192 335628 309198 335640
rect 310054 335628 310060 335640
rect 309192 335600 310060 335628
rect 309192 335588 309198 335600
rect 310054 335588 310060 335600
rect 310112 335588 310118 335640
rect 321646 335588 321652 335640
rect 321704 335628 321710 335640
rect 322198 335628 322204 335640
rect 321704 335600 322204 335628
rect 321704 335588 321710 335600
rect 322198 335588 322204 335600
rect 322256 335588 322262 335640
rect 329834 335588 329840 335640
rect 329892 335628 329898 335640
rect 330110 335628 330116 335640
rect 329892 335600 330116 335628
rect 329892 335588 329898 335600
rect 330110 335588 330116 335600
rect 330168 335588 330174 335640
rect 332594 335588 332600 335640
rect 332652 335628 332658 335640
rect 333054 335628 333060 335640
rect 332652 335600 333060 335628
rect 332652 335588 332658 335600
rect 333054 335588 333060 335600
rect 333112 335588 333118 335640
rect 333974 335588 333980 335640
rect 334032 335628 334038 335640
rect 334526 335628 334532 335640
rect 334032 335600 334532 335628
rect 334032 335588 334038 335600
rect 334526 335588 334532 335600
rect 334584 335588 334590 335640
rect 335354 335588 335360 335640
rect 335412 335628 335418 335640
rect 335998 335628 336004 335640
rect 335412 335600 336004 335628
rect 335412 335588 335418 335600
rect 335998 335588 336004 335600
rect 336056 335588 336062 335640
rect 338114 335588 338120 335640
rect 338172 335628 338178 335640
rect 338942 335628 338948 335640
rect 338172 335600 338948 335628
rect 338172 335588 338178 335600
rect 338942 335588 338948 335600
rect 339000 335588 339006 335640
rect 363046 335588 363052 335640
rect 363104 335628 363110 335640
rect 363782 335628 363788 335640
rect 363104 335600 363788 335628
rect 363104 335588 363110 335600
rect 363782 335588 363788 335600
rect 363840 335588 363846 335640
rect 367278 335588 367284 335640
rect 367336 335628 367342 335640
rect 367922 335628 367928 335640
rect 367336 335600 367928 335628
rect 367336 335588 367342 335600
rect 367922 335588 367928 335600
rect 367980 335588 367986 335640
rect 374086 335588 374092 335640
rect 374144 335628 374150 335640
rect 374638 335628 374644 335640
rect 374144 335600 374644 335628
rect 374144 335588 374150 335600
rect 374638 335588 374644 335600
rect 374696 335588 374702 335640
rect 465442 335588 465448 335640
rect 465500 335628 465506 335640
rect 466362 335628 466368 335640
rect 465500 335600 466368 335628
rect 465500 335588 465506 335600
rect 466362 335588 466368 335600
rect 466420 335588 466426 335640
rect 245838 335452 245844 335504
rect 245896 335492 245902 335504
rect 246666 335492 246672 335504
rect 245896 335464 246672 335492
rect 245896 335452 245902 335464
rect 246666 335452 246672 335464
rect 246724 335452 246730 335504
rect 438026 335452 438032 335504
rect 438084 335492 438090 335504
rect 438670 335492 438676 335504
rect 438084 335464 438676 335492
rect 438084 335452 438090 335464
rect 438670 335452 438676 335464
rect 438728 335452 438734 335504
rect 284389 335223 284447 335229
rect 284389 335189 284401 335223
rect 284435 335220 284447 335223
rect 284478 335220 284484 335232
rect 284435 335192 284484 335220
rect 284435 335189 284447 335192
rect 284389 335183 284447 335189
rect 284478 335180 284484 335192
rect 284536 335180 284542 335232
rect 258166 334704 258172 334756
rect 258224 334744 258230 334756
rect 258534 334744 258540 334756
rect 258224 334716 258540 334744
rect 258224 334704 258230 334716
rect 258534 334704 258540 334716
rect 258592 334704 258598 334756
rect 302513 334747 302571 334753
rect 302513 334713 302525 334747
rect 302559 334744 302571 334747
rect 303062 334744 303068 334756
rect 302559 334716 303068 334744
rect 302559 334713 302571 334716
rect 302513 334707 302571 334713
rect 303062 334704 303068 334716
rect 303120 334704 303126 334756
rect 234982 334500 234988 334552
rect 235040 334540 235046 334552
rect 235626 334540 235632 334552
rect 235040 334512 235632 334540
rect 235040 334500 235046 334512
rect 235626 334500 235632 334512
rect 235684 334500 235690 334552
rect 250165 334475 250223 334481
rect 250165 334441 250177 334475
rect 250211 334472 250223 334475
rect 250622 334472 250628 334484
rect 250211 334444 250628 334472
rect 250211 334441 250223 334444
rect 250165 334435 250223 334441
rect 250622 334432 250628 334444
rect 250680 334432 250686 334484
rect 270770 334296 270776 334348
rect 270828 334336 270834 334348
rect 271230 334336 271236 334348
rect 270828 334308 271236 334336
rect 270828 334296 270834 334308
rect 271230 334296 271236 334308
rect 271288 334296 271294 334348
rect 272242 334296 272248 334348
rect 272300 334336 272306 334348
rect 272702 334336 272708 334348
rect 272300 334308 272708 334336
rect 272300 334296 272306 334308
rect 272702 334296 272708 334308
rect 272760 334296 272766 334348
rect 247126 334160 247132 334212
rect 247184 334200 247190 334212
rect 248138 334200 248144 334212
rect 247184 334172 248144 334200
rect 247184 334160 247190 334172
rect 248138 334160 248144 334172
rect 248196 334160 248202 334212
rect 278774 333276 278780 333328
rect 278832 333316 278838 333328
rect 278958 333316 278964 333328
rect 278832 333288 278964 333316
rect 278832 333276 278838 333288
rect 278958 333276 278964 333288
rect 279016 333276 279022 333328
rect 325970 333276 325976 333328
rect 326028 333316 326034 333328
rect 326522 333316 326528 333328
rect 326028 333288 326528 333316
rect 326028 333276 326034 333288
rect 326522 333276 326528 333288
rect 326580 333276 326586 333328
rect 336734 333276 336740 333328
rect 336792 333316 336798 333328
rect 336918 333316 336924 333328
rect 336792 333288 336924 333316
rect 336792 333276 336798 333288
rect 336918 333276 336924 333288
rect 336976 333276 336982 333328
rect 361666 333276 361672 333328
rect 361724 333316 361730 333328
rect 362310 333316 362316 333328
rect 361724 333288 362316 333316
rect 361724 333276 361730 333288
rect 362310 333276 362316 333288
rect 362368 333276 362374 333328
rect 356146 332800 356152 332852
rect 356204 332840 356210 332852
rect 356606 332840 356612 332852
rect 356204 332812 356612 332840
rect 356204 332800 356210 332812
rect 356606 332800 356612 332812
rect 356664 332800 356670 332852
rect 284662 332528 284668 332580
rect 284720 332568 284726 332580
rect 285122 332568 285128 332580
rect 284720 332540 285128 332568
rect 284720 332528 284726 332540
rect 285122 332528 285128 332540
rect 285180 332528 285186 332580
rect 331214 332120 331220 332172
rect 331272 332160 331278 332172
rect 331490 332160 331496 332172
rect 331272 332132 331496 332160
rect 331272 332120 331278 332132
rect 331490 332120 331496 332132
rect 331548 332120 331554 332172
rect 242986 332052 242992 332104
rect 243044 332092 243050 332104
rect 243446 332092 243452 332104
rect 243044 332064 243452 332092
rect 243044 332052 243050 332064
rect 243446 332052 243452 332064
rect 243504 332052 243510 332104
rect 310514 332052 310520 332104
rect 310572 332092 310578 332104
rect 311526 332092 311532 332104
rect 310572 332064 311532 332092
rect 310572 332052 310578 332064
rect 311526 332052 311532 332064
rect 311584 332052 311590 332104
rect 301038 331848 301044 331900
rect 301096 331888 301102 331900
rect 301682 331888 301688 331900
rect 301096 331860 301688 331888
rect 301096 331848 301102 331860
rect 301682 331848 301688 331860
rect 301740 331848 301746 331900
rect 331306 331712 331312 331764
rect 331364 331752 331370 331764
rect 331950 331752 331956 331764
rect 331364 331724 331956 331752
rect 331364 331712 331370 331724
rect 331950 331712 331956 331724
rect 332008 331712 332014 331764
rect 328546 331304 328552 331356
rect 328604 331344 328610 331356
rect 329006 331344 329012 331356
rect 328604 331316 329012 331344
rect 328604 331304 328610 331316
rect 329006 331304 329012 331316
rect 329064 331304 329070 331356
rect 299566 331236 299572 331288
rect 299624 331236 299630 331288
rect 336826 331236 336832 331288
rect 336884 331236 336890 331288
rect 259638 331168 259644 331220
rect 259696 331208 259702 331220
rect 259822 331208 259828 331220
rect 259696 331180 259828 331208
rect 259696 331168 259702 331180
rect 259822 331168 259828 331180
rect 259880 331168 259886 331220
rect 299584 331152 299612 331236
rect 336844 331152 336872 331236
rect 341150 331168 341156 331220
rect 341208 331208 341214 331220
rect 341334 331208 341340 331220
rect 341208 331180 341340 331208
rect 341208 331168 341214 331180
rect 341334 331168 341340 331180
rect 341392 331168 341398 331220
rect 360286 331168 360292 331220
rect 360344 331208 360350 331220
rect 360470 331208 360476 331220
rect 360344 331180 360476 331208
rect 360344 331168 360350 331180
rect 360470 331168 360476 331180
rect 360528 331168 360534 331220
rect 459646 331168 459652 331220
rect 459704 331208 459710 331220
rect 460106 331208 460112 331220
rect 459704 331180 460112 331208
rect 459704 331168 459710 331180
rect 460106 331168 460112 331180
rect 460164 331168 460170 331220
rect 299566 331100 299572 331152
rect 299624 331100 299630 331152
rect 299750 331100 299756 331152
rect 299808 331140 299814 331152
rect 300210 331140 300216 331152
rect 299808 331112 300216 331140
rect 299808 331100 299814 331112
rect 300210 331100 300216 331112
rect 300268 331100 300274 331152
rect 336826 331100 336832 331152
rect 336884 331100 336890 331152
rect 299474 331032 299480 331084
rect 299532 331072 299538 331084
rect 299658 331072 299664 331084
rect 299532 331044 299664 331072
rect 299532 331032 299538 331044
rect 299658 331032 299664 331044
rect 299716 331032 299722 331084
rect 306466 331032 306472 331084
rect 306524 331072 306530 331084
rect 306650 331072 306656 331084
rect 306524 331044 306656 331072
rect 306524 331032 306530 331044
rect 306650 331032 306656 331044
rect 306708 331032 306714 331084
rect 284294 329536 284300 329588
rect 284352 329576 284358 329588
rect 284570 329576 284576 329588
rect 284352 329548 284576 329576
rect 284352 329536 284358 329548
rect 284570 329536 284576 329548
rect 284628 329536 284634 329588
rect 250162 328488 250168 328500
rect 250123 328460 250168 328488
rect 250162 328448 250168 328460
rect 250220 328448 250226 328500
rect 278866 328448 278872 328500
rect 278924 328488 278930 328500
rect 279050 328488 279056 328500
rect 278924 328460 279056 328488
rect 278924 328448 278930 328460
rect 279050 328448 279056 328460
rect 279108 328448 279114 328500
rect 302510 328488 302516 328500
rect 302471 328460 302516 328488
rect 302510 328448 302516 328460
rect 302568 328448 302574 328500
rect 303890 328448 303896 328500
rect 303948 328488 303954 328500
rect 304626 328488 304632 328500
rect 303948 328460 304632 328488
rect 303948 328448 303954 328460
rect 304626 328448 304632 328460
rect 304684 328448 304690 328500
rect 323302 328448 323308 328500
rect 323360 328488 323366 328500
rect 323670 328488 323676 328500
rect 323360 328460 323676 328488
rect 323360 328448 323366 328460
rect 323670 328448 323676 328460
rect 323728 328448 323734 328500
rect 324682 328448 324688 328500
rect 324740 328488 324746 328500
rect 325142 328488 325148 328500
rect 324740 328460 325148 328488
rect 324740 328448 324746 328460
rect 325142 328448 325148 328460
rect 325200 328448 325206 328500
rect 337286 328448 337292 328500
rect 337344 328488 337350 328500
rect 337378 328488 337384 328500
rect 337344 328460 337384 328488
rect 337344 328448 337350 328460
rect 337378 328448 337384 328460
rect 337436 328448 337442 328500
rect 372706 328448 372712 328500
rect 372764 328488 372770 328500
rect 373258 328488 373264 328500
rect 372764 328460 373264 328488
rect 372764 328448 372770 328460
rect 373258 328448 373264 328460
rect 373316 328448 373322 328500
rect 375650 328448 375656 328500
rect 375708 328488 375714 328500
rect 376110 328488 376116 328500
rect 375708 328460 376116 328488
rect 375708 328448 375714 328460
rect 376110 328448 376116 328460
rect 376168 328448 376174 328500
rect 259822 328420 259828 328432
rect 259783 328392 259828 328420
rect 259822 328380 259828 328392
rect 259880 328380 259886 328432
rect 295518 328380 295524 328432
rect 295576 328420 295582 328432
rect 295702 328420 295708 328432
rect 295576 328392 295708 328420
rect 295576 328380 295582 328392
rect 295702 328380 295708 328392
rect 295760 328380 295766 328432
rect 296806 328380 296812 328432
rect 296864 328420 296870 328432
rect 296990 328420 296996 328432
rect 296864 328392 296996 328420
rect 296864 328380 296870 328392
rect 296990 328380 296996 328392
rect 297048 328380 297054 328432
rect 341334 328420 341340 328432
rect 341295 328392 341340 328420
rect 341334 328380 341340 328392
rect 341392 328380 341398 328432
rect 358722 328420 358728 328432
rect 358683 328392 358728 328420
rect 358722 328380 358728 328392
rect 358780 328380 358786 328432
rect 470594 328420 470600 328432
rect 470555 328392 470600 328420
rect 470594 328380 470600 328392
rect 470652 328380 470658 328432
rect 330478 327196 330484 327208
rect 330128 327168 330484 327196
rect 330128 327140 330156 327168
rect 330478 327156 330484 327168
rect 330536 327156 330542 327208
rect 327258 327128 327264 327140
rect 327219 327100 327264 327128
rect 327258 327088 327264 327100
rect 327316 327088 327322 327140
rect 330110 327088 330116 327140
rect 330168 327088 330174 327140
rect 421190 327128 421196 327140
rect 421151 327100 421196 327128
rect 421190 327088 421196 327100
rect 421248 327088 421254 327140
rect 299842 327060 299848 327072
rect 299803 327032 299848 327060
rect 299842 327020 299848 327032
rect 299900 327020 299906 327072
rect 301130 327020 301136 327072
rect 301188 327060 301194 327072
rect 301314 327060 301320 327072
rect 301188 327032 301320 327060
rect 301188 327020 301194 327032
rect 301314 327020 301320 327032
rect 301372 327020 301378 327072
rect 359182 327060 359188 327072
rect 359143 327032 359188 327060
rect 359182 327020 359188 327032
rect 359240 327020 359246 327072
rect 272150 324300 272156 324352
rect 272208 324340 272214 324352
rect 272242 324340 272248 324352
rect 272208 324312 272248 324340
rect 272208 324300 272214 324312
rect 272242 324300 272248 324312
rect 272300 324300 272306 324352
rect 3326 324232 3332 324284
rect 3384 324272 3390 324284
rect 14458 324272 14464 324284
rect 3384 324244 14464 324272
rect 3384 324232 3390 324244
rect 14458 324232 14464 324244
rect 14516 324232 14522 324284
rect 470134 322872 470140 322924
rect 470192 322912 470198 322924
rect 579982 322912 579988 322924
rect 470192 322884 579988 322912
rect 470192 322872 470198 322884
rect 579982 322872 579988 322884
rect 580040 322872 580046 322924
rect 262677 322303 262735 322309
rect 262677 322269 262689 322303
rect 262723 322300 262735 322303
rect 262766 322300 262772 322312
rect 262723 322272 262772 322300
rect 262723 322269 262735 322272
rect 262677 322263 262735 322269
rect 262766 322260 262772 322272
rect 262824 322260 262830 322312
rect 251450 321580 251456 321632
rect 251508 321580 251514 321632
rect 266633 321623 266691 321629
rect 266633 321589 266645 321623
rect 266679 321620 266691 321623
rect 266722 321620 266728 321632
rect 266679 321592 266728 321620
rect 266679 321589 266691 321592
rect 266633 321583 266691 321589
rect 266722 321580 266728 321592
rect 266780 321580 266786 321632
rect 267737 321623 267795 321629
rect 267737 321589 267749 321623
rect 267783 321620 267795 321623
rect 267826 321620 267832 321632
rect 267783 321592 267832 321620
rect 267783 321589 267795 321592
rect 267737 321583 267795 321589
rect 267826 321580 267832 321592
rect 267884 321580 267890 321632
rect 310790 321580 310796 321632
rect 310848 321580 310854 321632
rect 337286 321580 337292 321632
rect 337344 321580 337350 321632
rect 377122 321580 377128 321632
rect 377180 321580 377186 321632
rect 232222 321512 232228 321564
rect 232280 321552 232286 321564
rect 232406 321552 232412 321564
rect 232280 321524 232412 321552
rect 232280 321512 232286 321524
rect 232406 321512 232412 321524
rect 232464 321512 232470 321564
rect 251468 321416 251496 321580
rect 310808 321484 310836 321580
rect 310882 321484 310888 321496
rect 310808 321456 310888 321484
rect 310882 321444 310888 321456
rect 310940 321444 310946 321496
rect 337304 321484 337332 321580
rect 337378 321484 337384 321496
rect 337304 321456 337384 321484
rect 337378 321444 337384 321456
rect 337436 321444 337442 321496
rect 251542 321416 251548 321428
rect 251468 321388 251548 321416
rect 251542 321376 251548 321388
rect 251600 321376 251606 321428
rect 377140 321416 377168 321580
rect 377214 321416 377220 321428
rect 377140 321388 377220 321416
rect 377214 321376 377220 321388
rect 377272 321376 377278 321428
rect 288802 319104 288808 319116
rect 288763 319076 288808 319104
rect 288802 319064 288808 319076
rect 288860 319064 288866 319116
rect 265250 318900 265256 318912
rect 265211 318872 265256 318900
rect 265250 318860 265256 318872
rect 265308 318860 265314 318912
rect 259825 318835 259883 318841
rect 259825 318801 259837 318835
rect 259871 318832 259883 318835
rect 259914 318832 259920 318844
rect 259871 318804 259920 318832
rect 259871 318801 259883 318804
rect 259825 318795 259883 318801
rect 259914 318792 259920 318804
rect 259972 318792 259978 318844
rect 266630 318832 266636 318844
rect 266591 318804 266636 318832
rect 266630 318792 266636 318804
rect 266688 318792 266694 318844
rect 267734 318832 267740 318844
rect 267695 318804 267740 318832
rect 267734 318792 267740 318804
rect 267792 318792 267798 318844
rect 284662 318792 284668 318844
rect 284720 318832 284726 318844
rect 284754 318832 284760 318844
rect 284720 318804 284760 318832
rect 284720 318792 284726 318804
rect 284754 318792 284760 318804
rect 284812 318792 284818 318844
rect 302510 318792 302516 318844
rect 302568 318832 302574 318844
rect 302602 318832 302608 318844
rect 302568 318804 302608 318832
rect 302568 318792 302574 318804
rect 302602 318792 302608 318804
rect 302660 318792 302666 318844
rect 306742 318792 306748 318844
rect 306800 318832 306806 318844
rect 306834 318832 306840 318844
rect 306800 318804 306840 318832
rect 306800 318792 306806 318804
rect 306834 318792 306840 318804
rect 306892 318792 306898 318844
rect 330110 318792 330116 318844
rect 330168 318792 330174 318844
rect 339770 318832 339776 318844
rect 339731 318804 339776 318832
rect 339770 318792 339776 318804
rect 339828 318792 339834 318844
rect 341337 318835 341395 318841
rect 341337 318801 341349 318835
rect 341383 318832 341395 318835
rect 341426 318832 341432 318844
rect 341383 318804 341432 318832
rect 341383 318801 341395 318804
rect 341337 318795 341395 318801
rect 341426 318792 341432 318804
rect 341484 318792 341490 318844
rect 358722 318832 358728 318844
rect 358683 318804 358728 318832
rect 358722 318792 358728 318804
rect 358780 318792 358786 318844
rect 470594 318832 470600 318844
rect 470555 318804 470600 318832
rect 470594 318792 470600 318804
rect 470652 318792 470658 318844
rect 330128 318696 330156 318792
rect 372706 318764 372712 318776
rect 372667 318736 372712 318764
rect 372706 318724 372712 318736
rect 372764 318724 372770 318776
rect 330202 318696 330208 318708
rect 330128 318668 330208 318696
rect 330202 318656 330208 318668
rect 330260 318656 330266 318708
rect 359182 317744 359188 317756
rect 359143 317716 359188 317744
rect 359182 317704 359188 317716
rect 359240 317704 359246 317756
rect 262674 317472 262680 317484
rect 262635 317444 262680 317472
rect 262674 317432 262680 317444
rect 262732 317432 262738 317484
rect 265250 317472 265256 317484
rect 265211 317444 265256 317472
rect 265250 317432 265256 317444
rect 265308 317432 265314 317484
rect 299842 317472 299848 317484
rect 299803 317444 299848 317472
rect 299842 317432 299848 317444
rect 299900 317432 299906 317484
rect 358722 317404 358728 317416
rect 358683 317376 358728 317404
rect 358722 317364 358728 317376
rect 358780 317364 358786 317416
rect 421190 317404 421196 317416
rect 421151 317376 421196 317404
rect 421190 317364 421196 317376
rect 421248 317364 421254 317416
rect 460198 317404 460204 317416
rect 460159 317376 460204 317404
rect 460198 317364 460204 317376
rect 460256 317364 460262 317416
rect 386782 316072 386788 316124
rect 386840 316112 386846 316124
rect 386966 316112 386972 316124
rect 386840 316084 386972 316112
rect 386840 316072 386846 316084
rect 386966 316072 386972 316084
rect 387024 316072 387030 316124
rect 270494 316004 270500 316056
rect 270552 316044 270558 316056
rect 270678 316044 270684 316056
rect 270552 316016 270684 316044
rect 270552 316004 270558 316016
rect 270678 316004 270684 316016
rect 270736 316004 270742 316056
rect 273530 316004 273536 316056
rect 273588 316044 273594 316056
rect 273622 316044 273628 316056
rect 273588 316016 273628 316044
rect 273588 316004 273594 316016
rect 273622 316004 273628 316016
rect 273680 316004 273686 316056
rect 294138 316004 294144 316056
rect 294196 316044 294202 316056
rect 294230 316044 294236 316056
rect 294196 316016 294236 316044
rect 294196 316004 294202 316016
rect 294230 316004 294236 316016
rect 294288 316004 294294 316056
rect 262674 315976 262680 315988
rect 262635 315948 262680 315976
rect 262674 315936 262680 315948
rect 262732 315936 262738 315988
rect 386782 315976 386788 315988
rect 386743 315948 386788 315976
rect 386782 315936 386788 315948
rect 386840 315936 386846 315988
rect 272150 314616 272156 314628
rect 272111 314588 272156 314616
rect 272150 314576 272156 314588
rect 272208 314576 272214 314628
rect 250162 313964 250168 314016
rect 250220 313964 250226 314016
rect 250180 313880 250208 313964
rect 250162 313828 250168 313880
rect 250220 313828 250226 313880
rect 232406 311964 232412 311976
rect 232332 311936 232412 311964
rect 232332 311840 232360 311936
rect 232406 311924 232412 311936
rect 232464 311924 232470 311976
rect 288713 311967 288771 311973
rect 288713 311933 288725 311967
rect 288759 311964 288771 311967
rect 288802 311964 288808 311976
rect 288759 311936 288808 311964
rect 288759 311933 288771 311936
rect 288713 311927 288771 311933
rect 288802 311924 288808 311936
rect 288860 311924 288866 311976
rect 310882 311964 310888 311976
rect 310843 311936 310888 311964
rect 310882 311924 310888 311936
rect 310940 311924 310946 311976
rect 323302 311964 323308 311976
rect 323228 311936 323308 311964
rect 323228 311908 323256 311936
rect 323302 311924 323308 311936
rect 323360 311924 323366 311976
rect 259730 311856 259736 311908
rect 259788 311896 259794 311908
rect 259914 311896 259920 311908
rect 259788 311868 259920 311896
rect 259788 311856 259794 311868
rect 259914 311856 259920 311868
rect 259972 311856 259978 311908
rect 284573 311899 284631 311905
rect 284573 311865 284585 311899
rect 284619 311896 284631 311899
rect 284662 311896 284668 311908
rect 284619 311868 284668 311896
rect 284619 311865 284631 311868
rect 284573 311859 284631 311865
rect 284662 311856 284668 311868
rect 284720 311856 284726 311908
rect 285950 311896 285956 311908
rect 285911 311868 285956 311896
rect 285950 311856 285956 311868
rect 286008 311856 286014 311908
rect 323210 311856 323216 311908
rect 323268 311856 323274 311908
rect 337194 311856 337200 311908
rect 337252 311896 337258 311908
rect 337378 311896 337384 311908
rect 337252 311868 337384 311896
rect 337252 311856 337258 311868
rect 337378 311856 337384 311868
rect 337436 311856 337442 311908
rect 341242 311856 341248 311908
rect 341300 311896 341306 311908
rect 341426 311896 341432 311908
rect 341300 311868 341432 311896
rect 341300 311856 341306 311868
rect 341426 311856 341432 311868
rect 341484 311856 341490 311908
rect 232314 311788 232320 311840
rect 232372 311788 232378 311840
rect 244458 311828 244464 311840
rect 244419 311800 244464 311828
rect 244458 311788 244464 311800
rect 244516 311788 244522 311840
rect 339678 311788 339684 311840
rect 339736 311828 339742 311840
rect 339862 311828 339868 311840
rect 339736 311800 339868 311828
rect 339736 311788 339742 311800
rect 339862 311788 339868 311800
rect 339920 311788 339926 311840
rect 273438 309312 273444 309324
rect 273399 309284 273444 309312
rect 273438 309272 273444 309284
rect 273496 309272 273502 309324
rect 266630 309204 266636 309256
rect 266688 309204 266694 309256
rect 244458 309176 244464 309188
rect 244419 309148 244464 309176
rect 244458 309136 244464 309148
rect 244516 309136 244522 309188
rect 266648 309120 266676 309204
rect 289998 309136 290004 309188
rect 290056 309176 290062 309188
rect 290090 309176 290096 309188
rect 290056 309148 290096 309176
rect 290056 309136 290062 309148
rect 290090 309136 290096 309148
rect 290148 309136 290154 309188
rect 372706 309176 372712 309188
rect 372667 309148 372712 309176
rect 372706 309136 372712 309148
rect 372764 309136 372770 309188
rect 236270 309108 236276 309120
rect 236231 309080 236276 309108
rect 236270 309068 236276 309080
rect 236328 309068 236334 309120
rect 259641 309111 259699 309117
rect 259641 309077 259653 309111
rect 259687 309108 259699 309111
rect 259730 309108 259736 309120
rect 259687 309080 259736 309108
rect 259687 309077 259699 309080
rect 259641 309071 259699 309077
rect 259730 309068 259736 309080
rect 259788 309068 259794 309120
rect 265250 309108 265256 309120
rect 265211 309080 265256 309108
rect 265250 309068 265256 309080
rect 265308 309068 265314 309120
rect 266630 309068 266636 309120
rect 266688 309068 266694 309120
rect 339862 309108 339868 309120
rect 339823 309080 339868 309108
rect 339862 309068 339868 309080
rect 339920 309068 339926 309120
rect 341153 309111 341211 309117
rect 341153 309077 341165 309111
rect 341199 309108 341211 309111
rect 341242 309108 341248 309120
rect 341199 309080 341248 309108
rect 341199 309077 341211 309080
rect 341153 309071 341211 309077
rect 341242 309068 341248 309080
rect 341300 309068 341306 309120
rect 470594 309108 470600 309120
rect 470555 309080 470600 309108
rect 470594 309068 470600 309080
rect 470652 309068 470658 309120
rect 327258 309000 327264 309052
rect 327316 309040 327322 309052
rect 327350 309040 327356 309052
rect 327316 309012 327356 309040
rect 327316 309000 327322 309012
rect 327350 309000 327356 309012
rect 327408 309000 327414 309052
rect 2774 308796 2780 308848
rect 2832 308836 2838 308848
rect 5350 308836 5356 308848
rect 2832 308808 5356 308836
rect 2832 308796 2838 308808
rect 5350 308796 5356 308808
rect 5408 308796 5414 308848
rect 310698 307844 310704 307896
rect 310756 307884 310762 307896
rect 310885 307887 310943 307893
rect 310885 307884 310897 307887
rect 310756 307856 310897 307884
rect 310756 307844 310762 307856
rect 310885 307853 310897 307856
rect 310931 307853 310943 307887
rect 310885 307847 310943 307853
rect 301038 307776 301044 307828
rect 301096 307816 301102 307828
rect 301222 307816 301228 307828
rect 301096 307788 301228 307816
rect 301096 307776 301102 307788
rect 301222 307776 301228 307788
rect 301280 307776 301286 307828
rect 358722 307816 358728 307828
rect 358683 307788 358728 307816
rect 358722 307776 358728 307788
rect 358780 307776 358786 307828
rect 421190 307816 421196 307828
rect 421151 307788 421196 307816
rect 421190 307776 421196 307788
rect 421248 307776 421254 307828
rect 460198 307816 460204 307828
rect 460159 307788 460204 307816
rect 460198 307776 460204 307788
rect 460256 307776 460262 307828
rect 310698 307748 310704 307760
rect 310659 307720 310704 307748
rect 310698 307708 310704 307720
rect 310756 307708 310762 307760
rect 325602 307708 325608 307760
rect 325660 307748 325666 307760
rect 325970 307748 325976 307760
rect 325660 307720 325976 307748
rect 325660 307708 325666 307720
rect 325970 307708 325976 307720
rect 326028 307708 326034 307760
rect 337013 307751 337071 307757
rect 337013 307717 337025 307751
rect 337059 307748 337071 307751
rect 337194 307748 337200 307760
rect 337059 307720 337200 307748
rect 337059 307717 337071 307720
rect 337013 307711 337071 307717
rect 337194 307708 337200 307720
rect 337252 307708 337258 307760
rect 285766 306416 285772 306468
rect 285824 306456 285830 306468
rect 285953 306459 286011 306465
rect 285953 306456 285965 306459
rect 285824 306428 285965 306456
rect 285824 306416 285830 306428
rect 285953 306425 285965 306428
rect 285999 306425 286011 306459
rect 285953 306419 286011 306425
rect 262674 306348 262680 306400
rect 262732 306388 262738 306400
rect 284570 306388 284576 306400
rect 262732 306360 262777 306388
rect 284531 306360 284576 306388
rect 262732 306348 262738 306360
rect 284570 306348 284576 306360
rect 284628 306348 284634 306400
rect 317506 306348 317512 306400
rect 317564 306388 317570 306400
rect 317690 306388 317696 306400
rect 317564 306360 317696 306388
rect 317564 306348 317570 306360
rect 317690 306348 317696 306360
rect 317748 306348 317754 306400
rect 463694 306348 463700 306400
rect 463752 306388 463758 306400
rect 463878 306388 463884 306400
rect 463752 306360 463884 306388
rect 463752 306348 463758 306360
rect 463878 306348 463884 306360
rect 463936 306348 463942 306400
rect 357802 302268 357808 302320
rect 357860 302268 357866 302320
rect 295610 302132 295616 302184
rect 295668 302132 295674 302184
rect 327261 302175 327319 302181
rect 327261 302141 327273 302175
rect 327307 302172 327319 302175
rect 327350 302172 327356 302184
rect 327307 302144 327356 302172
rect 327307 302141 327319 302144
rect 327261 302135 327319 302141
rect 327350 302132 327356 302144
rect 327408 302132 327414 302184
rect 295628 302104 295656 302132
rect 295702 302104 295708 302116
rect 295628 302076 295708 302104
rect 295702 302064 295708 302076
rect 295760 302064 295766 302116
rect 357820 302104 357848 302268
rect 357894 302104 357900 302116
rect 357820 302076 357900 302104
rect 357894 302064 357900 302076
rect 357952 302064 357958 302116
rect 386782 302104 386788 302116
rect 386743 302076 386788 302104
rect 386782 302064 386788 302076
rect 386840 302064 386846 302116
rect 273441 301563 273499 301569
rect 273441 301529 273453 301563
rect 273487 301560 273499 301563
rect 273530 301560 273536 301572
rect 273487 301532 273536 301560
rect 273487 301529 273499 301532
rect 273441 301523 273499 301529
rect 273530 301520 273536 301532
rect 273588 301520 273594 301572
rect 339862 299928 339868 299940
rect 339823 299900 339868 299928
rect 339862 299888 339868 299900
rect 339920 299888 339926 299940
rect 259638 299588 259644 299600
rect 259599 299560 259644 299588
rect 259638 299548 259644 299560
rect 259696 299548 259702 299600
rect 267826 299588 267832 299600
rect 267752 299560 267832 299588
rect 236273 299523 236331 299529
rect 236273 299489 236285 299523
rect 236319 299520 236331 299523
rect 236454 299520 236460 299532
rect 236319 299492 236460 299520
rect 236319 299489 236331 299492
rect 236273 299483 236331 299489
rect 236454 299480 236460 299492
rect 236512 299480 236518 299532
rect 239122 299480 239128 299532
rect 239180 299520 239186 299532
rect 239306 299520 239312 299532
rect 239180 299492 239312 299520
rect 239180 299480 239186 299492
rect 239306 299480 239312 299492
rect 239364 299480 239370 299532
rect 262582 299480 262588 299532
rect 262640 299520 262646 299532
rect 265250 299520 265256 299532
rect 262640 299492 262720 299520
rect 265211 299492 265256 299520
rect 262640 299480 262646 299492
rect 262692 299464 262720 299492
rect 265250 299480 265256 299492
rect 265308 299480 265314 299532
rect 267752 299464 267780 299560
rect 267826 299548 267832 299560
rect 267884 299548 267890 299600
rect 359274 299588 359280 299600
rect 359108 299560 359280 299588
rect 341150 299520 341156 299532
rect 341111 299492 341156 299520
rect 341150 299480 341156 299492
rect 341208 299480 341214 299532
rect 359108 299464 359136 299560
rect 359274 299548 359280 299560
rect 359332 299548 359338 299600
rect 470594 299520 470600 299532
rect 470555 299492 470600 299520
rect 470594 299480 470600 299492
rect 470652 299480 470658 299532
rect 259638 299412 259644 299464
rect 259696 299452 259702 299464
rect 259822 299452 259828 299464
rect 259696 299424 259828 299452
rect 259696 299412 259702 299424
rect 259822 299412 259828 299424
rect 259880 299412 259886 299464
rect 262674 299412 262680 299464
rect 262732 299412 262738 299464
rect 267734 299412 267740 299464
rect 267792 299412 267798 299464
rect 323302 299452 323308 299464
rect 323263 299424 323308 299452
rect 323302 299412 323308 299424
rect 323360 299412 323366 299464
rect 324682 299452 324688 299464
rect 324643 299424 324688 299452
rect 324682 299412 324688 299424
rect 324740 299412 324746 299464
rect 359090 299412 359096 299464
rect 359148 299412 359154 299464
rect 372706 299452 372712 299464
rect 372667 299424 372712 299452
rect 372706 299412 372712 299424
rect 372764 299412 372770 299464
rect 375653 299455 375711 299461
rect 375653 299421 375665 299455
rect 375699 299452 375711 299455
rect 375742 299452 375748 299464
rect 375699 299424 375748 299452
rect 375699 299421 375711 299424
rect 375653 299415 375711 299421
rect 375742 299412 375748 299424
rect 375800 299412 375806 299464
rect 470042 299412 470048 299464
rect 470100 299452 470106 299464
rect 579798 299452 579804 299464
rect 470100 299424 579804 299452
rect 470100 299412 470106 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 337010 298228 337016 298240
rect 336971 298200 337016 298228
rect 337010 298188 337016 298200
rect 337068 298188 337074 298240
rect 266630 298160 266636 298172
rect 266591 298132 266636 298160
rect 266630 298120 266636 298132
rect 266688 298120 266694 298172
rect 310701 298163 310759 298169
rect 310701 298129 310713 298163
rect 310747 298160 310759 298163
rect 310882 298160 310888 298172
rect 310747 298132 310888 298160
rect 310747 298129 310759 298132
rect 310701 298123 310759 298129
rect 310882 298120 310888 298132
rect 310940 298120 310946 298172
rect 327258 298160 327264 298172
rect 327219 298132 327264 298160
rect 327258 298120 327264 298132
rect 327316 298120 327322 298172
rect 337010 298052 337016 298104
rect 337068 298092 337074 298104
rect 337197 298095 337255 298101
rect 337197 298092 337209 298095
rect 337068 298064 337209 298092
rect 337068 298052 337074 298064
rect 337197 298061 337209 298064
rect 337243 298061 337255 298095
rect 358722 298092 358728 298104
rect 358683 298064 358728 298092
rect 337197 298055 337255 298061
rect 358722 298052 358728 298064
rect 358780 298052 358786 298104
rect 359090 298092 359096 298104
rect 359051 298064 359096 298092
rect 359090 298052 359096 298064
rect 359148 298052 359154 298104
rect 421190 298092 421196 298104
rect 421151 298064 421196 298092
rect 421190 298052 421196 298064
rect 421248 298052 421254 298104
rect 460014 298092 460020 298104
rect 459975 298064 460020 298092
rect 460014 298052 460020 298064
rect 460072 298052 460078 298104
rect 329926 297712 329932 297764
rect 329984 297752 329990 297764
rect 330386 297752 330392 297764
rect 329984 297724 330392 297752
rect 329984 297712 329990 297724
rect 330386 297712 330392 297724
rect 330444 297712 330450 297764
rect 266630 296732 266636 296744
rect 266591 296704 266636 296732
rect 266630 296692 266636 296704
rect 266688 296692 266694 296744
rect 270770 296692 270776 296744
rect 270828 296732 270834 296744
rect 270954 296732 270960 296744
rect 270828 296704 270960 296732
rect 270828 296692 270834 296704
rect 270954 296692 270960 296704
rect 271012 296692 271018 296744
rect 272153 296735 272211 296741
rect 272153 296701 272165 296735
rect 272199 296732 272211 296735
rect 272242 296732 272248 296744
rect 272199 296704 272248 296732
rect 272199 296701 272211 296704
rect 272153 296695 272211 296701
rect 272242 296692 272248 296704
rect 272300 296692 272306 296744
rect 285766 296692 285772 296744
rect 285824 296732 285830 296744
rect 286042 296732 286048 296744
rect 285824 296704 286048 296732
rect 285824 296692 285830 296704
rect 286042 296692 286048 296704
rect 286100 296692 286106 296744
rect 294138 296692 294144 296744
rect 294196 296732 294202 296744
rect 294322 296732 294328 296744
rect 294196 296704 294328 296732
rect 294196 296692 294202 296704
rect 294322 296692 294328 296704
rect 294380 296692 294386 296744
rect 270770 295264 270776 295316
rect 270828 295304 270834 295316
rect 270954 295304 270960 295316
rect 270828 295276 270960 295304
rect 270828 295264 270834 295276
rect 270954 295264 270960 295276
rect 271012 295264 271018 295316
rect 272153 295307 272211 295313
rect 272153 295273 272165 295307
rect 272199 295304 272211 295307
rect 272242 295304 272248 295316
rect 272199 295276 272248 295304
rect 272199 295273 272211 295276
rect 272153 295267 272211 295273
rect 272242 295264 272248 295276
rect 272300 295264 272306 295316
rect 251453 294695 251511 294701
rect 251453 294661 251465 294695
rect 251499 294692 251511 294695
rect 251542 294692 251548 294704
rect 251499 294664 251548 294692
rect 251499 294661 251511 294664
rect 251453 294655 251511 294661
rect 251542 294652 251548 294664
rect 251600 294652 251606 294704
rect 289998 294584 290004 294636
rect 290056 294624 290062 294636
rect 290182 294624 290188 294636
rect 290056 294596 290188 294624
rect 290056 294584 290062 294596
rect 290182 294584 290188 294596
rect 290240 294584 290246 294636
rect 306742 294584 306748 294636
rect 306800 294624 306806 294636
rect 306926 294624 306932 294636
rect 306800 294596 306932 294624
rect 306800 294584 306806 294596
rect 306926 294584 306932 294596
rect 306984 294584 306990 294636
rect 310882 293060 310888 293072
rect 310843 293032 310888 293060
rect 310882 293020 310888 293032
rect 310940 293020 310946 293072
rect 386782 293060 386788 293072
rect 386743 293032 386788 293060
rect 386782 293020 386788 293032
rect 386840 293020 386846 293072
rect 236270 292544 236276 292596
rect 236328 292584 236334 292596
rect 236454 292584 236460 292596
rect 236328 292556 236460 292584
rect 236328 292544 236334 292556
rect 236454 292544 236460 292556
rect 236512 292544 236518 292596
rect 296806 292544 296812 292596
rect 296864 292544 296870 292596
rect 301038 292544 301044 292596
rect 301096 292544 301102 292596
rect 357434 292544 357440 292596
rect 357492 292584 357498 292596
rect 357894 292584 357900 292596
rect 357492 292556 357900 292584
rect 357492 292544 357498 292556
rect 357894 292544 357900 292556
rect 357952 292544 357958 292596
rect 239030 292476 239036 292528
rect 239088 292516 239094 292528
rect 239214 292516 239220 292528
rect 239088 292488 239220 292516
rect 239088 292476 239094 292488
rect 239214 292476 239220 292488
rect 239272 292476 239278 292528
rect 296824 292516 296852 292544
rect 296898 292516 296904 292528
rect 296824 292488 296904 292516
rect 296898 292476 296904 292488
rect 296956 292476 296962 292528
rect 301056 292516 301084 292544
rect 301130 292516 301136 292528
rect 301056 292488 301136 292516
rect 301130 292476 301136 292488
rect 301188 292476 301194 292528
rect 337194 292448 337200 292460
rect 337155 292420 337200 292448
rect 337194 292408 337200 292420
rect 337252 292408 337258 292460
rect 285766 291864 285772 291916
rect 285824 291904 285830 291916
rect 286042 291904 286048 291916
rect 285824 291876 286048 291904
rect 285824 291864 285830 291876
rect 286042 291864 286048 291876
rect 286100 291864 286106 291916
rect 288710 290000 288716 290012
rect 288671 289972 288716 290000
rect 288710 289960 288716 289972
rect 288768 289960 288774 290012
rect 251450 289864 251456 289876
rect 251411 289836 251456 289864
rect 251450 289824 251456 289836
rect 251508 289824 251514 289876
rect 299750 289824 299756 289876
rect 299808 289864 299814 289876
rect 299842 289864 299848 289876
rect 299808 289836 299848 289864
rect 299808 289824 299814 289836
rect 299842 289824 299848 289836
rect 299900 289824 299906 289876
rect 324682 289864 324688 289876
rect 324643 289836 324688 289864
rect 324682 289824 324688 289836
rect 324740 289824 324746 289876
rect 372706 289864 372712 289876
rect 372667 289836 372712 289864
rect 372706 289824 372712 289836
rect 372764 289824 372770 289876
rect 375650 289864 375656 289876
rect 375611 289836 375656 289864
rect 375650 289824 375656 289836
rect 375708 289824 375714 289876
rect 377122 289824 377128 289876
rect 377180 289864 377186 289876
rect 377214 289864 377220 289876
rect 377180 289836 377220 289864
rect 377180 289824 377186 289836
rect 377214 289824 377220 289836
rect 377272 289824 377278 289876
rect 250070 289756 250076 289808
rect 250128 289796 250134 289808
rect 250346 289796 250352 289808
rect 250128 289768 250352 289796
rect 250128 289756 250134 289768
rect 250346 289756 250352 289768
rect 250404 289756 250410 289808
rect 259730 289756 259736 289808
rect 259788 289796 259794 289808
rect 259914 289796 259920 289808
rect 259788 289768 259920 289796
rect 259788 289756 259794 289768
rect 259914 289756 259920 289768
rect 259972 289756 259978 289808
rect 284570 289756 284576 289808
rect 284628 289756 284634 289808
rect 288710 289756 288716 289808
rect 288768 289796 288774 289808
rect 288802 289796 288808 289808
rect 288768 289768 288808 289796
rect 288768 289756 288774 289768
rect 288802 289756 288808 289768
rect 288860 289756 288866 289808
rect 289998 289756 290004 289808
rect 290056 289796 290062 289808
rect 290182 289796 290188 289808
rect 290056 289768 290188 289796
rect 290056 289756 290062 289768
rect 290182 289756 290188 289768
rect 290240 289756 290246 289808
rect 302510 289756 302516 289808
rect 302568 289796 302574 289808
rect 302694 289796 302700 289808
rect 302568 289768 302700 289796
rect 302568 289756 302574 289768
rect 302694 289756 302700 289768
rect 302752 289756 302758 289808
rect 306742 289756 306748 289808
rect 306800 289796 306806 289808
rect 306926 289796 306932 289808
rect 306800 289768 306932 289796
rect 306800 289756 306806 289768
rect 306926 289756 306932 289768
rect 306984 289756 306990 289808
rect 327258 289756 327264 289808
rect 327316 289756 327322 289808
rect 341153 289799 341211 289805
rect 341153 289765 341165 289799
rect 341199 289796 341211 289799
rect 341242 289796 341248 289808
rect 341199 289768 341248 289796
rect 341199 289765 341211 289768
rect 341153 289759 341211 289765
rect 341242 289756 341248 289768
rect 341300 289756 341306 289808
rect 470594 289796 470600 289808
rect 470555 289768 470600 289796
rect 470594 289756 470600 289768
rect 470652 289756 470658 289808
rect 284588 289728 284616 289756
rect 284754 289728 284760 289740
rect 284588 289700 284760 289728
rect 284754 289688 284760 289700
rect 284812 289688 284818 289740
rect 327276 289728 327304 289756
rect 327350 289728 327356 289740
rect 327276 289700 327356 289728
rect 327350 289688 327356 289700
rect 327408 289688 327414 289740
rect 295521 288507 295579 288513
rect 295521 288473 295533 288507
rect 295567 288504 295579 288507
rect 295702 288504 295708 288516
rect 295567 288476 295708 288504
rect 295567 288473 295579 288476
rect 295521 288467 295579 288473
rect 295702 288464 295708 288476
rect 295760 288464 295766 288516
rect 323305 288507 323363 288513
rect 323305 288473 323317 288507
rect 323351 288504 323363 288507
rect 323486 288504 323492 288516
rect 323351 288476 323492 288504
rect 323351 288473 323363 288476
rect 323305 288467 323363 288473
rect 323486 288464 323492 288476
rect 323544 288464 323550 288516
rect 267734 288396 267740 288448
rect 267792 288436 267798 288448
rect 267826 288436 267832 288448
rect 267792 288408 267832 288436
rect 267792 288396 267798 288408
rect 267826 288396 267832 288408
rect 267884 288396 267890 288448
rect 359093 288439 359151 288445
rect 359093 288405 359105 288439
rect 359139 288436 359151 288439
rect 359182 288436 359188 288448
rect 359139 288408 359188 288436
rect 359139 288405 359151 288408
rect 359093 288399 359151 288405
rect 359182 288396 359188 288408
rect 359240 288396 359246 288448
rect 421190 288436 421196 288448
rect 421151 288408 421196 288436
rect 421190 288396 421196 288408
rect 421248 288396 421254 288448
rect 460017 288439 460075 288445
rect 460017 288405 460029 288439
rect 460063 288436 460075 288439
rect 460106 288436 460112 288448
rect 460063 288408 460112 288436
rect 460063 288405 460075 288408
rect 460017 288399 460075 288405
rect 460106 288396 460112 288408
rect 460164 288396 460170 288448
rect 325878 288328 325884 288380
rect 325936 288368 325942 288380
rect 326062 288368 326068 288380
rect 325936 288340 326068 288368
rect 325936 288328 325942 288340
rect 326062 288328 326068 288340
rect 326120 288328 326126 288380
rect 329926 288328 329932 288380
rect 329984 288368 329990 288380
rect 330294 288368 330300 288380
rect 329984 288340 330300 288368
rect 329984 288328 329990 288340
rect 330294 288328 330300 288340
rect 330352 288328 330358 288380
rect 266630 287036 266636 287088
rect 266688 287076 266694 287088
rect 266722 287076 266728 287088
rect 266688 287048 266728 287076
rect 266688 287036 266694 287048
rect 266722 287036 266728 287048
rect 266780 287036 266786 287088
rect 291562 287036 291568 287088
rect 291620 287076 291626 287088
rect 291746 287076 291752 287088
rect 291620 287048 291752 287076
rect 291620 287036 291626 287048
rect 291746 287036 291752 287048
rect 291804 287036 291810 287088
rect 294230 287036 294236 287088
rect 294288 287076 294294 287088
rect 294322 287076 294328 287088
rect 294288 287048 294328 287076
rect 294288 287036 294294 287048
rect 294322 287036 294328 287048
rect 294380 287036 294386 287088
rect 295518 287076 295524 287088
rect 295479 287048 295524 287076
rect 295518 287036 295524 287048
rect 295576 287036 295582 287088
rect 296809 287011 296867 287017
rect 296809 286977 296821 287011
rect 296855 287008 296867 287011
rect 296898 287008 296904 287020
rect 296855 286980 296904 287008
rect 296855 286977 296867 286980
rect 296809 286971 296867 286977
rect 296898 286968 296904 286980
rect 296956 286968 296962 287020
rect 272150 285716 272156 285728
rect 272111 285688 272156 285716
rect 272150 285676 272156 285688
rect 272208 285676 272214 285728
rect 266722 285648 266728 285660
rect 266683 285620 266728 285648
rect 266722 285608 266728 285620
rect 266780 285608 266786 285660
rect 301130 282996 301136 283008
rect 301056 282968 301136 282996
rect 236270 282888 236276 282940
rect 236328 282888 236334 282940
rect 236288 282792 236316 282888
rect 301056 282872 301084 282968
rect 301130 282956 301136 282968
rect 301188 282956 301194 283008
rect 460106 282956 460112 283008
rect 460164 282956 460170 283008
rect 337102 282928 337108 282940
rect 337063 282900 337108 282928
rect 337102 282888 337108 282900
rect 337160 282888 337166 282940
rect 339678 282888 339684 282940
rect 339736 282928 339742 282940
rect 339862 282928 339868 282940
rect 339736 282900 339868 282928
rect 339736 282888 339742 282900
rect 339862 282888 339868 282900
rect 339920 282888 339926 282940
rect 357434 282888 357440 282940
rect 357492 282928 357498 282940
rect 357492 282900 357756 282928
rect 357492 282888 357498 282900
rect 301038 282820 301044 282872
rect 301096 282820 301102 282872
rect 357728 282804 357756 282900
rect 360286 282888 360292 282940
rect 360344 282928 360350 282940
rect 360470 282928 360476 282940
rect 360344 282900 360476 282928
rect 360344 282888 360350 282900
rect 360470 282888 360476 282900
rect 360528 282888 360534 282940
rect 460124 282804 460152 282956
rect 236454 282792 236460 282804
rect 236288 282764 236460 282792
rect 236454 282752 236460 282764
rect 236512 282752 236518 282804
rect 310882 282792 310888 282804
rect 310843 282764 310888 282792
rect 310882 282752 310888 282764
rect 310940 282752 310946 282804
rect 357710 282752 357716 282804
rect 357768 282752 357774 282804
rect 386782 282792 386788 282804
rect 386743 282764 386788 282792
rect 386782 282752 386788 282764
rect 386840 282752 386846 282804
rect 460106 282752 460112 282804
rect 460164 282752 460170 282804
rect 270770 282208 270776 282260
rect 270828 282248 270834 282260
rect 270954 282248 270960 282260
rect 270828 282220 270960 282248
rect 270828 282208 270834 282220
rect 270954 282208 270960 282220
rect 271012 282208 271018 282260
rect 295518 280780 295524 280832
rect 295576 280820 295582 280832
rect 295794 280820 295800 280832
rect 295576 280792 295800 280820
rect 295576 280780 295582 280792
rect 295794 280780 295800 280792
rect 295852 280780 295858 280832
rect 358722 280276 358728 280288
rect 358683 280248 358728 280276
rect 358722 280236 358728 280248
rect 358780 280236 358786 280288
rect 325878 280208 325884 280220
rect 325839 280180 325884 280208
rect 325878 280168 325884 280180
rect 325936 280168 325942 280220
rect 341150 280208 341156 280220
rect 341111 280180 341156 280208
rect 341150 280168 341156 280180
rect 341208 280168 341214 280220
rect 470594 280208 470600 280220
rect 470555 280180 470600 280208
rect 470594 280168 470600 280180
rect 470652 280168 470658 280220
rect 236273 280143 236331 280149
rect 236273 280109 236285 280143
rect 236319 280140 236331 280143
rect 236454 280140 236460 280152
rect 236319 280112 236460 280140
rect 236319 280109 236331 280112
rect 236273 280103 236331 280109
rect 236454 280100 236460 280112
rect 236512 280100 236518 280152
rect 239122 280140 239128 280152
rect 239083 280112 239128 280140
rect 239122 280100 239128 280112
rect 239180 280100 239186 280152
rect 251450 280140 251456 280152
rect 251411 280112 251456 280140
rect 251450 280100 251456 280112
rect 251508 280100 251514 280152
rect 259546 280140 259552 280152
rect 259507 280112 259552 280140
rect 259546 280100 259552 280112
rect 259604 280100 259610 280152
rect 273530 280100 273536 280152
rect 273588 280140 273594 280152
rect 273622 280140 273628 280152
rect 273588 280112 273628 280140
rect 273588 280100 273594 280112
rect 273622 280100 273628 280112
rect 273680 280100 273686 280152
rect 284570 280100 284576 280152
rect 284628 280140 284634 280152
rect 284754 280140 284760 280152
rect 284628 280112 284760 280140
rect 284628 280100 284634 280112
rect 284754 280100 284760 280112
rect 284812 280100 284818 280152
rect 336918 280140 336924 280152
rect 336879 280112 336924 280140
rect 336918 280100 336924 280112
rect 336976 280100 336982 280152
rect 359090 280100 359096 280152
rect 359148 280140 359154 280152
rect 359182 280140 359188 280152
rect 359148 280112 359188 280140
rect 359148 280100 359154 280112
rect 359182 280100 359188 280112
rect 359240 280100 359246 280152
rect 372706 280140 372712 280152
rect 372667 280112 372712 280140
rect 372706 280100 372712 280112
rect 372764 280100 372770 280152
rect 377122 280140 377128 280152
rect 377083 280112 377128 280140
rect 377122 280100 377128 280112
rect 377180 280100 377186 280152
rect 460106 280140 460112 280152
rect 460067 280112 460112 280140
rect 460106 280100 460112 280112
rect 460164 280100 460170 280152
rect 265250 278916 265256 278928
rect 265176 278888 265256 278916
rect 250070 278740 250076 278792
rect 250128 278780 250134 278792
rect 250162 278780 250168 278792
rect 250128 278752 250168 278780
rect 250128 278740 250134 278752
rect 250162 278740 250168 278752
rect 250220 278740 250226 278792
rect 265176 278712 265204 278888
rect 265250 278876 265256 278888
rect 265308 278876 265314 278928
rect 285766 278740 285772 278792
rect 285824 278780 285830 278792
rect 286042 278780 286048 278792
rect 285824 278752 286048 278780
rect 285824 278740 285830 278752
rect 286042 278740 286048 278752
rect 286100 278740 286106 278792
rect 288710 278740 288716 278792
rect 288768 278780 288774 278792
rect 288802 278780 288808 278792
rect 288768 278752 288808 278780
rect 288768 278740 288774 278752
rect 288802 278740 288808 278752
rect 288860 278740 288866 278792
rect 294230 278740 294236 278792
rect 294288 278780 294294 278792
rect 294322 278780 294328 278792
rect 294288 278752 294328 278780
rect 294288 278740 294294 278752
rect 294322 278740 294328 278752
rect 294380 278740 294386 278792
rect 323210 278740 323216 278792
rect 323268 278780 323274 278792
rect 323302 278780 323308 278792
rect 323268 278752 323308 278780
rect 323268 278740 323274 278752
rect 323302 278740 323308 278752
rect 323360 278740 323366 278792
rect 325878 278780 325884 278792
rect 325839 278752 325884 278780
rect 325878 278740 325884 278752
rect 325936 278740 325942 278792
rect 337102 278780 337108 278792
rect 337063 278752 337108 278780
rect 337102 278740 337108 278752
rect 337160 278740 337166 278792
rect 265342 278712 265348 278724
rect 265176 278684 265348 278712
rect 265342 278672 265348 278684
rect 265400 278672 265406 278724
rect 310882 278712 310888 278724
rect 310843 278684 310888 278712
rect 310882 278672 310888 278684
rect 310940 278672 310946 278724
rect 386782 278712 386788 278724
rect 386743 278684 386788 278712
rect 386782 278672 386788 278684
rect 386840 278672 386846 278724
rect 291562 277448 291568 277500
rect 291620 277448 291626 277500
rect 291580 277364 291608 277448
rect 291562 277312 291568 277364
rect 291620 277312 291626 277364
rect 266722 276060 266728 276072
rect 266683 276032 266728 276060
rect 266722 276020 266728 276032
rect 266780 276020 266786 276072
rect 296809 276063 296867 276069
rect 296809 276029 296821 276063
rect 296855 276060 296867 276063
rect 297082 276060 297088 276072
rect 296855 276032 297088 276060
rect 296855 276029 296867 276032
rect 296809 276023 296867 276029
rect 297082 276020 297088 276032
rect 297140 276020 297146 276072
rect 463786 275312 463792 275324
rect 463747 275284 463792 275312
rect 463786 275272 463792 275284
rect 463844 275272 463850 275324
rect 266630 274632 266636 274644
rect 266591 274604 266636 274632
rect 266630 274592 266636 274604
rect 266688 274592 266694 274644
rect 330110 273952 330116 273964
rect 330071 273924 330116 273952
rect 330110 273912 330116 273924
rect 330168 273912 330174 273964
rect 250162 273340 250168 273352
rect 250088 273312 250168 273340
rect 250088 273216 250116 273312
rect 250162 273300 250168 273312
rect 250220 273300 250226 273352
rect 250070 273164 250076 273216
rect 250128 273164 250134 273216
rect 460106 273136 460112 273148
rect 460067 273108 460112 273136
rect 460106 273096 460112 273108
rect 460164 273096 460170 273148
rect 259546 273068 259552 273080
rect 259507 273040 259552 273068
rect 259546 273028 259552 273040
rect 259604 273028 259610 273080
rect 367002 270648 367008 270700
rect 367060 270648 367066 270700
rect 367020 270564 367048 270648
rect 236270 270552 236276 270564
rect 236231 270524 236276 270552
rect 236270 270512 236276 270524
rect 236328 270512 236334 270564
rect 239125 270555 239183 270561
rect 239125 270521 239137 270555
rect 239171 270552 239183 270555
rect 239214 270552 239220 270564
rect 239171 270524 239220 270552
rect 239171 270521 239183 270524
rect 239125 270515 239183 270521
rect 239214 270512 239220 270524
rect 239272 270512 239278 270564
rect 251450 270552 251456 270564
rect 251411 270524 251456 270552
rect 251450 270512 251456 270524
rect 251508 270512 251514 270564
rect 324682 270512 324688 270564
rect 324740 270552 324746 270564
rect 324774 270552 324780 270564
rect 324740 270524 324780 270552
rect 324740 270512 324746 270524
rect 324774 270512 324780 270524
rect 324832 270512 324838 270564
rect 325878 270512 325884 270564
rect 325936 270552 325942 270564
rect 325970 270552 325976 270564
rect 325936 270524 325976 270552
rect 325936 270512 325942 270524
rect 325970 270512 325976 270524
rect 326028 270512 326034 270564
rect 336918 270552 336924 270564
rect 336879 270524 336924 270552
rect 336918 270512 336924 270524
rect 336976 270512 336982 270564
rect 367002 270512 367008 270564
rect 367060 270512 367066 270564
rect 372706 270552 372712 270564
rect 372667 270524 372712 270552
rect 372706 270512 372712 270524
rect 372764 270512 372770 270564
rect 377122 270552 377128 270564
rect 377083 270524 377128 270552
rect 377122 270512 377128 270524
rect 377180 270512 377186 270564
rect 463789 270555 463847 270561
rect 463789 270521 463801 270555
rect 463835 270552 463847 270555
rect 463878 270552 463884 270564
rect 463835 270524 463884 270552
rect 463835 270521 463847 270524
rect 463789 270515 463847 270521
rect 463878 270512 463884 270524
rect 463936 270512 463942 270564
rect 341153 270487 341211 270493
rect 341153 270453 341165 270487
rect 341199 270484 341211 270487
rect 341242 270484 341248 270496
rect 341199 270456 341248 270484
rect 341199 270453 341211 270456
rect 341153 270447 341211 270453
rect 341242 270444 341248 270456
rect 341300 270444 341306 270496
rect 460017 270487 460075 270493
rect 460017 270453 460029 270487
rect 460063 270484 460075 270487
rect 460106 270484 460112 270496
rect 460063 270456 460112 270484
rect 460063 270453 460075 270456
rect 460017 270447 460075 270453
rect 460106 270444 460112 270456
rect 460164 270444 460170 270496
rect 470594 270484 470600 270496
rect 470555 270456 470600 270484
rect 470594 270444 470600 270456
rect 470652 270444 470658 270496
rect 302694 269192 302700 269204
rect 302620 269164 302700 269192
rect 302620 269136 302648 269164
rect 302694 269152 302700 269164
rect 302752 269152 302758 269204
rect 306926 269192 306932 269204
rect 306852 269164 306932 269192
rect 306852 269136 306880 269164
rect 306926 269152 306932 269164
rect 306984 269152 306990 269204
rect 262490 269084 262496 269136
rect 262548 269124 262554 269136
rect 262582 269124 262588 269136
rect 262548 269096 262588 269124
rect 262548 269084 262554 269096
rect 262582 269084 262588 269096
rect 262640 269084 262646 269136
rect 284570 269084 284576 269136
rect 284628 269124 284634 269136
rect 284754 269124 284760 269136
rect 284628 269096 284760 269124
rect 284628 269084 284634 269096
rect 284754 269084 284760 269096
rect 284812 269084 284818 269136
rect 290090 269084 290096 269136
rect 290148 269124 290154 269136
rect 290182 269124 290188 269136
rect 290148 269096 290188 269124
rect 290148 269084 290154 269096
rect 290182 269084 290188 269096
rect 290240 269084 290246 269136
rect 301038 269084 301044 269136
rect 301096 269124 301102 269136
rect 301222 269124 301228 269136
rect 301096 269096 301228 269124
rect 301096 269084 301102 269096
rect 301222 269084 301228 269096
rect 301280 269084 301286 269136
rect 302602 269084 302608 269136
rect 302660 269084 302666 269136
rect 306834 269084 306840 269136
rect 306892 269084 306898 269136
rect 358538 269084 358544 269136
rect 358596 269124 358602 269136
rect 358630 269124 358636 269136
rect 358596 269096 358636 269124
rect 358596 269084 358602 269096
rect 358630 269084 358636 269096
rect 358688 269084 358694 269136
rect 421190 269084 421196 269136
rect 421248 269124 421254 269136
rect 421374 269124 421380 269136
rect 421248 269096 421380 269124
rect 421248 269084 421254 269096
rect 421374 269084 421380 269096
rect 421432 269084 421438 269136
rect 250070 269056 250076 269068
rect 250031 269028 250076 269056
rect 250070 269016 250076 269028
rect 250128 269016 250134 269068
rect 288710 267724 288716 267776
rect 288768 267764 288774 267776
rect 288802 267764 288808 267776
rect 288768 267736 288808 267764
rect 288768 267724 288774 267736
rect 288802 267724 288808 267736
rect 288860 267724 288866 267776
rect 291562 267724 291568 267776
rect 291620 267764 291626 267776
rect 291654 267764 291660 267776
rect 291620 267736 291660 267764
rect 291620 267724 291626 267736
rect 291654 267724 291660 267736
rect 291712 267724 291718 267776
rect 295610 267724 295616 267776
rect 295668 267764 295674 267776
rect 295794 267764 295800 267776
rect 295668 267736 295800 267764
rect 295668 267724 295674 267736
rect 295794 267724 295800 267736
rect 295852 267724 295858 267776
rect 294230 264936 294236 264988
rect 294288 264976 294294 264988
rect 294322 264976 294328 264988
rect 294288 264948 294328 264976
rect 294288 264936 294294 264948
rect 294322 264936 294328 264948
rect 294380 264936 294386 264988
rect 270678 263576 270684 263628
rect 270736 263576 270742 263628
rect 339678 263576 339684 263628
rect 339736 263616 339742 263628
rect 339862 263616 339868 263628
rect 339736 263588 339868 263616
rect 339736 263576 339742 263588
rect 339862 263576 339868 263588
rect 339920 263576 339926 263628
rect 360286 263576 360292 263628
rect 360344 263616 360350 263628
rect 360470 263616 360476 263628
rect 360344 263588 360476 263616
rect 360344 263576 360350 263588
rect 360470 263576 360476 263588
rect 360528 263576 360534 263628
rect 270696 263492 270724 263576
rect 270678 263440 270684 263492
rect 270736 263440 270742 263492
rect 310882 263480 310888 263492
rect 310843 263452 310888 263480
rect 310882 263440 310888 263452
rect 310940 263440 310946 263492
rect 386782 263480 386788 263492
rect 386743 263452 386788 263480
rect 386782 263440 386788 263452
rect 386840 263440 386846 263492
rect 325970 260924 325976 260976
rect 326028 260924 326034 260976
rect 460014 260964 460020 260976
rect 459975 260936 460020 260964
rect 460014 260924 460020 260936
rect 460072 260924 460078 260976
rect 284570 260856 284576 260908
rect 284628 260896 284634 260908
rect 284754 260896 284760 260908
rect 284628 260868 284760 260896
rect 284628 260856 284634 260868
rect 284754 260856 284760 260868
rect 284812 260856 284818 260908
rect 236273 260831 236331 260837
rect 236273 260797 236285 260831
rect 236319 260828 236331 260831
rect 236454 260828 236460 260840
rect 236319 260800 236460 260828
rect 236319 260797 236331 260800
rect 236273 260791 236331 260797
rect 236454 260788 236460 260800
rect 236512 260788 236518 260840
rect 239122 260828 239128 260840
rect 239083 260800 239128 260828
rect 239122 260788 239128 260800
rect 239180 260788 239186 260840
rect 251450 260828 251456 260840
rect 251411 260800 251456 260828
rect 251450 260788 251456 260800
rect 251508 260788 251514 260840
rect 259546 260828 259552 260840
rect 259507 260800 259552 260828
rect 259546 260788 259552 260800
rect 259604 260788 259610 260840
rect 262582 260788 262588 260840
rect 262640 260788 262646 260840
rect 266630 260828 266636 260840
rect 266591 260800 266636 260828
rect 266630 260788 266636 260800
rect 266688 260788 266694 260840
rect 267734 260788 267740 260840
rect 267792 260788 267798 260840
rect 270678 260828 270684 260840
rect 270639 260800 270684 260828
rect 270678 260788 270684 260800
rect 270736 260788 270742 260840
rect 273530 260788 273536 260840
rect 273588 260828 273594 260840
rect 273622 260828 273628 260840
rect 273588 260800 273628 260828
rect 273588 260788 273594 260800
rect 273622 260788 273628 260800
rect 273680 260788 273686 260840
rect 262600 260760 262628 260788
rect 262674 260760 262680 260772
rect 262600 260732 262680 260760
rect 262674 260720 262680 260732
rect 262732 260720 262738 260772
rect 267752 260760 267780 260788
rect 325988 260772 326016 260924
rect 330110 260896 330116 260908
rect 330071 260868 330116 260896
rect 330110 260856 330116 260868
rect 330168 260856 330174 260908
rect 341150 260896 341156 260908
rect 341111 260868 341156 260896
rect 341150 260856 341156 260868
rect 341208 260856 341214 260908
rect 470594 260896 470600 260908
rect 470555 260868 470600 260896
rect 470594 260856 470600 260868
rect 470652 260856 470658 260908
rect 336918 260828 336924 260840
rect 336879 260800 336924 260828
rect 336918 260788 336924 260800
rect 336976 260788 336982 260840
rect 372706 260828 372712 260840
rect 372667 260800 372712 260828
rect 372706 260788 372712 260800
rect 372764 260788 372770 260840
rect 377122 260828 377128 260840
rect 377083 260800 377128 260828
rect 377122 260788 377128 260800
rect 377180 260788 377186 260840
rect 460014 260788 460020 260840
rect 460072 260828 460078 260840
rect 460198 260828 460204 260840
rect 460072 260800 460204 260828
rect 460072 260788 460078 260800
rect 460198 260788 460204 260800
rect 460256 260788 460262 260840
rect 463697 260831 463755 260837
rect 463697 260797 463709 260831
rect 463743 260828 463755 260831
rect 463786 260828 463792 260840
rect 463743 260800 463792 260828
rect 463743 260797 463755 260800
rect 463697 260791 463755 260797
rect 463786 260788 463792 260800
rect 463844 260788 463850 260840
rect 267826 260760 267832 260772
rect 267752 260732 267832 260760
rect 267826 260720 267832 260732
rect 267884 260720 267890 260772
rect 325970 260720 325976 260772
rect 326028 260720 326034 260772
rect 327258 259564 327264 259616
rect 327316 259564 327322 259616
rect 250073 259471 250131 259477
rect 250073 259437 250085 259471
rect 250119 259468 250131 259471
rect 250162 259468 250168 259480
rect 250119 259440 250168 259468
rect 250119 259437 250131 259440
rect 250073 259431 250131 259437
rect 250162 259428 250168 259440
rect 250220 259428 250226 259480
rect 272058 259428 272064 259480
rect 272116 259468 272122 259480
rect 272150 259468 272156 259480
rect 272116 259440 272156 259468
rect 272116 259428 272122 259440
rect 272150 259428 272156 259440
rect 272208 259428 272214 259480
rect 327276 259412 327304 259564
rect 336918 259428 336924 259480
rect 336976 259468 336982 259480
rect 337102 259468 337108 259480
rect 336976 259440 337108 259468
rect 336976 259428 336982 259440
rect 337102 259428 337108 259440
rect 337160 259428 337166 259480
rect 299842 259360 299848 259412
rect 299900 259400 299906 259412
rect 300026 259400 300032 259412
rect 299900 259372 300032 259400
rect 299900 259360 299906 259372
rect 300026 259360 300032 259372
rect 300084 259360 300090 259412
rect 302602 259360 302608 259412
rect 302660 259400 302666 259412
rect 302786 259400 302792 259412
rect 302660 259372 302792 259400
rect 302660 259360 302666 259372
rect 302786 259360 302792 259372
rect 302844 259360 302850 259412
rect 327258 259360 327264 259412
rect 327316 259360 327322 259412
rect 358722 259400 358728 259412
rect 358683 259372 358728 259400
rect 358722 259360 358728 259372
rect 358780 259360 358786 259412
rect 250162 259332 250168 259344
rect 250123 259304 250168 259332
rect 250162 259292 250168 259304
rect 250220 259292 250226 259344
rect 267826 258000 267832 258052
rect 267884 258000 267890 258052
rect 272426 258000 272432 258052
rect 272484 258040 272490 258052
rect 272521 258043 272579 258049
rect 272521 258040 272533 258043
rect 272484 258012 272533 258040
rect 272484 258000 272490 258012
rect 272521 258009 272533 258012
rect 272567 258009 272579 258043
rect 272521 258003 272579 258009
rect 267844 257972 267872 258000
rect 268010 257972 268016 257984
rect 267844 257944 268016 257972
rect 268010 257932 268016 257944
rect 268068 257932 268074 257984
rect 295702 256640 295708 256692
rect 295760 256680 295766 256692
rect 295886 256680 295892 256692
rect 295760 256652 295892 256680
rect 295760 256640 295766 256652
rect 295886 256640 295892 256652
rect 295944 256640 295950 256692
rect 310882 256068 310888 256080
rect 310843 256040 310888 256068
rect 310882 256028 310888 256040
rect 310940 256028 310946 256080
rect 265342 255932 265348 255944
rect 265303 255904 265348 255932
rect 265342 255892 265348 255904
rect 265400 255892 265406 255944
rect 337105 254643 337163 254649
rect 337105 254609 337117 254643
rect 337151 254640 337163 254643
rect 337286 254640 337292 254652
rect 337151 254612 337292 254640
rect 337151 254609 337163 254612
rect 337105 254603 337163 254609
rect 337286 254600 337292 254612
rect 337344 254600 337350 254652
rect 323394 254028 323400 254040
rect 323320 254000 323400 254028
rect 323320 253904 323348 254000
rect 323394 253988 323400 254000
rect 323452 253988 323458 254040
rect 386782 254028 386788 254040
rect 386708 254000 386788 254028
rect 327169 253963 327227 253969
rect 327169 253929 327181 253963
rect 327215 253960 327227 253963
rect 327258 253960 327264 253972
rect 327215 253932 327264 253960
rect 327215 253929 327227 253932
rect 327169 253923 327227 253929
rect 327258 253920 327264 253932
rect 327316 253920 327322 253972
rect 386708 253904 386736 254000
rect 386782 253988 386788 254000
rect 386840 253988 386846 254040
rect 323302 253852 323308 253904
rect 323360 253852 323366 253904
rect 357526 253852 357532 253904
rect 357584 253892 357590 253904
rect 357710 253892 357716 253904
rect 357584 253864 357716 253892
rect 357584 253852 357590 253864
rect 357710 253852 357716 253864
rect 357768 253852 357774 253904
rect 358998 253852 359004 253904
rect 359056 253892 359062 253904
rect 359182 253892 359188 253904
rect 359056 253864 359188 253892
rect 359056 253852 359062 253864
rect 359182 253852 359188 253864
rect 359240 253852 359246 253904
rect 386690 253852 386696 253904
rect 386748 253852 386754 253904
rect 259546 253756 259552 253768
rect 259507 253728 259552 253756
rect 259546 253716 259552 253728
rect 259604 253716 259610 253768
rect 2774 252492 2780 252544
rect 2832 252532 2838 252544
rect 5258 252532 5264 252544
rect 2832 252504 5264 252532
rect 2832 252492 2838 252504
rect 5258 252492 5264 252504
rect 5316 252492 5322 252544
rect 469950 252492 469956 252544
rect 470008 252532 470014 252544
rect 580166 252532 580172 252544
rect 470008 252504 580172 252532
rect 470008 252492 470014 252504
rect 580166 252492 580172 252504
rect 580224 252492 580230 252544
rect 296990 251308 296996 251320
rect 296824 251280 296996 251308
rect 236270 251240 236276 251252
rect 236231 251212 236276 251240
rect 236270 251200 236276 251212
rect 236328 251200 236334 251252
rect 239125 251243 239183 251249
rect 239125 251209 239137 251243
rect 239171 251240 239183 251243
rect 239214 251240 239220 251252
rect 239171 251212 239220 251240
rect 239171 251209 239183 251212
rect 239125 251203 239183 251209
rect 239214 251200 239220 251212
rect 239272 251200 239278 251252
rect 251450 251240 251456 251252
rect 251411 251212 251456 251240
rect 251450 251200 251456 251212
rect 251508 251200 251514 251252
rect 289998 251200 290004 251252
rect 290056 251240 290062 251252
rect 290090 251240 290096 251252
rect 290056 251212 290096 251240
rect 290056 251200 290062 251212
rect 290090 251200 290096 251212
rect 290148 251200 290154 251252
rect 259546 251172 259552 251184
rect 259507 251144 259552 251172
rect 259546 251132 259552 251144
rect 259604 251132 259610 251184
rect 266722 251132 266728 251184
rect 266780 251172 266786 251184
rect 266814 251172 266820 251184
rect 266780 251144 266820 251172
rect 266780 251132 266786 251144
rect 266814 251132 266820 251144
rect 266872 251132 266878 251184
rect 296824 251116 296852 251280
rect 296990 251268 296996 251280
rect 297048 251268 297054 251320
rect 310698 251268 310704 251320
rect 310756 251308 310762 251320
rect 310885 251311 310943 251317
rect 310885 251308 310897 251311
rect 310756 251280 310897 251308
rect 310756 251268 310762 251280
rect 310885 251277 310897 251280
rect 310931 251277 310943 251311
rect 310885 251271 310943 251277
rect 372706 251240 372712 251252
rect 372667 251212 372712 251240
rect 372706 251200 372712 251212
rect 372764 251200 372770 251252
rect 377122 251240 377128 251252
rect 377083 251212 377128 251240
rect 377122 251200 377128 251212
rect 377180 251200 377186 251252
rect 463694 251200 463700 251252
rect 463752 251240 463758 251252
rect 463752 251212 463797 251240
rect 463752 251200 463758 251212
rect 310698 251172 310704 251184
rect 310659 251144 310704 251172
rect 310698 251132 310704 251144
rect 310756 251132 310762 251184
rect 367002 251172 367008 251184
rect 366963 251144 367008 251172
rect 367002 251132 367008 251144
rect 367060 251132 367066 251184
rect 470594 251172 470600 251184
rect 470555 251144 470600 251172
rect 470594 251132 470600 251144
rect 470652 251132 470658 251184
rect 250165 251107 250223 251113
rect 250165 251073 250177 251107
rect 250211 251104 250223 251107
rect 250346 251104 250352 251116
rect 250211 251076 250352 251104
rect 250211 251073 250223 251076
rect 250165 251067 250223 251073
rect 250346 251064 250352 251076
rect 250404 251064 250410 251116
rect 296806 251064 296812 251116
rect 296864 251064 296870 251116
rect 284662 249840 284668 249892
rect 284720 249880 284726 249892
rect 284754 249880 284760 249892
rect 284720 249852 284760 249880
rect 284720 249840 284726 249852
rect 284754 249840 284760 249852
rect 284812 249840 284818 249892
rect 285950 249772 285956 249824
rect 286008 249812 286014 249824
rect 286042 249812 286048 249824
rect 286008 249784 286048 249812
rect 286008 249772 286014 249784
rect 286042 249772 286048 249784
rect 286100 249772 286106 249824
rect 336918 249812 336924 249824
rect 336879 249784 336924 249812
rect 336918 249772 336924 249784
rect 336976 249772 336982 249824
rect 421190 249772 421196 249824
rect 421248 249812 421254 249824
rect 421374 249812 421380 249824
rect 421248 249784 421380 249812
rect 421248 249772 421254 249784
rect 421374 249772 421380 249784
rect 421432 249772 421438 249824
rect 272426 249704 272432 249756
rect 272484 249744 272490 249756
rect 272521 249747 272579 249753
rect 272521 249744 272533 249747
rect 272484 249716 272533 249744
rect 272484 249704 272490 249716
rect 272521 249713 272533 249716
rect 272567 249713 272579 249747
rect 284662 249744 284668 249756
rect 284623 249716 284668 249744
rect 272521 249707 272579 249713
rect 284662 249704 284668 249716
rect 284720 249704 284726 249756
rect 265342 248248 265348 248260
rect 265303 248220 265348 248248
rect 265342 248208 265348 248220
rect 265400 248208 265406 248260
rect 289998 246984 290004 247036
rect 290056 247024 290062 247036
rect 290366 247024 290372 247036
rect 290056 246996 290372 247024
rect 290056 246984 290062 246996
rect 290366 246984 290372 246996
rect 290424 246984 290430 247036
rect 294230 246984 294236 247036
rect 294288 246984 294294 247036
rect 294248 246888 294276 246984
rect 294414 246888 294420 246900
rect 294248 246860 294420 246888
rect 294414 246848 294420 246860
rect 294472 246848 294478 246900
rect 288894 245596 288900 245608
rect 288855 245568 288900 245596
rect 288894 245556 288900 245568
rect 288952 245556 288958 245608
rect 285950 244984 285956 244996
rect 285911 244956 285956 244984
rect 285950 244944 285956 244956
rect 286008 244944 286014 244996
rect 341242 244372 341248 244384
rect 341168 244344 341248 244372
rect 339678 244264 339684 244316
rect 339736 244304 339742 244316
rect 339862 244304 339868 244316
rect 339736 244276 339868 244304
rect 339736 244264 339742 244276
rect 339862 244264 339868 244276
rect 339920 244264 339926 244316
rect 341168 244248 341196 244344
rect 341242 244332 341248 244344
rect 341300 244332 341306 244384
rect 460106 244372 460112 244384
rect 460032 244344 460112 244372
rect 360286 244264 360292 244316
rect 360344 244304 360350 244316
rect 360470 244304 360476 244316
rect 360344 244276 360476 244304
rect 360344 244264 360350 244276
rect 360470 244264 360476 244276
rect 360528 244264 360534 244316
rect 460032 244248 460060 244344
rect 460106 244332 460112 244344
rect 460164 244332 460170 244384
rect 341150 244196 341156 244248
rect 341208 244196 341214 244248
rect 460014 244196 460020 244248
rect 460072 244196 460078 244248
rect 259549 244171 259607 244177
rect 259549 244137 259561 244171
rect 259595 244168 259607 244171
rect 259638 244168 259644 244180
rect 259595 244140 259644 244168
rect 259595 244137 259607 244140
rect 259549 244131 259607 244137
rect 259638 244128 259644 244140
rect 259696 244128 259702 244180
rect 271874 243040 271880 243092
rect 271932 243080 271938 243092
rect 272426 243080 272432 243092
rect 271932 243052 272432 243080
rect 271932 243040 271938 243052
rect 272426 243040 272432 243052
rect 272484 243040 272490 243092
rect 306834 241544 306840 241596
rect 306892 241544 306898 241596
rect 324682 241584 324688 241596
rect 324608 241556 324688 241584
rect 236546 241476 236552 241528
rect 236604 241516 236610 241528
rect 236638 241516 236644 241528
rect 236604 241488 236644 241516
rect 236604 241476 236610 241488
rect 236638 241476 236644 241488
rect 236696 241476 236702 241528
rect 266722 241476 266728 241528
rect 266780 241516 266786 241528
rect 266814 241516 266820 241528
rect 266780 241488 266820 241516
rect 266780 241476 266786 241488
rect 266814 241476 266820 241488
rect 266872 241476 266878 241528
rect 306852 241460 306880 241544
rect 324608 241528 324636 241556
rect 324682 241544 324688 241556
rect 324740 241544 324746 241596
rect 325970 241584 325976 241596
rect 325896 241556 325976 241584
rect 325896 241528 325924 241556
rect 325970 241544 325976 241556
rect 326028 241544 326034 241596
rect 337102 241584 337108 241596
rect 337063 241556 337108 241584
rect 337102 241544 337108 241556
rect 337160 241544 337166 241596
rect 310701 241519 310759 241525
rect 310701 241485 310713 241519
rect 310747 241516 310759 241519
rect 310882 241516 310888 241528
rect 310747 241488 310888 241516
rect 310747 241485 310759 241488
rect 310701 241479 310759 241485
rect 310882 241476 310888 241488
rect 310940 241476 310946 241528
rect 323302 241476 323308 241528
rect 323360 241516 323366 241528
rect 323394 241516 323400 241528
rect 323360 241488 323400 241516
rect 323360 241476 323366 241488
rect 323394 241476 323400 241488
rect 323452 241476 323458 241528
rect 324590 241476 324596 241528
rect 324648 241476 324654 241528
rect 325878 241476 325884 241528
rect 325936 241476 325942 241528
rect 357618 241476 357624 241528
rect 357676 241516 357682 241528
rect 357710 241516 357716 241528
rect 357676 241488 357716 241516
rect 357676 241476 357682 241488
rect 357710 241476 357716 241488
rect 357768 241476 357774 241528
rect 359090 241476 359096 241528
rect 359148 241516 359154 241528
rect 359182 241516 359188 241528
rect 359148 241488 359188 241516
rect 359148 241476 359154 241488
rect 359182 241476 359188 241488
rect 359240 241476 359246 241528
rect 367002 241516 367008 241528
rect 366963 241488 367008 241516
rect 367002 241476 367008 241488
rect 367060 241476 367066 241528
rect 470594 241516 470600 241528
rect 470555 241488 470600 241516
rect 470594 241476 470600 241488
rect 470652 241476 470658 241528
rect 299474 241408 299480 241460
rect 299532 241448 299538 241460
rect 299532 241420 299577 241448
rect 299532 241408 299538 241420
rect 306834 241408 306840 241460
rect 306892 241408 306898 241460
rect 259638 241340 259644 241392
rect 259696 241380 259702 241392
rect 259822 241380 259828 241392
rect 259696 241352 259828 241380
rect 259696 241340 259702 241352
rect 259822 241340 259828 241352
rect 259880 241340 259886 241392
rect 270678 240224 270684 240236
rect 270639 240196 270684 240224
rect 270678 240184 270684 240196
rect 270736 240184 270742 240236
rect 327166 240224 327172 240236
rect 327127 240196 327172 240224
rect 327166 240184 327172 240196
rect 327224 240184 327230 240236
rect 284665 240159 284723 240165
rect 284665 240125 284677 240159
rect 284711 240156 284723 240159
rect 284846 240156 284852 240168
rect 284711 240128 284852 240156
rect 284711 240125 284723 240128
rect 284665 240119 284723 240125
rect 284846 240116 284852 240128
rect 284904 240116 284910 240168
rect 299934 240116 299940 240168
rect 299992 240156 299998 240168
rect 300026 240156 300032 240168
rect 299992 240128 300032 240156
rect 299992 240116 299998 240128
rect 300026 240116 300032 240128
rect 300084 240116 300090 240168
rect 302694 240116 302700 240168
rect 302752 240156 302758 240168
rect 302786 240156 302792 240168
rect 302752 240128 302792 240156
rect 302752 240116 302758 240128
rect 302786 240116 302792 240128
rect 302844 240116 302850 240168
rect 358722 240156 358728 240168
rect 358683 240128 358728 240156
rect 358722 240116 358728 240128
rect 358780 240116 358786 240168
rect 267734 240048 267740 240100
rect 267792 240088 267798 240100
rect 267918 240088 267924 240100
rect 267792 240060 267924 240088
rect 267792 240048 267798 240060
rect 267918 240048 267924 240060
rect 267976 240048 267982 240100
rect 291562 240048 291568 240100
rect 291620 240088 291626 240100
rect 291838 240088 291844 240100
rect 291620 240060 291844 240088
rect 291620 240048 291626 240060
rect 291838 240048 291844 240060
rect 291896 240048 291902 240100
rect 324590 240088 324596 240100
rect 324551 240060 324596 240088
rect 324590 240048 324596 240060
rect 324648 240048 324654 240100
rect 327166 240088 327172 240100
rect 327127 240060 327172 240088
rect 327166 240048 327172 240060
rect 327224 240048 327230 240100
rect 270678 238728 270684 238740
rect 270639 238700 270684 238728
rect 270678 238688 270684 238700
rect 270736 238688 270742 238740
rect 3050 237328 3056 237380
rect 3108 237368 3114 237380
rect 15838 237368 15844 237380
rect 3108 237340 15844 237368
rect 3108 237328 3114 237340
rect 15838 237328 15844 237340
rect 15896 237328 15902 237380
rect 288897 236011 288955 236017
rect 288897 235977 288909 236011
rect 288943 236008 288955 236011
rect 288986 236008 288992 236020
rect 288943 235980 288992 236008
rect 288943 235977 288955 235980
rect 288897 235971 288955 235977
rect 288986 235968 288992 235980
rect 289044 235968 289050 236020
rect 262585 235943 262643 235949
rect 262585 235909 262597 235943
rect 262631 235940 262643 235943
rect 262766 235940 262772 235952
rect 262631 235912 262772 235940
rect 262631 235909 262643 235912
rect 262585 235903 262643 235909
rect 262766 235900 262772 235912
rect 262824 235900 262830 235952
rect 265158 234676 265164 234728
rect 265216 234716 265222 234728
rect 265342 234716 265348 234728
rect 265216 234688 265348 234716
rect 265216 234676 265222 234688
rect 265342 234676 265348 234688
rect 265400 234676 265406 234728
rect 310882 234716 310888 234728
rect 310808 234688 310888 234716
rect 310808 234592 310836 234688
rect 310882 234676 310888 234688
rect 310940 234676 310946 234728
rect 323394 234716 323400 234728
rect 323355 234688 323400 234716
rect 323394 234676 323400 234688
rect 323452 234676 323458 234728
rect 337105 234651 337163 234657
rect 337105 234617 337117 234651
rect 337151 234648 337163 234651
rect 337194 234648 337200 234660
rect 337151 234620 337200 234648
rect 337151 234617 337163 234620
rect 337105 234611 337163 234617
rect 337194 234608 337200 234620
rect 337252 234608 337258 234660
rect 273438 234540 273444 234592
rect 273496 234580 273502 234592
rect 273622 234580 273628 234592
rect 273496 234552 273628 234580
rect 273496 234540 273502 234552
rect 273622 234540 273628 234552
rect 273680 234540 273686 234592
rect 310790 234540 310796 234592
rect 310848 234540 310854 234592
rect 357526 234540 357532 234592
rect 357584 234580 357590 234592
rect 357710 234580 357716 234592
rect 357584 234552 357716 234580
rect 357584 234540 357590 234552
rect 357710 234540 357716 234552
rect 357768 234540 357774 234592
rect 358998 234540 359004 234592
rect 359056 234580 359062 234592
rect 359182 234580 359188 234592
rect 359056 234552 359188 234580
rect 359056 234540 359062 234552
rect 359182 234540 359188 234552
rect 359240 234540 359246 234592
rect 285950 234512 285956 234524
rect 285911 234484 285956 234512
rect 285950 234472 285956 234484
rect 286008 234472 286014 234524
rect 270678 233832 270684 233844
rect 270639 233804 270684 233832
rect 270678 233792 270684 233804
rect 270736 233792 270742 233844
rect 301130 231928 301136 231940
rect 301056 231900 301136 231928
rect 244274 231820 244280 231872
rect 244332 231860 244338 231872
rect 244458 231860 244464 231872
rect 244332 231832 244464 231860
rect 244332 231820 244338 231832
rect 244458 231820 244464 231832
rect 244516 231820 244522 231872
rect 250070 231820 250076 231872
rect 250128 231860 250134 231872
rect 250346 231860 250352 231872
rect 250128 231832 250352 231860
rect 250128 231820 250134 231832
rect 250346 231820 250352 231832
rect 250404 231820 250410 231872
rect 251450 231820 251456 231872
rect 251508 231860 251514 231872
rect 251634 231860 251640 231872
rect 251508 231832 251640 231860
rect 251508 231820 251514 231832
rect 251634 231820 251640 231832
rect 251692 231820 251698 231872
rect 299474 231820 299480 231872
rect 299532 231860 299538 231872
rect 299934 231860 299940 231872
rect 299532 231832 299577 231860
rect 299768 231832 299940 231860
rect 299532 231820 299538 231832
rect 299768 231804 299796 231832
rect 299934 231820 299940 231832
rect 299992 231820 299998 231872
rect 301056 231804 301084 231900
rect 301130 231888 301136 231900
rect 301188 231888 301194 231940
rect 372522 231820 372528 231872
rect 372580 231860 372586 231872
rect 372706 231860 372712 231872
rect 372580 231832 372712 231860
rect 372580 231820 372586 231832
rect 372706 231820 372712 231832
rect 372764 231820 372770 231872
rect 376938 231820 376944 231872
rect 376996 231860 377002 231872
rect 377122 231860 377128 231872
rect 376996 231832 377128 231860
rect 376996 231820 377002 231832
rect 377122 231820 377128 231832
rect 377180 231820 377186 231872
rect 299750 231752 299756 231804
rect 299808 231752 299814 231804
rect 301038 231752 301044 231804
rect 301096 231752 301102 231804
rect 310790 231792 310796 231804
rect 310751 231764 310796 231792
rect 310790 231752 310796 231764
rect 310848 231752 310854 231804
rect 323394 231792 323400 231804
rect 323355 231764 323400 231792
rect 323394 231752 323400 231764
rect 323452 231752 323458 231804
rect 324593 231795 324651 231801
rect 324593 231761 324605 231795
rect 324639 231792 324651 231795
rect 324774 231792 324780 231804
rect 324639 231764 324780 231792
rect 324639 231761 324651 231764
rect 324593 231755 324651 231761
rect 324774 231752 324780 231764
rect 324832 231752 324838 231804
rect 327166 230568 327172 230580
rect 327127 230540 327172 230568
rect 327166 230528 327172 230540
rect 327224 230528 327230 230580
rect 325970 230460 325976 230512
rect 326028 230500 326034 230512
rect 326154 230500 326160 230512
rect 326028 230472 326160 230500
rect 326028 230460 326034 230472
rect 326154 230460 326160 230472
rect 326212 230460 326218 230512
rect 336734 230460 336740 230512
rect 336792 230500 336798 230512
rect 336918 230500 336924 230512
rect 336792 230472 336924 230500
rect 336792 230460 336798 230472
rect 336918 230460 336924 230472
rect 336976 230460 336982 230512
rect 337102 230500 337108 230512
rect 337063 230472 337108 230500
rect 337102 230460 337108 230472
rect 337160 230460 337166 230512
rect 341242 230460 341248 230512
rect 341300 230500 341306 230512
rect 341426 230500 341432 230512
rect 341300 230472 341432 230500
rect 341300 230460 341306 230472
rect 341426 230460 341432 230472
rect 341484 230460 341490 230512
rect 358446 230460 358452 230512
rect 358504 230500 358510 230512
rect 358630 230500 358636 230512
rect 358504 230472 358636 230500
rect 358504 230460 358510 230472
rect 358630 230460 358636 230472
rect 358688 230460 358694 230512
rect 421190 230460 421196 230512
rect 421248 230500 421254 230512
rect 421374 230500 421380 230512
rect 421248 230472 421380 230500
rect 421248 230460 421254 230472
rect 421374 230460 421380 230472
rect 421432 230460 421438 230512
rect 459830 230460 459836 230512
rect 459888 230500 459894 230512
rect 460106 230500 460112 230512
rect 459888 230472 460112 230500
rect 459888 230460 459894 230472
rect 460106 230460 460112 230472
rect 460164 230460 460170 230512
rect 358538 230392 358544 230444
rect 358596 230432 358602 230444
rect 358725 230435 358783 230441
rect 358725 230432 358737 230435
rect 358596 230404 358737 230432
rect 358596 230392 358602 230404
rect 358725 230401 358737 230404
rect 358771 230401 358783 230435
rect 358725 230395 358783 230401
rect 265158 229032 265164 229084
rect 265216 229072 265222 229084
rect 265526 229072 265532 229084
rect 265216 229044 265532 229072
rect 265216 229032 265222 229044
rect 265526 229032 265532 229044
rect 265584 229032 265590 229084
rect 272058 229072 272064 229084
rect 272019 229044 272064 229072
rect 272058 229032 272064 229044
rect 272116 229032 272122 229084
rect 262582 226352 262588 226364
rect 262543 226324 262588 226352
rect 262582 226312 262588 226324
rect 262640 226312 262646 226364
rect 336734 225428 336740 225480
rect 336792 225468 336798 225480
rect 336918 225468 336924 225480
rect 336792 225440 336924 225468
rect 336792 225428 336798 225440
rect 336918 225428 336924 225440
rect 336976 225428 336982 225480
rect 284846 225020 284852 225072
rect 284904 225020 284910 225072
rect 341242 225060 341248 225072
rect 341168 225032 341248 225060
rect 236270 224952 236276 225004
rect 236328 224952 236334 225004
rect 236288 224856 236316 224952
rect 284864 224936 284892 225020
rect 339678 224952 339684 225004
rect 339736 224992 339742 225004
rect 339862 224992 339868 225004
rect 339736 224964 339868 224992
rect 339736 224952 339742 224964
rect 339862 224952 339868 224964
rect 339920 224952 339926 225004
rect 341168 224936 341196 225032
rect 341242 225020 341248 225032
rect 341300 225020 341306 225072
rect 460106 225060 460112 225072
rect 460032 225032 460112 225060
rect 360286 224952 360292 225004
rect 360344 224992 360350 225004
rect 360470 224992 360476 225004
rect 360344 224964 360476 224992
rect 360344 224952 360350 224964
rect 360470 224952 360476 224964
rect 360528 224952 360534 225004
rect 460032 224936 460060 225032
rect 460106 225020 460112 225032
rect 460164 225020 460170 225072
rect 284846 224884 284852 224936
rect 284904 224884 284910 224936
rect 341150 224884 341156 224936
rect 341208 224884 341214 224936
rect 460014 224884 460020 224936
rect 460072 224884 460078 224936
rect 236454 224856 236460 224868
rect 236288 224828 236460 224856
rect 236454 224816 236460 224828
rect 236512 224816 236518 224868
rect 306834 222300 306840 222352
rect 306892 222340 306898 222352
rect 306926 222340 306932 222352
rect 306892 222312 306932 222340
rect 306892 222300 306898 222312
rect 306926 222300 306932 222312
rect 306984 222300 306990 222352
rect 259638 222164 259644 222216
rect 259696 222204 259702 222216
rect 259822 222204 259828 222216
rect 259696 222176 259828 222204
rect 259696 222164 259702 222176
rect 259822 222164 259828 222176
rect 259880 222164 259886 222216
rect 294322 222164 294328 222216
rect 294380 222204 294386 222216
rect 294414 222204 294420 222216
rect 294380 222176 294420 222204
rect 294380 222164 294386 222176
rect 294414 222164 294420 222176
rect 294472 222164 294478 222216
rect 295518 222164 295524 222216
rect 295576 222204 295582 222216
rect 295610 222204 295616 222216
rect 295576 222176 295616 222204
rect 295576 222164 295582 222176
rect 295610 222164 295616 222176
rect 295668 222164 295674 222216
rect 296806 222164 296812 222216
rect 296864 222204 296870 222216
rect 296898 222204 296904 222216
rect 296864 222176 296904 222204
rect 296864 222164 296870 222176
rect 296898 222164 296904 222176
rect 296956 222164 296962 222216
rect 299750 222164 299756 222216
rect 299808 222204 299814 222216
rect 299934 222204 299940 222216
rect 299808 222176 299940 222204
rect 299808 222164 299814 222176
rect 299934 222164 299940 222176
rect 299992 222164 299998 222216
rect 310793 222207 310851 222213
rect 310793 222173 310805 222207
rect 310839 222204 310851 222207
rect 310882 222204 310888 222216
rect 310839 222176 310888 222204
rect 310839 222173 310851 222176
rect 310793 222167 310851 222173
rect 310882 222164 310888 222176
rect 310940 222164 310946 222216
rect 325878 222164 325884 222216
rect 325936 222204 325942 222216
rect 326062 222204 326068 222216
rect 325936 222176 326068 222204
rect 325936 222164 325942 222176
rect 326062 222164 326068 222176
rect 326120 222164 326126 222216
rect 359090 222164 359096 222216
rect 359148 222204 359154 222216
rect 359182 222204 359188 222216
rect 359148 222176 359188 222204
rect 359148 222164 359154 222176
rect 359182 222164 359188 222176
rect 359240 222164 359246 222216
rect 386598 222164 386604 222216
rect 386656 222204 386662 222216
rect 386782 222204 386788 222216
rect 386656 222176 386788 222204
rect 386656 222164 386662 222176
rect 386782 222164 386788 222176
rect 386840 222164 386846 222216
rect 463786 222164 463792 222216
rect 463844 222204 463850 222216
rect 464062 222204 464068 222216
rect 463844 222176 464068 222204
rect 463844 222164 463850 222176
rect 464062 222164 464068 222176
rect 464120 222164 464126 222216
rect 470410 222164 470416 222216
rect 470468 222204 470474 222216
rect 470594 222204 470600 222216
rect 470468 222176 470600 222204
rect 470468 222164 470474 222176
rect 470594 222164 470600 222176
rect 470652 222164 470658 222216
rect 299474 222096 299480 222148
rect 299532 222136 299538 222148
rect 299532 222108 299577 222136
rect 299532 222096 299538 222108
rect 259638 222028 259644 222080
rect 259696 222068 259702 222080
rect 259822 222068 259828 222080
rect 259696 222040 259828 222068
rect 259696 222028 259702 222040
rect 259822 222028 259828 222040
rect 259880 222028 259886 222080
rect 273530 220804 273536 220856
rect 273588 220844 273594 220856
rect 273622 220844 273628 220856
rect 273588 220816 273628 220844
rect 273588 220804 273594 220816
rect 273622 220804 273628 220816
rect 273680 220804 273686 220856
rect 327350 220804 327356 220856
rect 327408 220844 327414 220856
rect 327534 220844 327540 220856
rect 327408 220816 327540 220844
rect 327408 220804 327414 220816
rect 327534 220804 327540 220816
rect 327592 220804 327598 220856
rect 330202 220804 330208 220856
rect 330260 220844 330266 220856
rect 330386 220844 330392 220856
rect 330260 220816 330392 220844
rect 330260 220804 330266 220816
rect 330386 220804 330392 220816
rect 330444 220804 330450 220856
rect 358722 220844 358728 220856
rect 358683 220816 358728 220844
rect 358722 220804 358728 220816
rect 358780 220804 358786 220856
rect 272061 220779 272119 220785
rect 272061 220745 272073 220779
rect 272107 220776 272119 220779
rect 272150 220776 272156 220788
rect 272107 220748 272156 220776
rect 272107 220745 272119 220748
rect 272061 220739 272119 220745
rect 272150 220736 272156 220748
rect 272208 220736 272214 220788
rect 341150 220776 341156 220788
rect 341111 220748 341156 220776
rect 341150 220736 341156 220748
rect 341208 220736 341214 220788
rect 262582 219444 262588 219496
rect 262640 219444 262646 219496
rect 262600 219348 262628 219444
rect 270770 219376 270776 219428
rect 270828 219416 270834 219428
rect 270954 219416 270960 219428
rect 270828 219388 270960 219416
rect 270828 219376 270834 219388
rect 270954 219376 270960 219388
rect 271012 219376 271018 219428
rect 317506 219376 317512 219428
rect 317564 219416 317570 219428
rect 317690 219416 317696 219428
rect 317564 219388 317696 219416
rect 317564 219376 317570 219388
rect 317690 219376 317696 219388
rect 317748 219376 317754 219428
rect 262674 219348 262680 219360
rect 262600 219320 262680 219348
rect 262674 219308 262680 219320
rect 262732 219308 262738 219360
rect 290090 217988 290096 218000
rect 290051 217960 290096 217988
rect 290090 217948 290096 217960
rect 290148 217948 290154 218000
rect 310882 215404 310888 215416
rect 310808 215376 310888 215404
rect 310808 215280 310836 215376
rect 310882 215364 310888 215376
rect 310940 215364 310946 215416
rect 464062 215404 464068 215416
rect 463988 215376 464068 215404
rect 386414 215296 386420 215348
rect 386472 215336 386478 215348
rect 386598 215336 386604 215348
rect 386472 215308 386604 215336
rect 386472 215296 386478 215308
rect 386598 215296 386604 215308
rect 386656 215296 386662 215348
rect 463988 215280 464016 215376
rect 464062 215364 464068 215376
rect 464120 215364 464126 215416
rect 273438 215228 273444 215280
rect 273496 215268 273502 215280
rect 273622 215268 273628 215280
rect 273496 215240 273628 215268
rect 273496 215228 273502 215240
rect 273622 215228 273628 215240
rect 273680 215228 273686 215280
rect 310790 215228 310796 215280
rect 310848 215228 310854 215280
rect 341150 215268 341156 215280
rect 341111 215240 341156 215268
rect 341150 215228 341156 215240
rect 341208 215228 341214 215280
rect 459830 215228 459836 215280
rect 459888 215268 459894 215280
rect 460014 215268 460020 215280
rect 459888 215240 460020 215268
rect 459888 215228 459894 215240
rect 460014 215228 460020 215240
rect 460072 215228 460078 215280
rect 463970 215228 463976 215280
rect 464028 215228 464034 215280
rect 291654 214588 291660 214600
rect 291615 214560 291660 214588
rect 291654 214548 291660 214560
rect 291712 214548 291718 214600
rect 299934 212616 299940 212628
rect 299768 212588 299940 212616
rect 244274 212508 244280 212560
rect 244332 212548 244338 212560
rect 244458 212548 244464 212560
rect 244332 212520 244464 212548
rect 244332 212508 244338 212520
rect 244458 212508 244464 212520
rect 244516 212508 244522 212560
rect 250070 212508 250076 212560
rect 250128 212548 250134 212560
rect 250346 212548 250352 212560
rect 250128 212520 250352 212548
rect 250128 212508 250134 212520
rect 250346 212508 250352 212520
rect 250404 212508 250410 212560
rect 251450 212508 251456 212560
rect 251508 212548 251514 212560
rect 251634 212548 251640 212560
rect 251508 212520 251640 212548
rect 251508 212508 251514 212520
rect 251634 212508 251640 212520
rect 251692 212508 251698 212560
rect 299474 212508 299480 212560
rect 299532 212548 299538 212560
rect 299532 212520 299577 212548
rect 299532 212508 299538 212520
rect 299768 212492 299796 212588
rect 299934 212576 299940 212588
rect 299992 212576 299998 212628
rect 301130 212616 301136 212628
rect 301056 212588 301136 212616
rect 301056 212492 301084 212588
rect 301130 212576 301136 212588
rect 301188 212576 301194 212628
rect 324682 212508 324688 212560
rect 324740 212548 324746 212560
rect 324774 212548 324780 212560
rect 324740 212520 324780 212548
rect 324740 212508 324746 212520
rect 324774 212508 324780 212520
rect 324832 212508 324838 212560
rect 325878 212508 325884 212560
rect 325936 212548 325942 212560
rect 325970 212548 325976 212560
rect 325936 212520 325976 212548
rect 325936 212508 325942 212520
rect 325970 212508 325976 212520
rect 326028 212508 326034 212560
rect 336734 212508 336740 212560
rect 336792 212548 336798 212560
rect 336918 212548 336924 212560
rect 336792 212520 336924 212548
rect 336792 212508 336798 212520
rect 336918 212508 336924 212520
rect 336976 212508 336982 212560
rect 357618 212508 357624 212560
rect 357676 212548 357682 212560
rect 357710 212548 357716 212560
rect 357676 212520 357716 212548
rect 357676 212508 357682 212520
rect 357710 212508 357716 212520
rect 357768 212508 357774 212560
rect 359090 212508 359096 212560
rect 359148 212548 359154 212560
rect 359182 212548 359188 212560
rect 359148 212520 359188 212548
rect 359148 212508 359154 212520
rect 359182 212508 359188 212520
rect 359240 212508 359246 212560
rect 372522 212508 372528 212560
rect 372580 212548 372586 212560
rect 372706 212548 372712 212560
rect 372580 212520 372712 212548
rect 372580 212508 372586 212520
rect 372706 212508 372712 212520
rect 372764 212508 372770 212560
rect 376938 212508 376944 212560
rect 376996 212548 377002 212560
rect 377122 212548 377128 212560
rect 376996 212520 377128 212548
rect 376996 212508 377002 212520
rect 377122 212508 377128 212520
rect 377180 212508 377186 212560
rect 284662 212440 284668 212492
rect 284720 212480 284726 212492
rect 284846 212480 284852 212492
rect 284720 212452 284852 212480
rect 284720 212440 284726 212452
rect 284846 212440 284852 212452
rect 284904 212440 284910 212492
rect 299750 212440 299756 212492
rect 299808 212440 299814 212492
rect 301038 212440 301044 212492
rect 301096 212440 301102 212492
rect 310790 212480 310796 212492
rect 310751 212452 310796 212480
rect 310790 212440 310796 212452
rect 310848 212440 310854 212492
rect 330202 212440 330208 212492
rect 330260 212480 330266 212492
rect 330294 212480 330300 212492
rect 330260 212452 330300 212480
rect 330260 212440 330266 212452
rect 330294 212440 330300 212452
rect 330352 212440 330358 212492
rect 250070 211080 250076 211132
rect 250128 211120 250134 211132
rect 250254 211120 250260 211132
rect 250128 211092 250260 211120
rect 250128 211080 250134 211092
rect 250254 211080 250260 211092
rect 250312 211080 250318 211132
rect 284662 211080 284668 211132
rect 284720 211120 284726 211132
rect 284938 211120 284944 211132
rect 284720 211092 284944 211120
rect 284720 211080 284726 211092
rect 284938 211080 284944 211092
rect 284996 211080 285002 211132
rect 317506 209788 317512 209840
rect 317564 209828 317570 209840
rect 317690 209828 317696 209840
rect 317564 209800 317696 209828
rect 317564 209788 317570 209800
rect 317690 209788 317696 209800
rect 317748 209788 317754 209840
rect 290090 208400 290096 208412
rect 290051 208372 290096 208400
rect 290090 208360 290096 208372
rect 290148 208360 290154 208412
rect 460106 205748 460112 205760
rect 460032 205720 460112 205748
rect 323302 205640 323308 205692
rect 323360 205640 323366 205692
rect 339678 205640 339684 205692
rect 339736 205680 339742 205692
rect 339862 205680 339868 205692
rect 339736 205652 339868 205680
rect 339736 205640 339742 205652
rect 339862 205640 339868 205652
rect 339920 205640 339926 205692
rect 360286 205640 360292 205692
rect 360344 205680 360350 205692
rect 360470 205680 360476 205692
rect 360344 205652 360476 205680
rect 360344 205640 360350 205652
rect 360470 205640 360476 205652
rect 360528 205640 360534 205692
rect 323320 205544 323348 205640
rect 460032 205624 460060 205720
rect 460106 205708 460112 205720
rect 460164 205708 460170 205760
rect 460014 205572 460020 205624
rect 460072 205572 460078 205624
rect 323394 205544 323400 205556
rect 323320 205516 323400 205544
rect 323394 205504 323400 205516
rect 323452 205504 323458 205556
rect 291654 204048 291660 204060
rect 291615 204020 291660 204048
rect 291654 204008 291660 204020
rect 291712 204008 291718 204060
rect 262582 202852 262588 202904
rect 262640 202892 262646 202904
rect 262674 202892 262680 202904
rect 262640 202864 262680 202892
rect 262640 202852 262646 202864
rect 262674 202852 262680 202864
rect 262732 202852 262738 202904
rect 266630 202852 266636 202904
rect 266688 202892 266694 202904
rect 266722 202892 266728 202904
rect 266688 202864 266728 202892
rect 266688 202852 266694 202864
rect 266722 202852 266728 202864
rect 266780 202852 266786 202904
rect 285950 202852 285956 202904
rect 286008 202892 286014 202904
rect 286134 202892 286140 202904
rect 286008 202864 286140 202892
rect 286008 202852 286014 202864
rect 286134 202852 286140 202864
rect 286192 202852 286198 202904
rect 294230 202852 294236 202904
rect 294288 202892 294294 202904
rect 294322 202892 294328 202904
rect 294288 202864 294328 202892
rect 294288 202852 294294 202864
rect 294322 202852 294328 202864
rect 294380 202852 294386 202904
rect 295518 202852 295524 202904
rect 295576 202892 295582 202904
rect 295610 202892 295616 202904
rect 295576 202864 295616 202892
rect 295576 202852 295582 202864
rect 295610 202852 295616 202864
rect 295668 202852 295674 202904
rect 296806 202852 296812 202904
rect 296864 202892 296870 202904
rect 296898 202892 296904 202904
rect 296864 202864 296904 202892
rect 296864 202852 296870 202864
rect 296898 202852 296904 202864
rect 296956 202852 296962 202904
rect 299750 202852 299756 202904
rect 299808 202892 299814 202904
rect 299934 202892 299940 202904
rect 299808 202864 299940 202892
rect 299808 202852 299814 202864
rect 299934 202852 299940 202864
rect 299992 202852 299998 202904
rect 310793 202895 310851 202901
rect 310793 202861 310805 202895
rect 310839 202892 310851 202895
rect 310882 202892 310888 202904
rect 310839 202864 310888 202892
rect 310839 202861 310851 202864
rect 310793 202855 310851 202861
rect 310882 202852 310888 202864
rect 310940 202852 310946 202904
rect 324590 202852 324596 202904
rect 324648 202892 324654 202904
rect 324682 202892 324688 202904
rect 324648 202864 324688 202892
rect 324648 202852 324654 202864
rect 324682 202852 324688 202864
rect 324740 202852 324746 202904
rect 325878 202852 325884 202904
rect 325936 202892 325942 202904
rect 325970 202892 325976 202904
rect 325936 202864 325976 202892
rect 325936 202852 325942 202864
rect 325970 202852 325976 202864
rect 326028 202852 326034 202904
rect 341150 202852 341156 202904
rect 341208 202892 341214 202904
rect 341242 202892 341248 202904
rect 341208 202864 341248 202892
rect 341208 202852 341214 202864
rect 341242 202852 341248 202864
rect 341300 202852 341306 202904
rect 463786 202852 463792 202904
rect 463844 202892 463850 202904
rect 464062 202892 464068 202904
rect 463844 202864 464068 202892
rect 463844 202852 463850 202864
rect 464062 202852 464068 202864
rect 464120 202852 464126 202904
rect 470410 202852 470416 202904
rect 470468 202892 470474 202904
rect 470594 202892 470600 202904
rect 470468 202864 470600 202892
rect 470468 202852 470474 202864
rect 470594 202852 470600 202864
rect 470652 202852 470658 202904
rect 239122 202784 239128 202836
rect 239180 202824 239186 202836
rect 239214 202824 239220 202836
rect 239180 202796 239220 202824
rect 239180 202784 239186 202796
rect 239214 202784 239220 202796
rect 239272 202784 239278 202836
rect 273530 202784 273536 202836
rect 273588 202824 273594 202836
rect 273622 202824 273628 202836
rect 273588 202796 273628 202824
rect 273588 202784 273594 202796
rect 273622 202784 273628 202796
rect 273680 202784 273686 202836
rect 299474 202784 299480 202836
rect 299532 202824 299538 202836
rect 336918 202824 336924 202836
rect 299532 202796 299577 202824
rect 336879 202796 336924 202824
rect 299532 202784 299538 202796
rect 336918 202784 336924 202796
rect 336976 202784 336982 202836
rect 270494 202104 270500 202156
rect 270552 202144 270558 202156
rect 270954 202144 270960 202156
rect 270552 202116 270960 202144
rect 270552 202104 270558 202116
rect 270954 202104 270960 202116
rect 271012 202104 271018 202156
rect 290090 201492 290096 201544
rect 290148 201492 290154 201544
rect 250070 201424 250076 201476
rect 250128 201464 250134 201476
rect 250346 201464 250352 201476
rect 250128 201436 250352 201464
rect 250128 201424 250134 201436
rect 250346 201424 250352 201436
rect 250404 201424 250410 201476
rect 262582 201424 262588 201476
rect 262640 201464 262646 201476
rect 262766 201464 262772 201476
rect 262640 201436 262772 201464
rect 262640 201424 262646 201436
rect 262766 201424 262772 201436
rect 262824 201424 262830 201476
rect 272334 201464 272340 201476
rect 272295 201436 272340 201464
rect 272334 201424 272340 201436
rect 272392 201424 272398 201476
rect 267734 201356 267740 201408
rect 267792 201396 267798 201408
rect 267918 201396 267924 201408
rect 267792 201368 267924 201396
rect 267792 201356 267798 201368
rect 267918 201356 267924 201368
rect 267976 201356 267982 201408
rect 290108 201396 290136 201492
rect 358446 201424 358452 201476
rect 358504 201464 358510 201476
rect 358722 201464 358728 201476
rect 358504 201436 358728 201464
rect 358504 201424 358510 201436
rect 358722 201424 358728 201436
rect 358780 201424 358786 201476
rect 421190 201424 421196 201476
rect 421248 201464 421254 201476
rect 421374 201464 421380 201476
rect 421248 201436 421380 201464
rect 421248 201424 421254 201436
rect 421374 201424 421380 201436
rect 421432 201424 421438 201476
rect 290182 201396 290188 201408
rect 290108 201368 290188 201396
rect 290182 201356 290188 201368
rect 290240 201356 290246 201408
rect 250070 200104 250076 200116
rect 250031 200076 250076 200104
rect 250070 200064 250076 200076
rect 250128 200064 250134 200116
rect 265158 200104 265164 200116
rect 265119 200076 265164 200104
rect 265158 200064 265164 200076
rect 265216 200064 265222 200116
rect 317506 200064 317512 200116
rect 317564 200104 317570 200116
rect 317690 200104 317696 200116
rect 317564 200076 317696 200104
rect 317564 200064 317570 200076
rect 317690 200064 317696 200076
rect 317748 200064 317754 200116
rect 285766 198024 285772 198076
rect 285824 198064 285830 198076
rect 285950 198064 285956 198076
rect 285824 198036 285956 198064
rect 285824 198024 285830 198036
rect 285950 198024 285956 198036
rect 286008 198024 286014 198076
rect 294230 198024 294236 198076
rect 294288 198064 294294 198076
rect 294414 198064 294420 198076
rect 294288 198036 294420 198064
rect 294288 198024 294294 198036
rect 294414 198024 294420 198036
rect 294472 198024 294478 198076
rect 310882 196092 310888 196104
rect 310808 196064 310888 196092
rect 232222 195984 232228 196036
rect 232280 195984 232286 196036
rect 232240 195956 232268 195984
rect 310808 195968 310836 196064
rect 310882 196052 310888 196064
rect 310940 196052 310946 196104
rect 464062 196092 464068 196104
rect 463988 196064 464068 196092
rect 337102 195984 337108 196036
rect 337160 195984 337166 196036
rect 460014 195984 460020 196036
rect 460072 195984 460078 196036
rect 232314 195956 232320 195968
rect 232240 195928 232320 195956
rect 232314 195916 232320 195928
rect 232372 195916 232378 195968
rect 310790 195916 310796 195968
rect 310848 195916 310854 195968
rect 337120 195956 337148 195984
rect 337194 195956 337200 195968
rect 337120 195928 337200 195956
rect 337194 195916 337200 195928
rect 337252 195916 337258 195968
rect 357526 195916 357532 195968
rect 357584 195956 357590 195968
rect 357710 195956 357716 195968
rect 357584 195928 357716 195956
rect 357584 195916 357590 195928
rect 357710 195916 357716 195928
rect 357768 195916 357774 195968
rect 358998 195916 359004 195968
rect 359056 195956 359062 195968
rect 359182 195956 359188 195968
rect 359056 195928 359188 195956
rect 359056 195916 359062 195928
rect 359182 195916 359188 195928
rect 359240 195916 359246 195968
rect 460032 195888 460060 195984
rect 463988 195968 464016 196064
rect 464062 196052 464068 196064
rect 464120 196052 464126 196104
rect 463970 195916 463976 195968
rect 464028 195916 464034 195968
rect 460106 195888 460112 195900
rect 460032 195860 460112 195888
rect 460106 195848 460112 195860
rect 460164 195848 460170 195900
rect 270494 195780 270500 195832
rect 270552 195820 270558 195832
rect 270678 195820 270684 195832
rect 270552 195792 270684 195820
rect 270552 195780 270558 195792
rect 270678 195780 270684 195792
rect 270736 195780 270742 195832
rect 265158 195276 265164 195288
rect 265119 195248 265164 195276
rect 265158 195236 265164 195248
rect 265216 195236 265222 195288
rect 290182 193304 290188 193316
rect 290108 193276 290188 193304
rect 244274 193196 244280 193248
rect 244332 193236 244338 193248
rect 244458 193236 244464 193248
rect 244332 193208 244464 193236
rect 244332 193196 244338 193208
rect 244458 193196 244464 193208
rect 244516 193196 244522 193248
rect 251450 193196 251456 193248
rect 251508 193236 251514 193248
rect 251634 193236 251640 193248
rect 251508 193208 251640 193236
rect 251508 193196 251514 193208
rect 251634 193196 251640 193208
rect 251692 193196 251698 193248
rect 259730 193196 259736 193248
rect 259788 193236 259794 193248
rect 259914 193236 259920 193248
rect 259788 193208 259920 193236
rect 259788 193196 259794 193208
rect 259914 193196 259920 193208
rect 259972 193196 259978 193248
rect 290108 193180 290136 193276
rect 290182 193264 290188 193276
rect 290240 193264 290246 193316
rect 302694 193304 302700 193316
rect 302528 193276 302700 193304
rect 299474 193196 299480 193248
rect 299532 193236 299538 193248
rect 299532 193208 299577 193236
rect 299532 193196 299538 193208
rect 302528 193180 302556 193276
rect 302694 193264 302700 193276
rect 302752 193264 302758 193316
rect 323302 193196 323308 193248
rect 323360 193236 323366 193248
rect 323486 193236 323492 193248
rect 323360 193208 323492 193236
rect 323360 193196 323366 193208
rect 323486 193196 323492 193208
rect 323544 193196 323550 193248
rect 324590 193196 324596 193248
rect 324648 193236 324654 193248
rect 324682 193236 324688 193248
rect 324648 193208 324688 193236
rect 324648 193196 324654 193208
rect 324682 193196 324688 193208
rect 324740 193196 324746 193248
rect 325878 193196 325884 193248
rect 325936 193236 325942 193248
rect 325970 193236 325976 193248
rect 325936 193208 325976 193236
rect 325936 193196 325942 193208
rect 325970 193196 325976 193208
rect 326028 193196 326034 193248
rect 336918 193236 336924 193248
rect 336879 193208 336924 193236
rect 336918 193196 336924 193208
rect 336976 193196 336982 193248
rect 341242 193196 341248 193248
rect 341300 193236 341306 193248
rect 341426 193236 341432 193248
rect 341300 193208 341432 193236
rect 341300 193196 341306 193208
rect 341426 193196 341432 193208
rect 341484 193196 341490 193248
rect 372522 193196 372528 193248
rect 372580 193236 372586 193248
rect 372706 193236 372712 193248
rect 372580 193208 372712 193236
rect 372580 193196 372586 193208
rect 372706 193196 372712 193208
rect 372764 193196 372770 193248
rect 376938 193196 376944 193248
rect 376996 193236 377002 193248
rect 377122 193236 377128 193248
rect 376996 193208 377128 193236
rect 376996 193196 377002 193208
rect 377122 193196 377128 193208
rect 377180 193196 377186 193248
rect 386690 193196 386696 193248
rect 386748 193236 386754 193248
rect 386874 193236 386880 193248
rect 386748 193208 386880 193236
rect 386748 193196 386754 193208
rect 386874 193196 386880 193208
rect 386932 193196 386938 193248
rect 272334 193168 272340 193180
rect 272295 193140 272340 193168
rect 272334 193128 272340 193140
rect 272392 193128 272398 193180
rect 290090 193128 290096 193180
rect 290148 193128 290154 193180
rect 302510 193128 302516 193180
rect 302568 193128 302574 193180
rect 367002 193168 367008 193180
rect 366963 193140 367008 193168
rect 367002 193128 367008 193140
rect 367060 193128 367066 193180
rect 266630 191808 266636 191820
rect 266591 191780 266636 191808
rect 266630 191768 266636 191780
rect 266688 191768 266694 191820
rect 270678 191768 270684 191820
rect 270736 191808 270742 191820
rect 270862 191808 270868 191820
rect 270736 191780 270868 191808
rect 270736 191768 270742 191780
rect 270862 191768 270868 191780
rect 270920 191768 270926 191820
rect 288802 191808 288808 191820
rect 288763 191780 288808 191808
rect 288802 191768 288808 191780
rect 288860 191768 288866 191820
rect 291562 191768 291568 191820
rect 291620 191808 291626 191820
rect 291654 191808 291660 191820
rect 291620 191780 291660 191808
rect 291620 191768 291626 191780
rect 291654 191768 291660 191780
rect 291712 191768 291718 191820
rect 317506 190476 317512 190528
rect 317564 190516 317570 190528
rect 317690 190516 317696 190528
rect 317564 190488 317696 190516
rect 317564 190476 317570 190488
rect 317690 190476 317696 190488
rect 317748 190476 317754 190528
rect 270862 190408 270868 190460
rect 270920 190448 270926 190460
rect 271046 190448 271052 190460
rect 270920 190420 271052 190448
rect 270920 190408 270926 190420
rect 271046 190408 271052 190420
rect 271104 190408 271110 190460
rect 290001 188683 290059 188689
rect 290001 188649 290013 188683
rect 290047 188680 290059 188683
rect 290090 188680 290096 188692
rect 290047 188652 290096 188680
rect 290047 188649 290059 188652
rect 290001 188643 290059 188649
rect 290090 188640 290096 188652
rect 290148 188640 290154 188692
rect 299842 188476 299848 188488
rect 299803 188448 299848 188476
rect 299842 188436 299848 188448
rect 299900 188436 299906 188488
rect 306834 188476 306840 188488
rect 306795 188448 306840 188476
rect 306834 188436 306840 188448
rect 306892 188436 306898 188488
rect 264974 186940 264980 186992
rect 265032 186980 265038 186992
rect 265158 186980 265164 186992
rect 265032 186952 265164 186980
rect 265032 186940 265038 186952
rect 265158 186940 265164 186952
rect 265216 186940 265222 186992
rect 295610 186436 295616 186448
rect 295536 186408 295616 186436
rect 295536 186312 295564 186408
rect 295610 186396 295616 186408
rect 295668 186396 295674 186448
rect 296898 186436 296904 186448
rect 296824 186408 296904 186436
rect 296824 186312 296852 186408
rect 296898 186396 296904 186408
rect 296956 186396 296962 186448
rect 327258 186436 327264 186448
rect 327184 186408 327264 186436
rect 327184 186312 327212 186408
rect 327258 186396 327264 186408
rect 327316 186396 327322 186448
rect 330202 186396 330208 186448
rect 330260 186396 330266 186448
rect 250070 186300 250076 186312
rect 250031 186272 250076 186300
rect 250070 186260 250076 186272
rect 250128 186260 250134 186312
rect 266630 186300 266636 186312
rect 266591 186272 266636 186300
rect 266630 186260 266636 186272
rect 266688 186260 266694 186312
rect 272150 186260 272156 186312
rect 272208 186300 272214 186312
rect 272426 186300 272432 186312
rect 272208 186272 272432 186300
rect 272208 186260 272214 186272
rect 272426 186260 272432 186272
rect 272484 186260 272490 186312
rect 295518 186260 295524 186312
rect 295576 186260 295582 186312
rect 296806 186260 296812 186312
rect 296864 186260 296870 186312
rect 327166 186260 327172 186312
rect 327224 186260 327230 186312
rect 330220 186244 330248 186396
rect 460014 186328 460020 186380
rect 460072 186368 460078 186380
rect 460072 186340 460152 186368
rect 460072 186328 460078 186340
rect 460124 186312 460152 186340
rect 460106 186260 460112 186312
rect 460164 186260 460170 186312
rect 330202 186192 330208 186244
rect 330260 186192 330266 186244
rect 294325 184263 294383 184269
rect 294325 184229 294337 184263
rect 294371 184260 294383 184263
rect 294414 184260 294420 184272
rect 294371 184232 294420 184260
rect 294371 184229 294383 184232
rect 294325 184223 294383 184229
rect 294414 184220 294420 184232
rect 294472 184220 294478 184272
rect 285950 183676 285956 183728
rect 286008 183676 286014 183728
rect 284662 183608 284668 183660
rect 284720 183608 284726 183660
rect 236454 183540 236460 183592
rect 236512 183580 236518 183592
rect 236546 183580 236552 183592
rect 236512 183552 236552 183580
rect 236512 183540 236518 183552
rect 236546 183540 236552 183552
rect 236604 183540 236610 183592
rect 284680 183524 284708 183608
rect 285968 183592 285996 183676
rect 302510 183608 302516 183660
rect 302568 183648 302574 183660
rect 302568 183620 302648 183648
rect 302568 183608 302574 183620
rect 302620 183592 302648 183620
rect 285950 183540 285956 183592
rect 286008 183540 286014 183592
rect 299842 183580 299848 183592
rect 299803 183552 299848 183580
rect 299842 183540 299848 183552
rect 299900 183540 299906 183592
rect 301038 183540 301044 183592
rect 301096 183580 301102 183592
rect 301222 183580 301228 183592
rect 301096 183552 301228 183580
rect 301096 183540 301102 183552
rect 301222 183540 301228 183552
rect 301280 183540 301286 183592
rect 302602 183540 302608 183592
rect 302660 183540 302666 183592
rect 306834 183580 306840 183592
rect 306795 183552 306840 183580
rect 306834 183540 306840 183552
rect 306892 183540 306898 183592
rect 310882 183540 310888 183592
rect 310940 183580 310946 183592
rect 311066 183580 311072 183592
rect 310940 183552 311072 183580
rect 310940 183540 310946 183552
rect 311066 183540 311072 183552
rect 311124 183540 311130 183592
rect 358630 183540 358636 183592
rect 358688 183580 358694 183592
rect 358722 183580 358728 183592
rect 358688 183552 358728 183580
rect 358688 183540 358694 183552
rect 358722 183540 358728 183552
rect 358780 183540 358786 183592
rect 359090 183540 359096 183592
rect 359148 183580 359154 183592
rect 359182 183580 359188 183592
rect 359148 183552 359188 183580
rect 359148 183540 359154 183552
rect 359182 183540 359188 183552
rect 359240 183540 359246 183592
rect 360470 183540 360476 183592
rect 360528 183580 360534 183592
rect 360654 183580 360660 183592
rect 360528 183552 360660 183580
rect 360528 183540 360534 183552
rect 360654 183540 360660 183552
rect 360712 183540 360718 183592
rect 367002 183580 367008 183592
rect 366963 183552 367008 183580
rect 367002 183540 367008 183552
rect 367060 183540 367066 183592
rect 463786 183540 463792 183592
rect 463844 183580 463850 183592
rect 464062 183580 464068 183592
rect 463844 183552 464068 183580
rect 463844 183540 463850 183552
rect 464062 183540 464068 183552
rect 464120 183540 464126 183592
rect 470410 183540 470416 183592
rect 470468 183580 470474 183592
rect 470594 183580 470600 183592
rect 470468 183552 470600 183580
rect 470468 183540 470474 183552
rect 470594 183540 470600 183552
rect 470652 183540 470658 183592
rect 239122 183472 239128 183524
rect 239180 183512 239186 183524
rect 239214 183512 239220 183524
rect 239180 183484 239220 183512
rect 239180 183472 239186 183484
rect 239214 183472 239220 183484
rect 239272 183472 239278 183524
rect 273530 183472 273536 183524
rect 273588 183512 273594 183524
rect 273622 183512 273628 183524
rect 273588 183484 273628 183512
rect 273588 183472 273594 183484
rect 273622 183472 273628 183484
rect 273680 183472 273686 183524
rect 284662 183472 284668 183524
rect 284720 183472 284726 183524
rect 337102 183512 337108 183524
rect 337063 183484 337108 183512
rect 337102 183472 337108 183484
rect 337160 183472 337166 183524
rect 460106 183512 460112 183524
rect 460067 183484 460112 183512
rect 460106 183472 460112 183484
rect 460164 183472 460170 183524
rect 341150 182112 341156 182164
rect 341208 182152 341214 182164
rect 341242 182152 341248 182164
rect 341208 182124 341248 182152
rect 341208 182112 341214 182124
rect 341242 182112 341248 182124
rect 341300 182112 341306 182164
rect 358538 182112 358544 182164
rect 358596 182152 358602 182164
rect 358722 182152 358728 182164
rect 358596 182124 358728 182152
rect 358596 182112 358602 182124
rect 358722 182112 358728 182124
rect 358780 182112 358786 182164
rect 360470 182112 360476 182164
rect 360528 182152 360534 182164
rect 360654 182152 360660 182164
rect 360528 182124 360660 182152
rect 360528 182112 360534 182124
rect 360654 182112 360660 182124
rect 360712 182112 360718 182164
rect 421190 182112 421196 182164
rect 421248 182152 421254 182164
rect 421374 182152 421380 182164
rect 421248 182124 421380 182152
rect 421248 182112 421254 182124
rect 421374 182112 421380 182124
rect 421432 182112 421438 182164
rect 469858 182112 469864 182164
rect 469916 182152 469922 182164
rect 580166 182152 580172 182164
rect 469916 182124 580172 182152
rect 469916 182112 469922 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 357618 180820 357624 180872
rect 357676 180860 357682 180872
rect 357710 180860 357716 180872
rect 357676 180832 357716 180860
rect 357676 180820 357682 180832
rect 357710 180820 357716 180832
rect 357768 180820 357774 180872
rect 284662 180792 284668 180804
rect 284623 180764 284668 180792
rect 284662 180752 284668 180764
rect 284720 180752 284726 180804
rect 299842 180792 299848 180804
rect 299803 180764 299848 180792
rect 299842 180752 299848 180764
rect 299900 180752 299906 180804
rect 301038 180792 301044 180804
rect 300999 180764 301044 180792
rect 301038 180752 301044 180764
rect 301096 180752 301102 180804
rect 302602 180792 302608 180804
rect 302563 180764 302608 180792
rect 302602 180752 302608 180764
rect 302660 180752 302666 180804
rect 317506 180752 317512 180804
rect 317564 180792 317570 180804
rect 317690 180792 317696 180804
rect 317564 180764 317696 180792
rect 317564 180752 317570 180764
rect 317690 180752 317696 180764
rect 317748 180752 317754 180804
rect 259638 179568 259644 179580
rect 259599 179540 259644 179568
rect 259638 179528 259644 179540
rect 259696 179528 259702 179580
rect 288802 179432 288808 179444
rect 288763 179404 288808 179432
rect 288802 179392 288808 179404
rect 288860 179392 288866 179444
rect 289998 179432 290004 179444
rect 289959 179404 290004 179432
rect 289998 179392 290004 179404
rect 290056 179392 290062 179444
rect 294322 179432 294328 179444
rect 294283 179404 294328 179432
rect 294322 179392 294328 179404
rect 294380 179392 294386 179444
rect 295518 178712 295524 178764
rect 295576 178752 295582 178764
rect 295702 178752 295708 178764
rect 295576 178724 295708 178752
rect 295576 178712 295582 178724
rect 295702 178712 295708 178724
rect 295760 178712 295766 178764
rect 296806 178712 296812 178764
rect 296864 178752 296870 178764
rect 296990 178752 296996 178764
rect 296864 178724 296996 178752
rect 296864 178712 296870 178724
rect 296990 178712 296996 178724
rect 297048 178712 297054 178764
rect 294322 177964 294328 178016
rect 294380 178004 294386 178016
rect 294417 178007 294475 178013
rect 294417 178004 294429 178007
rect 294380 177976 294429 178004
rect 294380 177964 294386 177976
rect 294417 177973 294429 177976
rect 294463 177973 294475 178007
rect 294417 177967 294475 177973
rect 250070 177284 250076 177336
rect 250128 177324 250134 177336
rect 250346 177324 250352 177336
rect 250128 177296 250352 177324
rect 250128 177284 250134 177296
rect 250346 177284 250352 177296
rect 250404 177284 250410 177336
rect 310882 176780 310888 176792
rect 310808 176752 310888 176780
rect 232222 176672 232228 176724
rect 232280 176672 232286 176724
rect 232240 176644 232268 176672
rect 310808 176656 310836 176752
rect 310882 176740 310888 176752
rect 310940 176740 310946 176792
rect 357618 176740 357624 176792
rect 357676 176740 357682 176792
rect 357636 176656 357664 176740
rect 463878 176672 463884 176724
rect 463936 176712 463942 176724
rect 464062 176712 464068 176724
rect 463936 176684 464068 176712
rect 463936 176672 463942 176684
rect 464062 176672 464068 176684
rect 464120 176672 464126 176724
rect 232314 176644 232320 176656
rect 232240 176616 232320 176644
rect 232314 176604 232320 176616
rect 232372 176604 232378 176656
rect 288802 176644 288808 176656
rect 288763 176616 288808 176644
rect 288802 176604 288808 176616
rect 288860 176604 288866 176656
rect 310790 176604 310796 176656
rect 310848 176604 310854 176656
rect 357618 176604 357624 176656
rect 357676 176604 357682 176656
rect 372706 176604 372712 176656
rect 372764 176604 372770 176656
rect 372724 176576 372752 176604
rect 372798 176576 372804 176588
rect 372724 176548 372804 176576
rect 372798 176536 372804 176548
rect 372856 176536 372862 176588
rect 460106 176508 460112 176520
rect 460067 176480 460112 176508
rect 460106 176468 460112 176480
rect 460164 176468 460170 176520
rect 259641 173995 259699 174001
rect 259641 173961 259653 173995
rect 259687 173992 259699 173995
rect 259730 173992 259736 174004
rect 259687 173964 259736 173992
rect 259687 173961 259699 173964
rect 259641 173955 259699 173961
rect 259730 173952 259736 173964
rect 259788 173952 259794 174004
rect 236270 173884 236276 173936
rect 236328 173924 236334 173936
rect 236638 173924 236644 173936
rect 236328 173896 236644 173924
rect 236328 173884 236334 173896
rect 236638 173884 236644 173896
rect 236696 173884 236702 173936
rect 251450 173884 251456 173936
rect 251508 173924 251514 173936
rect 251634 173924 251640 173936
rect 251508 173896 251640 173924
rect 251508 173884 251514 173896
rect 251634 173884 251640 173896
rect 251692 173884 251698 173936
rect 262582 173884 262588 173936
rect 262640 173924 262646 173936
rect 262674 173924 262680 173936
rect 262640 173896 262680 173924
rect 262640 173884 262646 173896
rect 262674 173884 262680 173896
rect 262732 173884 262738 173936
rect 266630 173884 266636 173936
rect 266688 173924 266694 173936
rect 266814 173924 266820 173936
rect 266688 173896 266820 173924
rect 266688 173884 266694 173896
rect 266814 173884 266820 173896
rect 266872 173884 266878 173936
rect 267734 173884 267740 173936
rect 267792 173924 267798 173936
rect 267826 173924 267832 173936
rect 267792 173896 267832 173924
rect 267792 173884 267798 173896
rect 267826 173884 267832 173896
rect 267884 173884 267890 173936
rect 323302 173884 323308 173936
rect 323360 173924 323366 173936
rect 323486 173924 323492 173936
rect 323360 173896 323492 173924
rect 323360 173884 323366 173896
rect 323486 173884 323492 173896
rect 323544 173884 323550 173936
rect 324682 173884 324688 173936
rect 324740 173924 324746 173936
rect 324774 173924 324780 173936
rect 324740 173896 324780 173924
rect 324740 173884 324746 173896
rect 324774 173884 324780 173896
rect 324832 173884 324838 173936
rect 325878 173884 325884 173936
rect 325936 173924 325942 173936
rect 325970 173924 325976 173936
rect 325936 173896 325976 173924
rect 325936 173884 325942 173896
rect 325970 173884 325976 173896
rect 326028 173884 326034 173936
rect 327166 173884 327172 173936
rect 327224 173924 327230 173936
rect 327258 173924 327264 173936
rect 327224 173896 327264 173924
rect 327224 173884 327230 173896
rect 327258 173884 327264 173896
rect 327316 173884 327322 173936
rect 336734 173884 336740 173936
rect 336792 173924 336798 173936
rect 336918 173924 336924 173936
rect 336792 173896 336924 173924
rect 336792 173884 336798 173896
rect 336918 173884 336924 173896
rect 336976 173884 336982 173936
rect 376938 173884 376944 173936
rect 376996 173924 377002 173936
rect 377030 173924 377036 173936
rect 376996 173896 377036 173924
rect 376996 173884 377002 173896
rect 377030 173884 377036 173896
rect 377088 173884 377094 173936
rect 386782 173884 386788 173936
rect 386840 173924 386846 173936
rect 386966 173924 386972 173936
rect 386840 173896 386972 173924
rect 386840 173884 386846 173896
rect 386966 173884 386972 173896
rect 387024 173884 387030 173936
rect 339678 173816 339684 173868
rect 339736 173856 339742 173868
rect 339954 173856 339960 173868
rect 339736 173828 339960 173856
rect 339736 173816 339742 173828
rect 339954 173816 339960 173828
rect 340012 173816 340018 173868
rect 270770 172524 270776 172576
rect 270828 172524 270834 172576
rect 272242 172524 272248 172576
rect 272300 172564 272306 172576
rect 272334 172564 272340 172576
rect 272300 172536 272340 172564
rect 272300 172524 272306 172536
rect 272334 172524 272340 172536
rect 272392 172524 272398 172576
rect 337102 172564 337108 172576
rect 337063 172536 337108 172564
rect 337102 172524 337108 172536
rect 337160 172524 337166 172576
rect 270788 172428 270816 172524
rect 330110 172496 330116 172508
rect 330071 172468 330116 172496
rect 330110 172456 330116 172468
rect 330168 172456 330174 172508
rect 270862 172428 270868 172440
rect 270788 172400 270868 172428
rect 270862 172388 270868 172400
rect 270920 172388 270926 172440
rect 284665 171139 284723 171145
rect 284665 171105 284677 171139
rect 284711 171136 284723 171139
rect 284754 171136 284760 171148
rect 284711 171108 284760 171136
rect 284711 171105 284723 171108
rect 284665 171099 284723 171105
rect 284754 171096 284760 171108
rect 284812 171096 284818 171148
rect 299842 171136 299848 171148
rect 299803 171108 299848 171136
rect 299842 171096 299848 171108
rect 299900 171096 299906 171148
rect 301038 171136 301044 171148
rect 300999 171108 301044 171136
rect 301038 171096 301044 171108
rect 301096 171096 301102 171148
rect 302602 171136 302608 171148
rect 302563 171108 302608 171136
rect 302602 171096 302608 171108
rect 302660 171096 302666 171148
rect 306650 171096 306656 171148
rect 306708 171136 306714 171148
rect 306926 171136 306932 171148
rect 306708 171108 306932 171136
rect 306708 171096 306714 171108
rect 306926 171096 306932 171108
rect 306984 171096 306990 171148
rect 285953 171071 286011 171077
rect 285953 171037 285965 171071
rect 285999 171068 286011 171071
rect 286042 171068 286048 171080
rect 285999 171040 286048 171068
rect 285999 171037 286011 171040
rect 285953 171031 286011 171037
rect 286042 171028 286048 171040
rect 286100 171028 286106 171080
rect 337102 169260 337108 169312
rect 337160 169300 337166 169312
rect 337378 169300 337384 169312
rect 337160 169272 337384 169300
rect 337160 169260 337166 169272
rect 337378 169260 337384 169272
rect 337436 169260 337442 169312
rect 259730 169056 259736 169108
rect 259788 169096 259794 169108
rect 259914 169096 259920 169108
rect 259788 169068 259920 169096
rect 259788 169056 259794 169068
rect 259914 169056 259920 169068
rect 259972 169056 259978 169108
rect 294322 168376 294328 168428
rect 294380 168416 294386 168428
rect 294417 168419 294475 168425
rect 294417 168416 294429 168419
rect 294380 168388 294429 168416
rect 294380 168376 294386 168388
rect 294417 168385 294429 168388
rect 294463 168385 294475 168419
rect 294417 168379 294475 168385
rect 272058 167628 272064 167680
rect 272116 167668 272122 167680
rect 272242 167668 272248 167680
rect 272116 167640 272248 167668
rect 272116 167628 272122 167640
rect 272242 167628 272248 167640
rect 272300 167628 272306 167680
rect 357434 167628 357440 167680
rect 357492 167668 357498 167680
rect 357618 167668 357624 167680
rect 357492 167640 357624 167668
rect 357492 167628 357498 167640
rect 357618 167628 357624 167640
rect 357676 167628 357682 167680
rect 270862 167124 270868 167136
rect 270696 167096 270868 167124
rect 270696 167000 270724 167096
rect 270862 167084 270868 167096
rect 270920 167084 270926 167136
rect 288802 167056 288808 167068
rect 288763 167028 288808 167056
rect 288802 167016 288808 167028
rect 288860 167016 288866 167068
rect 310790 167016 310796 167068
rect 310848 167016 310854 167068
rect 270678 166948 270684 167000
rect 270736 166948 270742 167000
rect 310808 166920 310836 167016
rect 460106 166988 460112 167000
rect 460067 166960 460112 166988
rect 460106 166948 460112 166960
rect 460164 166948 460170 167000
rect 310882 166920 310888 166932
rect 310808 166892 310888 166920
rect 310882 166880 310888 166892
rect 310940 166880 310946 166932
rect 2774 165452 2780 165504
rect 2832 165492 2838 165504
rect 5166 165492 5172 165504
rect 2832 165464 5172 165492
rect 2832 165452 2838 165464
rect 5166 165452 5172 165464
rect 5224 165452 5230 165504
rect 262674 164336 262680 164348
rect 262600 164308 262680 164336
rect 262600 164280 262628 164308
rect 262674 164296 262680 164308
rect 262732 164296 262738 164348
rect 265250 164336 265256 164348
rect 265176 164308 265256 164336
rect 265176 164280 265204 164308
rect 265250 164296 265256 164308
rect 265308 164296 265314 164348
rect 267826 164336 267832 164348
rect 267752 164308 267832 164336
rect 267752 164280 267780 164308
rect 267826 164296 267832 164308
rect 267884 164296 267890 164348
rect 262582 164228 262588 164280
rect 262640 164228 262646 164280
rect 265158 164228 265164 164280
rect 265216 164228 265222 164280
rect 267734 164228 267740 164280
rect 267792 164228 267798 164280
rect 239122 164160 239128 164212
rect 239180 164200 239186 164212
rect 239214 164200 239220 164212
rect 239180 164172 239220 164200
rect 239180 164160 239186 164172
rect 239214 164160 239220 164172
rect 239272 164160 239278 164212
rect 244274 164160 244280 164212
rect 244332 164200 244338 164212
rect 244458 164200 244464 164212
rect 244332 164172 244464 164200
rect 244332 164160 244338 164172
rect 244458 164160 244464 164172
rect 244516 164160 244522 164212
rect 251450 164160 251456 164212
rect 251508 164200 251514 164212
rect 251634 164200 251640 164212
rect 251508 164172 251640 164200
rect 251508 164160 251514 164172
rect 251634 164160 251640 164172
rect 251692 164160 251698 164212
rect 259638 164160 259644 164212
rect 259696 164200 259702 164212
rect 259822 164200 259828 164212
rect 259696 164172 259828 164200
rect 259696 164160 259702 164172
rect 259822 164160 259828 164172
rect 259880 164160 259886 164212
rect 372798 164200 372804 164212
rect 372759 164172 372804 164200
rect 372798 164160 372804 164172
rect 372856 164160 372862 164212
rect 386506 164160 386512 164212
rect 386564 164200 386570 164212
rect 386690 164200 386696 164212
rect 386564 164172 386696 164200
rect 386564 164160 386570 164172
rect 386690 164160 386696 164172
rect 386748 164160 386754 164212
rect 330110 162976 330116 162988
rect 330071 162948 330116 162976
rect 330110 162936 330116 162948
rect 330168 162936 330174 162988
rect 232130 162800 232136 162852
rect 232188 162840 232194 162852
rect 232222 162840 232228 162852
rect 232188 162812 232228 162840
rect 232188 162800 232194 162812
rect 232222 162800 232228 162812
rect 232280 162800 232286 162852
rect 358538 162800 358544 162852
rect 358596 162840 358602 162852
rect 358722 162840 358728 162852
rect 358596 162812 358728 162840
rect 358596 162800 358602 162812
rect 358722 162800 358728 162812
rect 358780 162800 358786 162852
rect 421190 162840 421196 162852
rect 421151 162812 421196 162840
rect 421190 162800 421196 162812
rect 421248 162800 421254 162852
rect 357526 162732 357532 162784
rect 357584 162772 357590 162784
rect 357618 162772 357624 162784
rect 357584 162744 357624 162772
rect 357584 162732 357590 162744
rect 357618 162732 357624 162744
rect 357676 162732 357682 162784
rect 285950 161480 285956 161492
rect 285911 161452 285956 161480
rect 285950 161440 285956 161452
rect 286008 161440 286014 161492
rect 460106 161480 460112 161492
rect 460067 161452 460112 161480
rect 460106 161440 460112 161452
rect 460164 161440 460170 161492
rect 302510 161372 302516 161424
rect 302568 161412 302574 161424
rect 302602 161412 302608 161424
rect 302568 161384 302608 161412
rect 302568 161372 302574 161384
rect 302602 161372 302608 161384
rect 302660 161372 302666 161424
rect 330110 161412 330116 161424
rect 330071 161384 330116 161412
rect 330110 161372 330116 161384
rect 330168 161372 330174 161424
rect 295610 160080 295616 160132
rect 295668 160120 295674 160132
rect 295702 160120 295708 160132
rect 295668 160092 295708 160120
rect 295668 160080 295674 160092
rect 295702 160080 295708 160092
rect 295760 160080 295766 160132
rect 296898 160080 296904 160132
rect 296956 160120 296962 160132
rect 296990 160120 296996 160132
rect 296956 160092 296996 160120
rect 296956 160080 296962 160092
rect 296990 160080 296996 160092
rect 297048 160080 297054 160132
rect 306374 160012 306380 160064
rect 306432 160052 306438 160064
rect 306834 160052 306840 160064
rect 306432 160024 306840 160052
rect 306432 160012 306438 160024
rect 306834 160012 306840 160024
rect 306892 160012 306898 160064
rect 285950 158652 285956 158704
rect 286008 158692 286014 158704
rect 286045 158695 286103 158701
rect 286045 158692 286057 158695
rect 286008 158664 286057 158692
rect 286008 158652 286014 158664
rect 286045 158661 286057 158664
rect 286091 158661 286103 158695
rect 294322 158692 294328 158704
rect 294283 158664 294328 158692
rect 286045 158655 286103 158661
rect 294322 158652 294328 158664
rect 294380 158652 294386 158704
rect 272150 158012 272156 158024
rect 272111 157984 272156 158012
rect 272150 157972 272156 157984
rect 272208 157972 272214 158024
rect 337010 157972 337016 158024
rect 337068 158012 337074 158024
rect 337194 158012 337200 158024
rect 337068 157984 337200 158012
rect 337068 157972 337074 157984
rect 337194 157972 337200 157984
rect 337252 157972 337258 158024
rect 364334 157564 364340 157616
rect 364392 157604 364398 157616
rect 373810 157604 373816 157616
rect 364392 157576 373816 157604
rect 364392 157564 364398 157576
rect 373810 157564 373816 157576
rect 373868 157564 373874 157616
rect 396074 157496 396080 157548
rect 396132 157536 396138 157548
rect 400766 157536 400772 157548
rect 396132 157508 400772 157536
rect 396132 157496 396138 157508
rect 400766 157496 400772 157508
rect 400824 157496 400830 157548
rect 417878 157496 417884 157548
rect 417936 157536 417942 157548
rect 418154 157536 418160 157548
rect 417936 157508 418160 157536
rect 417936 157496 417942 157508
rect 418154 157496 418160 157508
rect 418212 157496 418218 157548
rect 437198 157496 437204 157548
rect 437256 157536 437262 157548
rect 437474 157536 437480 157548
rect 437256 157508 437480 157536
rect 437256 157496 437262 157508
rect 437474 157496 437480 157508
rect 437532 157496 437538 157548
rect 456518 157496 456524 157548
rect 456576 157536 456582 157548
rect 458266 157536 458272 157548
rect 456576 157508 458272 157536
rect 456576 157496 456582 157508
rect 458266 157496 458272 157508
rect 458324 157496 458330 157548
rect 267734 157428 267740 157480
rect 267792 157428 267798 157480
rect 265158 157360 265164 157412
rect 265216 157360 265222 157412
rect 265176 157264 265204 157360
rect 267752 157344 267780 157428
rect 325878 157360 325884 157412
rect 325936 157360 325942 157412
rect 327166 157360 327172 157412
rect 327224 157360 327230 157412
rect 267734 157292 267740 157344
rect 267792 157292 267798 157344
rect 265250 157264 265256 157276
rect 265176 157236 265256 157264
rect 265250 157224 265256 157236
rect 265308 157224 265314 157276
rect 325896 157196 325924 157360
rect 327184 157264 327212 157360
rect 359090 157292 359096 157344
rect 359148 157292 359154 157344
rect 372798 157332 372804 157344
rect 372759 157304 372804 157332
rect 372798 157292 372804 157304
rect 372856 157292 372862 157344
rect 377122 157292 377128 157344
rect 377180 157292 377186 157344
rect 327258 157264 327264 157276
rect 327184 157236 327264 157264
rect 327258 157224 327264 157236
rect 327316 157224 327322 157276
rect 359108 157264 359136 157292
rect 359182 157264 359188 157276
rect 359108 157236 359188 157264
rect 359182 157224 359188 157236
rect 359240 157224 359246 157276
rect 377140 157264 377168 157292
rect 377214 157264 377220 157276
rect 377140 157236 377220 157264
rect 377214 157224 377220 157236
rect 377272 157224 377278 157276
rect 325970 157196 325976 157208
rect 325896 157168 325976 157196
rect 325970 157156 325976 157168
rect 326028 157156 326034 157208
rect 247218 154572 247224 154624
rect 247276 154612 247282 154624
rect 247310 154612 247316 154624
rect 247276 154584 247316 154612
rect 247276 154572 247282 154584
rect 247310 154572 247316 154584
rect 247368 154572 247374 154624
rect 299750 154504 299756 154556
rect 299808 154544 299814 154556
rect 299842 154544 299848 154556
rect 299808 154516 299848 154544
rect 299808 154504 299814 154516
rect 299842 154504 299848 154516
rect 299900 154504 299906 154556
rect 470410 154504 470416 154556
rect 470468 154544 470474 154556
rect 470594 154544 470600 154556
rect 470468 154516 470600 154544
rect 470468 154504 470474 154516
rect 470594 154504 470600 154516
rect 470652 154504 470658 154556
rect 301038 154436 301044 154488
rect 301096 154476 301102 154488
rect 301222 154476 301228 154488
rect 301096 154448 301228 154476
rect 301096 154436 301102 154448
rect 301222 154436 301228 154448
rect 301280 154436 301286 154488
rect 259641 154207 259699 154213
rect 259641 154173 259653 154207
rect 259687 154204 259699 154207
rect 259822 154204 259828 154216
rect 259687 154176 259828 154204
rect 259687 154173 259699 154176
rect 259641 154167 259699 154173
rect 259822 154164 259828 154176
rect 259880 154164 259886 154216
rect 421190 153252 421196 153264
rect 421151 153224 421196 153252
rect 421190 153212 421196 153224
rect 421248 153212 421254 153264
rect 289998 153144 290004 153196
rect 290056 153184 290062 153196
rect 290090 153184 290096 153196
rect 290056 153156 290096 153184
rect 290056 153144 290062 153156
rect 290090 153144 290096 153156
rect 290148 153144 290154 153196
rect 291470 153144 291476 153196
rect 291528 153184 291534 153196
rect 291562 153184 291568 153196
rect 291528 153156 291568 153184
rect 291528 153144 291534 153156
rect 291562 153144 291568 153156
rect 291620 153144 291626 153196
rect 295518 153144 295524 153196
rect 295576 153184 295582 153196
rect 295610 153184 295616 153196
rect 295576 153156 295616 153184
rect 295576 153144 295582 153156
rect 295610 153144 295616 153156
rect 295668 153144 295674 153196
rect 310790 153184 310796 153196
rect 310751 153156 310796 153184
rect 310790 153144 310796 153156
rect 310848 153144 310854 153196
rect 341150 153184 341156 153196
rect 341111 153156 341156 153184
rect 341150 153144 341156 153156
rect 341208 153144 341214 153196
rect 330110 151824 330116 151836
rect 330071 151796 330116 151824
rect 330110 151784 330116 151796
rect 330168 151784 330174 151836
rect 3326 151716 3332 151768
rect 3384 151756 3390 151768
rect 17218 151756 17224 151768
rect 3384 151728 17224 151756
rect 3384 151716 3390 151728
rect 17218 151716 17224 151728
rect 17276 151716 17282 151768
rect 460106 151756 460112 151768
rect 460067 151728 460112 151756
rect 460106 151716 460112 151728
rect 460164 151716 460170 151768
rect 339494 149676 339500 149728
rect 339552 149716 339558 149728
rect 339770 149716 339776 149728
rect 339552 149688 339776 149716
rect 339552 149676 339558 149688
rect 339770 149676 339776 149688
rect 339828 149676 339834 149728
rect 294322 149104 294328 149116
rect 294283 149076 294328 149104
rect 294322 149064 294328 149076
rect 294380 149064 294386 149116
rect 272150 148968 272156 148980
rect 272111 148940 272156 148968
rect 272150 148928 272156 148940
rect 272208 148928 272214 148980
rect 360197 147747 360255 147753
rect 360197 147713 360209 147747
rect 360243 147744 360255 147747
rect 360378 147744 360384 147756
rect 360243 147716 360384 147744
rect 360243 147713 360255 147716
rect 360197 147707 360255 147713
rect 360378 147704 360384 147716
rect 360436 147704 360442 147756
rect 463697 147747 463755 147753
rect 463697 147713 463709 147747
rect 463743 147744 463755 147747
rect 463786 147744 463792 147756
rect 463743 147716 463792 147744
rect 463743 147713 463755 147716
rect 463697 147707 463755 147713
rect 463786 147704 463792 147716
rect 463844 147704 463850 147756
rect 330110 147636 330116 147688
rect 330168 147636 330174 147688
rect 310790 147608 310796 147620
rect 310751 147580 310796 147608
rect 310790 147568 310796 147580
rect 310848 147568 310854 147620
rect 330128 147608 330156 147636
rect 330202 147608 330208 147620
rect 330128 147580 330208 147608
rect 330202 147568 330208 147580
rect 330260 147568 330266 147620
rect 266722 144916 266728 144968
rect 266780 144916 266786 144968
rect 463694 144916 463700 144968
rect 463752 144956 463758 144968
rect 463752 144928 463797 144956
rect 463752 144916 463758 144928
rect 244274 144848 244280 144900
rect 244332 144888 244338 144900
rect 244458 144888 244464 144900
rect 244332 144860 244464 144888
rect 244332 144848 244338 144860
rect 244458 144848 244464 144860
rect 244516 144848 244522 144900
rect 247126 144848 247132 144900
rect 247184 144888 247190 144900
rect 247218 144888 247224 144900
rect 247184 144860 247224 144888
rect 247184 144848 247190 144860
rect 247218 144848 247224 144860
rect 247276 144848 247282 144900
rect 262582 144848 262588 144900
rect 262640 144888 262646 144900
rect 262766 144888 262772 144900
rect 262640 144860 262772 144888
rect 262640 144848 262646 144860
rect 262766 144848 262772 144860
rect 262824 144848 262830 144900
rect 266740 144832 266768 144916
rect 267734 144848 267740 144900
rect 267792 144888 267798 144900
rect 267918 144888 267924 144900
rect 267792 144860 267924 144888
rect 267792 144848 267798 144860
rect 267918 144848 267924 144860
rect 267976 144848 267982 144900
rect 270678 144888 270684 144900
rect 270639 144860 270684 144888
rect 270678 144848 270684 144860
rect 270736 144848 270742 144900
rect 272150 144848 272156 144900
rect 272208 144888 272214 144900
rect 272426 144888 272432 144900
rect 272208 144860 272432 144888
rect 272208 144848 272214 144860
rect 272426 144848 272432 144860
rect 272484 144848 272490 144900
rect 323302 144848 323308 144900
rect 323360 144888 323366 144900
rect 323394 144888 323400 144900
rect 323360 144860 323400 144888
rect 323360 144848 323366 144860
rect 323394 144848 323400 144860
rect 323452 144848 323458 144900
rect 325878 144848 325884 144900
rect 325936 144888 325942 144900
rect 326062 144888 326068 144900
rect 325936 144860 326068 144888
rect 325936 144848 325942 144860
rect 326062 144848 326068 144860
rect 326120 144848 326126 144900
rect 327166 144848 327172 144900
rect 327224 144888 327230 144900
rect 327350 144888 327356 144900
rect 327224 144860 327356 144888
rect 327224 144848 327230 144860
rect 327350 144848 327356 144860
rect 327408 144848 327414 144900
rect 341153 144891 341211 144897
rect 341153 144857 341165 144891
rect 341199 144888 341211 144891
rect 341334 144888 341340 144900
rect 341199 144860 341340 144888
rect 341199 144857 341211 144860
rect 341153 144851 341211 144857
rect 341334 144848 341340 144860
rect 341392 144848 341398 144900
rect 360194 144888 360200 144900
rect 360155 144860 360200 144888
rect 360194 144848 360200 144860
rect 360252 144848 360258 144900
rect 367002 144888 367008 144900
rect 366963 144860 367008 144888
rect 367002 144848 367008 144860
rect 367060 144848 367066 144900
rect 386506 144848 386512 144900
rect 386564 144888 386570 144900
rect 386690 144888 386696 144900
rect 386564 144860 386696 144888
rect 386564 144848 386570 144860
rect 386690 144848 386696 144860
rect 386748 144848 386754 144900
rect 266722 144780 266728 144832
rect 266780 144780 266786 144832
rect 339678 144780 339684 144832
rect 339736 144820 339742 144832
rect 339862 144820 339868 144832
rect 339736 144792 339868 144820
rect 339736 144780 339742 144792
rect 339862 144780 339868 144792
rect 339920 144780 339926 144832
rect 232314 143528 232320 143540
rect 232275 143500 232320 143528
rect 232314 143488 232320 143500
rect 232372 143488 232378 143540
rect 272426 143528 272432 143540
rect 272387 143500 272432 143528
rect 272426 143488 272432 143500
rect 272484 143488 272490 143540
rect 301038 143488 301044 143540
rect 301096 143528 301102 143540
rect 301222 143528 301228 143540
rect 301096 143500 301228 143528
rect 301096 143488 301102 143500
rect 301222 143488 301228 143500
rect 301280 143488 301286 143540
rect 323302 143528 323308 143540
rect 323263 143500 323308 143528
rect 323302 143488 323308 143500
rect 323360 143488 323366 143540
rect 324590 143528 324596 143540
rect 324551 143500 324596 143528
rect 324590 143488 324596 143500
rect 324648 143488 324654 143540
rect 330113 143531 330171 143537
rect 330113 143497 330125 143531
rect 330159 143528 330171 143531
rect 330202 143528 330208 143540
rect 330159 143500 330208 143528
rect 330159 143497 330171 143500
rect 330113 143491 330171 143497
rect 330202 143488 330208 143500
rect 330260 143488 330266 143540
rect 421190 143528 421196 143540
rect 421151 143500 421196 143528
rect 421190 143488 421196 143500
rect 421248 143488 421254 143540
rect 460106 142236 460112 142248
rect 460067 142208 460112 142236
rect 460106 142196 460112 142208
rect 460164 142196 460170 142248
rect 259638 142168 259644 142180
rect 259599 142140 259644 142168
rect 259638 142128 259644 142140
rect 259696 142128 259702 142180
rect 306374 142128 306380 142180
rect 306432 142168 306438 142180
rect 307018 142168 307024 142180
rect 306432 142140 307024 142168
rect 306432 142128 306438 142140
rect 307018 142128 307024 142140
rect 307076 142128 307082 142180
rect 317506 142128 317512 142180
rect 317564 142168 317570 142180
rect 317690 142168 317696 142180
rect 317564 142140 317696 142168
rect 317564 142128 317570 142140
rect 317690 142128 317696 142140
rect 317748 142128 317754 142180
rect 460106 142100 460112 142112
rect 460067 142072 460112 142100
rect 460106 142060 460112 142072
rect 460164 142060 460170 142112
rect 259730 141992 259736 142044
rect 259788 142032 259794 142044
rect 259825 142035 259883 142041
rect 259825 142032 259837 142035
rect 259788 142004 259837 142032
rect 259788 141992 259794 142004
rect 259825 142001 259837 142004
rect 259871 142001 259883 142035
rect 259825 141995 259883 142001
rect 286042 140808 286048 140820
rect 286003 140780 286048 140808
rect 286042 140768 286048 140780
rect 286100 140768 286106 140820
rect 288621 140743 288679 140749
rect 288621 140709 288633 140743
rect 288667 140740 288679 140743
rect 288802 140740 288808 140752
rect 288667 140712 288808 140740
rect 288667 140709 288679 140712
rect 288621 140703 288679 140709
rect 288802 140700 288808 140712
rect 288860 140700 288866 140752
rect 294230 140700 294236 140752
rect 294288 140740 294294 140752
rect 294414 140740 294420 140752
rect 294288 140712 294420 140740
rect 294288 140700 294294 140712
rect 294414 140700 294420 140712
rect 294472 140700 294478 140752
rect 295518 140740 295524 140752
rect 295479 140712 295524 140740
rect 295518 140700 295524 140712
rect 295576 140700 295582 140752
rect 377125 140063 377183 140069
rect 377125 140029 377137 140063
rect 377171 140060 377183 140063
rect 377214 140060 377220 140072
rect 377171 140032 377220 140060
rect 377171 140029 377183 140032
rect 377125 140023 377183 140029
rect 377214 140020 377220 140032
rect 377272 140020 377278 140072
rect 270678 139992 270684 140004
rect 270639 139964 270684 139992
rect 270678 139952 270684 139964
rect 270736 139952 270742 140004
rect 294414 139380 294420 139392
rect 294375 139352 294420 139380
rect 294414 139340 294420 139352
rect 294472 139340 294478 139392
rect 372709 138159 372767 138165
rect 372709 138125 372721 138159
rect 372755 138156 372767 138159
rect 372798 138156 372804 138168
rect 372755 138128 372804 138156
rect 372755 138125 372767 138128
rect 372709 138119 372767 138125
rect 372798 138116 372804 138128
rect 372856 138116 372862 138168
rect 289909 138091 289967 138097
rect 289909 138057 289921 138091
rect 289955 138088 289967 138091
rect 290090 138088 290096 138100
rect 289955 138060 290096 138088
rect 289955 138057 289967 138060
rect 289909 138051 289967 138057
rect 290090 138048 290096 138060
rect 290148 138048 290154 138100
rect 375742 138088 375748 138100
rect 375668 138060 375748 138088
rect 375668 138032 375696 138060
rect 375742 138048 375748 138060
rect 375800 138048 375806 138100
rect 239122 137980 239128 138032
rect 239180 137980 239186 138032
rect 296806 137980 296812 138032
rect 296864 138020 296870 138032
rect 297266 138020 297272 138032
rect 296864 137992 297272 138020
rect 296864 137980 296870 137992
rect 297266 137980 297272 137992
rect 297324 137980 297330 138032
rect 337102 137980 337108 138032
rect 337160 137980 337166 138032
rect 375650 137980 375656 138032
rect 375708 137980 375714 138032
rect 463694 137980 463700 138032
rect 463752 137980 463758 138032
rect 239030 137912 239036 137964
rect 239088 137952 239094 137964
rect 239140 137952 239168 137980
rect 239088 137924 239168 137952
rect 239088 137912 239094 137924
rect 317506 137912 317512 137964
rect 317564 137952 317570 137964
rect 317782 137952 317788 137964
rect 317564 137924 317788 137952
rect 317564 137912 317570 137924
rect 317782 137912 317788 137924
rect 317840 137912 317846 137964
rect 330110 137952 330116 137964
rect 330071 137924 330116 137952
rect 330110 137912 330116 137924
rect 330168 137912 330174 137964
rect 337120 137952 337148 137980
rect 337194 137952 337200 137964
rect 337120 137924 337200 137952
rect 337194 137912 337200 137924
rect 337252 137912 337258 137964
rect 463712 137952 463740 137980
rect 463878 137952 463884 137964
rect 463712 137924 463884 137952
rect 463878 137912 463884 137924
rect 463936 137912 463942 137964
rect 2774 136484 2780 136536
rect 2832 136524 2838 136536
rect 5074 136524 5080 136536
rect 2832 136496 5080 136524
rect 2832 136484 2838 136496
rect 5074 136484 5080 136496
rect 5132 136484 5138 136536
rect 367002 135300 367008 135312
rect 366963 135272 367008 135300
rect 367002 135260 367008 135272
rect 367060 135260 367066 135312
rect 372706 135300 372712 135312
rect 372667 135272 372712 135300
rect 372706 135260 372712 135272
rect 372764 135260 372770 135312
rect 377122 135300 377128 135312
rect 377083 135272 377128 135300
rect 377122 135260 377128 135272
rect 377180 135260 377186 135312
rect 266630 135192 266636 135244
rect 266688 135232 266694 135244
rect 266722 135232 266728 135244
rect 266688 135204 266728 135232
rect 266688 135192 266694 135204
rect 266722 135192 266728 135204
rect 266780 135192 266786 135244
rect 272426 135232 272432 135244
rect 272387 135204 272432 135232
rect 272426 135192 272432 135204
rect 272484 135192 272490 135244
rect 358722 135232 358728 135244
rect 358683 135204 358728 135232
rect 358722 135192 358728 135204
rect 358780 135192 358786 135244
rect 470410 135192 470416 135244
rect 470468 135232 470474 135244
rect 470594 135232 470600 135244
rect 470468 135204 470600 135232
rect 470468 135192 470474 135204
rect 470594 135192 470600 135204
rect 470652 135192 470658 135244
rect 232314 133940 232320 133952
rect 232275 133912 232320 133940
rect 232314 133900 232320 133912
rect 232372 133900 232378 133952
rect 307018 133900 307024 133952
rect 307076 133900 307082 133952
rect 323302 133940 323308 133952
rect 323263 133912 323308 133940
rect 323302 133900 323308 133912
rect 323360 133900 323366 133952
rect 421190 133940 421196 133952
rect 421151 133912 421196 133940
rect 421190 133900 421196 133912
rect 421248 133900 421254 133952
rect 265250 133872 265256 133884
rect 265211 133844 265256 133872
rect 265250 133832 265256 133844
rect 265308 133832 265314 133884
rect 307036 133816 307064 133900
rect 307018 133764 307024 133816
rect 307076 133764 307082 133816
rect 324593 132515 324651 132521
rect 324593 132481 324605 132515
rect 324639 132512 324651 132515
rect 324682 132512 324688 132524
rect 324639 132484 324688 132512
rect 324639 132481 324651 132484
rect 324593 132475 324651 132481
rect 324682 132472 324688 132484
rect 324740 132472 324746 132524
rect 460109 132515 460167 132521
rect 460109 132481 460121 132515
rect 460155 132512 460167 132515
rect 460198 132512 460204 132524
rect 460155 132484 460204 132512
rect 460155 132481 460167 132484
rect 460109 132475 460167 132481
rect 460198 132472 460204 132484
rect 460256 132472 460262 132524
rect 463694 132472 463700 132524
rect 463752 132512 463758 132524
rect 463878 132512 463884 132524
rect 463752 132484 463884 132512
rect 463752 132472 463758 132484
rect 463878 132472 463884 132484
rect 463936 132472 463942 132524
rect 289906 132444 289912 132456
rect 289867 132416 289912 132444
rect 289906 132404 289912 132416
rect 289964 132404 289970 132456
rect 337194 132444 337200 132456
rect 337155 132416 337200 132444
rect 337194 132404 337200 132416
rect 337252 132404 337258 132456
rect 288618 131152 288624 131164
rect 288579 131124 288624 131152
rect 288618 131112 288624 131124
rect 288676 131112 288682 131164
rect 295521 131155 295579 131161
rect 295521 131121 295533 131155
rect 295567 131152 295579 131155
rect 295610 131152 295616 131164
rect 295567 131124 295616 131152
rect 295567 131121 295579 131124
rect 295521 131115 295579 131121
rect 295610 131112 295616 131124
rect 295668 131112 295674 131164
rect 291470 131084 291476 131096
rect 291431 131056 291476 131084
rect 291470 131044 291476 131056
rect 291528 131044 291534 131096
rect 296901 131087 296959 131093
rect 296901 131053 296913 131087
rect 296947 131084 296959 131087
rect 297174 131084 297180 131096
rect 296947 131056 297180 131084
rect 296947 131053 296959 131056
rect 296901 131047 296959 131053
rect 297174 131044 297180 131056
rect 297232 131044 297238 131096
rect 270494 130364 270500 130416
rect 270552 130404 270558 130416
rect 270678 130404 270684 130416
rect 270552 130376 270684 130404
rect 270552 130364 270558 130376
rect 270678 130364 270684 130376
rect 270736 130364 270742 130416
rect 294414 129792 294420 129804
rect 294375 129764 294420 129792
rect 294414 129752 294420 129764
rect 294472 129752 294478 129804
rect 325970 128432 325976 128444
rect 325896 128404 325976 128432
rect 250070 128324 250076 128376
rect 250128 128324 250134 128376
rect 284662 128324 284668 128376
rect 284720 128324 284726 128376
rect 302602 128324 302608 128376
rect 302660 128324 302666 128376
rect 250088 128296 250116 128324
rect 250162 128296 250168 128308
rect 250088 128268 250168 128296
rect 250162 128256 250168 128268
rect 250220 128256 250226 128308
rect 284680 128296 284708 128324
rect 284754 128296 284760 128308
rect 284680 128268 284760 128296
rect 284754 128256 284760 128268
rect 284812 128256 284818 128308
rect 302620 128240 302648 128324
rect 325896 128308 325924 128404
rect 325970 128392 325976 128404
rect 326028 128392 326034 128444
rect 327258 128432 327264 128444
rect 327184 128404 327264 128432
rect 327184 128308 327212 128404
rect 327258 128392 327264 128404
rect 327316 128392 327322 128444
rect 341242 128392 341248 128444
rect 341300 128392 341306 128444
rect 339678 128324 339684 128376
rect 339736 128364 339742 128376
rect 339862 128364 339868 128376
rect 339736 128336 339868 128364
rect 339736 128324 339742 128336
rect 339862 128324 339868 128336
rect 339920 128324 339926 128376
rect 341260 128308 341288 128392
rect 325878 128256 325884 128308
rect 325936 128256 325942 128308
rect 327166 128256 327172 128308
rect 327224 128256 327230 128308
rect 341242 128256 341248 128308
rect 341300 128256 341306 128308
rect 302602 128188 302608 128240
rect 302660 128188 302666 128240
rect 272150 125808 272156 125860
rect 272208 125848 272214 125860
rect 272426 125848 272432 125860
rect 272208 125820 272432 125848
rect 272208 125808 272214 125820
rect 272426 125808 272432 125820
rect 272484 125808 272490 125860
rect 358722 125644 358728 125656
rect 358683 125616 358728 125644
rect 358722 125604 358728 125616
rect 358780 125604 358786 125656
rect 239122 125576 239128 125588
rect 239083 125548 239128 125576
rect 239122 125536 239128 125548
rect 239180 125536 239186 125588
rect 251450 125576 251456 125588
rect 251411 125548 251456 125576
rect 251450 125536 251456 125548
rect 251508 125536 251514 125588
rect 262582 125536 262588 125588
rect 262640 125576 262646 125588
rect 262766 125576 262772 125588
rect 262640 125548 262772 125576
rect 262640 125536 262646 125548
rect 262766 125536 262772 125548
rect 262824 125536 262830 125588
rect 267734 125536 267740 125588
rect 267792 125576 267798 125588
rect 267918 125576 267924 125588
rect 267792 125548 267924 125576
rect 267792 125536 267798 125548
rect 267918 125536 267924 125548
rect 267976 125536 267982 125588
rect 270678 125576 270684 125588
rect 270639 125548 270684 125576
rect 270678 125536 270684 125548
rect 270736 125536 270742 125588
rect 272150 125536 272156 125588
rect 272208 125576 272214 125588
rect 272426 125576 272432 125588
rect 272208 125548 272432 125576
rect 272208 125536 272214 125548
rect 272426 125536 272432 125548
rect 272484 125536 272490 125588
rect 317690 125536 317696 125588
rect 317748 125576 317754 125588
rect 317966 125576 317972 125588
rect 317748 125548 317972 125576
rect 317748 125536 317754 125548
rect 317966 125536 317972 125548
rect 318024 125536 318030 125588
rect 325878 125536 325884 125588
rect 325936 125576 325942 125588
rect 326062 125576 326068 125588
rect 325936 125548 326068 125576
rect 325936 125536 325942 125548
rect 326062 125536 326068 125548
rect 326120 125536 326126 125588
rect 327166 125536 327172 125588
rect 327224 125576 327230 125588
rect 327350 125576 327356 125588
rect 327224 125548 327356 125576
rect 327224 125536 327230 125548
rect 327350 125536 327356 125548
rect 327408 125536 327414 125588
rect 336734 125536 336740 125588
rect 336792 125576 336798 125588
rect 336918 125576 336924 125588
rect 336792 125548 336924 125576
rect 336792 125536 336798 125548
rect 336918 125536 336924 125548
rect 336976 125536 336982 125588
rect 339770 125576 339776 125588
rect 339731 125548 339776 125576
rect 339770 125536 339776 125548
rect 339828 125536 339834 125588
rect 341153 125579 341211 125585
rect 341153 125545 341165 125579
rect 341199 125576 341211 125579
rect 341242 125576 341248 125588
rect 341199 125548 341248 125576
rect 341199 125545 341211 125548
rect 341153 125539 341211 125545
rect 341242 125536 341248 125548
rect 341300 125536 341306 125588
rect 259822 124216 259828 124228
rect 259783 124188 259828 124216
rect 259822 124176 259828 124188
rect 259880 124176 259886 124228
rect 265250 124216 265256 124228
rect 265211 124188 265256 124216
rect 265250 124176 265256 124188
rect 265308 124176 265314 124228
rect 360194 124176 360200 124228
rect 360252 124216 360258 124228
rect 360378 124216 360384 124228
rect 360252 124188 360384 124216
rect 360252 124176 360258 124188
rect 360378 124176 360384 124188
rect 360436 124176 360442 124228
rect 232314 124148 232320 124160
rect 232275 124120 232320 124148
rect 232314 124108 232320 124120
rect 232372 124108 232378 124160
rect 249981 124151 250039 124157
rect 249981 124117 249993 124151
rect 250027 124148 250039 124151
rect 250162 124148 250168 124160
rect 250027 124120 250168 124148
rect 250027 124117 250039 124120
rect 249981 124111 250039 124117
rect 250162 124108 250168 124120
rect 250220 124108 250226 124160
rect 272426 124148 272432 124160
rect 272387 124120 272432 124148
rect 272426 124108 272432 124120
rect 272484 124108 272490 124160
rect 299842 124148 299848 124160
rect 299803 124120 299848 124148
rect 299842 124108 299848 124120
rect 299900 124108 299906 124160
rect 306834 124148 306840 124160
rect 306795 124120 306840 124148
rect 306834 124108 306840 124120
rect 306892 124108 306898 124160
rect 359090 124108 359096 124160
rect 359148 124148 359154 124160
rect 359182 124148 359188 124160
rect 359148 124120 359188 124148
rect 359148 124108 359154 124120
rect 359182 124108 359188 124120
rect 359240 124108 359246 124160
rect 421190 124148 421196 124160
rect 421151 124120 421196 124148
rect 421190 124108 421196 124120
rect 421248 124108 421254 124160
rect 460014 124040 460020 124092
rect 460072 124080 460078 124092
rect 460198 124080 460204 124092
rect 460072 124052 460204 124080
rect 460072 124040 460078 124052
rect 460198 124040 460204 124052
rect 460256 124040 460262 124092
rect 284754 122748 284760 122800
rect 284812 122748 284818 122800
rect 324682 122788 324688 122800
rect 324643 122760 324688 122788
rect 324682 122748 324688 122760
rect 324740 122748 324746 122800
rect 284772 122664 284800 122748
rect 291473 122723 291531 122729
rect 291473 122689 291485 122723
rect 291519 122720 291531 122723
rect 291562 122720 291568 122732
rect 291519 122692 291568 122720
rect 291519 122689 291531 122692
rect 291473 122683 291531 122689
rect 291562 122680 291568 122692
rect 291620 122680 291626 122732
rect 284754 122612 284760 122664
rect 284812 122612 284818 122664
rect 2774 122272 2780 122324
rect 2832 122312 2838 122324
rect 4982 122312 4988 122324
rect 2832 122284 4988 122312
rect 2832 122272 2838 122284
rect 4982 122272 4988 122284
rect 5040 122272 5046 122324
rect 288618 121456 288624 121508
rect 288676 121496 288682 121508
rect 288894 121496 288900 121508
rect 288676 121468 288900 121496
rect 288676 121456 288682 121468
rect 288894 121456 288900 121468
rect 288952 121456 288958 121508
rect 294322 121456 294328 121508
rect 294380 121496 294386 121508
rect 294414 121496 294420 121508
rect 294380 121468 294420 121496
rect 294380 121456 294386 121468
rect 294414 121456 294420 121468
rect 294472 121456 294478 121508
rect 296898 121496 296904 121508
rect 296859 121468 296904 121496
rect 296898 121456 296904 121468
rect 296956 121456 296962 121508
rect 270678 120680 270684 120692
rect 270639 120652 270684 120680
rect 270678 120640 270684 120652
rect 270736 120640 270742 120692
rect 273530 118668 273536 118720
rect 273588 118668 273594 118720
rect 372706 118668 372712 118720
rect 372764 118668 372770 118720
rect 377122 118668 377128 118720
rect 377180 118668 377186 118720
rect 273548 118640 273576 118668
rect 273622 118640 273628 118652
rect 273548 118612 273628 118640
rect 273622 118600 273628 118612
rect 273680 118600 273686 118652
rect 339770 118640 339776 118652
rect 339731 118612 339776 118640
rect 339770 118600 339776 118612
rect 339828 118600 339834 118652
rect 341150 118640 341156 118652
rect 341111 118612 341156 118640
rect 341150 118600 341156 118612
rect 341208 118600 341214 118652
rect 372724 118584 372752 118668
rect 377140 118584 377168 118668
rect 372706 118532 372712 118584
rect 372764 118532 372770 118584
rect 377122 118532 377128 118584
rect 377180 118532 377186 118584
rect 327258 118464 327264 118516
rect 327316 118504 327322 118516
rect 327350 118504 327356 118516
rect 327316 118476 327356 118504
rect 327316 118464 327322 118476
rect 327350 118464 327356 118476
rect 327408 118464 327414 118516
rect 262582 117988 262588 118040
rect 262640 118028 262646 118040
rect 262766 118028 262772 118040
rect 262640 118000 262772 118028
rect 262640 117988 262646 118000
rect 262766 117988 262772 118000
rect 262824 117988 262830 118040
rect 239122 115988 239128 116000
rect 239083 115960 239128 115988
rect 239122 115948 239128 115960
rect 239180 115948 239186 116000
rect 251450 115988 251456 116000
rect 251411 115960 251456 115988
rect 251450 115948 251456 115960
rect 251508 115948 251514 116000
rect 341153 115923 341211 115929
rect 341153 115889 341165 115923
rect 341199 115920 341211 115923
rect 341242 115920 341248 115932
rect 341199 115892 341248 115920
rect 341199 115889 341211 115892
rect 341153 115883 341211 115889
rect 341242 115880 341248 115892
rect 341300 115880 341306 115932
rect 367002 115920 367008 115932
rect 366963 115892 367008 115920
rect 367002 115880 367008 115892
rect 367060 115880 367066 115932
rect 376938 115880 376944 115932
rect 376996 115920 377002 115932
rect 377122 115920 377128 115932
rect 376996 115892 377128 115920
rect 376996 115880 377002 115892
rect 377122 115880 377128 115892
rect 377180 115880 377186 115932
rect 470594 115920 470600 115932
rect 470555 115892 470600 115920
rect 470594 115880 470600 115892
rect 470652 115880 470658 115932
rect 259822 115404 259828 115456
rect 259880 115404 259886 115456
rect 259840 115320 259868 115404
rect 259822 115268 259828 115320
rect 259880 115268 259886 115320
rect 296898 114628 296904 114640
rect 296824 114600 296904 114628
rect 232314 114560 232320 114572
rect 232275 114532 232320 114560
rect 232314 114520 232320 114532
rect 232372 114520 232378 114572
rect 249978 114560 249984 114572
rect 249939 114532 249984 114560
rect 249978 114520 249984 114532
rect 250036 114520 250042 114572
rect 272426 114560 272432 114572
rect 272387 114532 272432 114560
rect 272426 114520 272432 114532
rect 272484 114520 272490 114572
rect 296824 114504 296852 114600
rect 296898 114588 296904 114600
rect 296956 114588 296962 114640
rect 357526 114628 357532 114640
rect 357452 114600 357532 114628
rect 357452 114572 357480 114600
rect 357526 114588 357532 114600
rect 357584 114588 357590 114640
rect 299842 114560 299848 114572
rect 299803 114532 299848 114560
rect 299842 114520 299848 114532
rect 299900 114520 299906 114572
rect 337194 114560 337200 114572
rect 337155 114532 337200 114560
rect 337194 114520 337200 114532
rect 337252 114520 337258 114572
rect 357434 114520 357440 114572
rect 357492 114520 357498 114572
rect 358630 114520 358636 114572
rect 358688 114560 358694 114572
rect 358722 114560 358728 114572
rect 358688 114532 358728 114560
rect 358688 114520 358694 114532
rect 358722 114520 358728 114532
rect 358780 114520 358786 114572
rect 421190 114560 421196 114572
rect 421151 114532 421196 114560
rect 421190 114520 421196 114532
rect 421248 114520 421254 114572
rect 296806 114452 296812 114504
rect 296864 114452 296870 114504
rect 327169 114495 327227 114501
rect 327169 114461 327181 114495
rect 327215 114492 327227 114495
rect 327258 114492 327264 114504
rect 327215 114464 327264 114492
rect 327215 114461 327227 114464
rect 327169 114455 327227 114461
rect 327258 114452 327264 114464
rect 327316 114452 327322 114504
rect 306742 113228 306748 113280
rect 306800 113268 306806 113280
rect 306837 113271 306895 113277
rect 306837 113268 306849 113271
rect 306800 113240 306849 113268
rect 306800 113228 306806 113240
rect 306837 113237 306849 113240
rect 306883 113237 306895 113271
rect 306837 113231 306895 113237
rect 286042 113160 286048 113212
rect 286100 113200 286106 113212
rect 286226 113200 286232 113212
rect 286100 113172 286232 113200
rect 286100 113160 286106 113172
rect 286226 113160 286232 113172
rect 286284 113160 286290 113212
rect 324682 113200 324688 113212
rect 324643 113172 324688 113200
rect 324682 113160 324688 113172
rect 324740 113160 324746 113212
rect 265250 113132 265256 113144
rect 265211 113104 265256 113132
rect 265250 113092 265256 113104
rect 265308 113092 265314 113144
rect 284662 113132 284668 113144
rect 284623 113104 284668 113132
rect 284662 113092 284668 113104
rect 284720 113092 284726 113144
rect 291562 113132 291568 113144
rect 291523 113104 291568 113132
rect 291562 113092 291568 113104
rect 291620 113092 291626 113144
rect 296806 113132 296812 113144
rect 296767 113104 296812 113132
rect 296806 113092 296812 113104
rect 296864 113092 296870 113144
rect 306834 113092 306840 113144
rect 306892 113132 306898 113144
rect 307018 113132 307024 113144
rect 306892 113104 307024 113132
rect 306892 113092 306898 113104
rect 307018 113092 307024 113104
rect 307076 113092 307082 113144
rect 329926 113092 329932 113144
rect 329984 113132 329990 113144
rect 330202 113132 330208 113144
rect 329984 113104 330208 113132
rect 329984 113092 329990 113104
rect 330202 113092 330208 113104
rect 330260 113092 330266 113144
rect 286042 113024 286048 113076
rect 286100 113064 286106 113076
rect 286226 113064 286232 113076
rect 286100 113036 286232 113064
rect 286100 113024 286106 113036
rect 286226 113024 286232 113036
rect 286284 113024 286290 113076
rect 270678 111052 270684 111104
rect 270736 111092 270742 111104
rect 270862 111092 270868 111104
rect 270736 111064 270868 111092
rect 270736 111052 270742 111064
rect 270862 111052 270868 111064
rect 270920 111052 270926 111104
rect 463878 111052 463884 111104
rect 463936 111092 463942 111104
rect 464062 111092 464068 111104
rect 463936 111064 464068 111092
rect 463936 111052 463942 111064
rect 464062 111052 464068 111064
rect 464120 111052 464126 111104
rect 294322 109732 294328 109744
rect 294283 109704 294328 109732
rect 294322 109692 294328 109704
rect 294380 109692 294386 109744
rect 247218 109052 247224 109064
rect 247179 109024 247224 109052
rect 247218 109012 247224 109024
rect 247276 109012 247282 109064
rect 310790 109012 310796 109064
rect 310848 109012 310854 109064
rect 375650 109012 375656 109064
rect 375708 109012 375714 109064
rect 310808 108984 310836 109012
rect 310882 108984 310888 108996
rect 310808 108956 310888 108984
rect 310882 108944 310888 108956
rect 310940 108944 310946 108996
rect 375558 108944 375564 108996
rect 375616 108984 375622 108996
rect 375668 108984 375696 109012
rect 375616 108956 375696 108984
rect 375616 108944 375622 108956
rect 272150 106496 272156 106548
rect 272208 106536 272214 106548
rect 272426 106536 272432 106548
rect 272208 106508 272432 106536
rect 272208 106496 272214 106508
rect 272426 106496 272432 106508
rect 272484 106496 272490 106548
rect 247218 106332 247224 106344
rect 247179 106304 247224 106332
rect 247218 106292 247224 106304
rect 247276 106292 247282 106344
rect 325970 106332 325976 106344
rect 325931 106304 325976 106332
rect 325970 106292 325976 106304
rect 326028 106292 326034 106344
rect 341150 106332 341156 106344
rect 341111 106304 341156 106332
rect 341150 106292 341156 106304
rect 341208 106292 341214 106344
rect 358630 106292 358636 106344
rect 358688 106292 358694 106344
rect 367002 106332 367008 106344
rect 366963 106304 367008 106332
rect 367002 106292 367008 106304
rect 367060 106292 367066 106344
rect 470594 106332 470600 106344
rect 470555 106304 470600 106332
rect 470594 106292 470600 106304
rect 470652 106292 470658 106344
rect 236454 106224 236460 106276
rect 236512 106264 236518 106276
rect 236638 106264 236644 106276
rect 236512 106236 236644 106264
rect 236512 106224 236518 106236
rect 236638 106224 236644 106236
rect 236696 106224 236702 106276
rect 239122 106224 239128 106276
rect 239180 106264 239186 106276
rect 239306 106264 239312 106276
rect 239180 106236 239312 106264
rect 239180 106224 239186 106236
rect 239306 106224 239312 106236
rect 239364 106224 239370 106276
rect 251450 106264 251456 106276
rect 251411 106236 251456 106264
rect 251450 106224 251456 106236
rect 251508 106224 251514 106276
rect 259730 106224 259736 106276
rect 259788 106264 259794 106276
rect 259822 106264 259828 106276
rect 259788 106236 259828 106264
rect 259788 106224 259794 106236
rect 259822 106224 259828 106236
rect 259880 106224 259886 106276
rect 266722 106224 266728 106276
rect 266780 106264 266786 106276
rect 266814 106264 266820 106276
rect 266780 106236 266820 106264
rect 266780 106224 266786 106236
rect 266814 106224 266820 106236
rect 266872 106224 266878 106276
rect 267826 106224 267832 106276
rect 267884 106264 267890 106276
rect 267918 106264 267924 106276
rect 267884 106236 267924 106264
rect 267884 106224 267890 106236
rect 267918 106224 267924 106236
rect 267976 106224 267982 106276
rect 270678 106264 270684 106276
rect 270639 106236 270684 106264
rect 270678 106224 270684 106236
rect 270736 106224 270742 106276
rect 272150 106224 272156 106276
rect 272208 106264 272214 106276
rect 272426 106264 272432 106276
rect 272208 106236 272432 106264
rect 272208 106224 272214 106236
rect 272426 106224 272432 106236
rect 272484 106224 272490 106276
rect 358648 106196 358676 106292
rect 360378 106224 360384 106276
rect 360436 106264 360442 106276
rect 360562 106264 360568 106276
rect 360436 106236 360568 106264
rect 360436 106224 360442 106236
rect 360562 106224 360568 106236
rect 360620 106224 360626 106276
rect 372706 106224 372712 106276
rect 372764 106264 372770 106276
rect 372798 106264 372804 106276
rect 372764 106236 372804 106264
rect 372764 106224 372770 106236
rect 372798 106224 372804 106236
rect 372856 106224 372862 106276
rect 386506 106264 386512 106276
rect 386467 106236 386512 106264
rect 386506 106224 386512 106236
rect 386564 106224 386570 106276
rect 358722 106196 358728 106208
rect 358648 106168 358728 106196
rect 358722 106156 358728 106168
rect 358780 106156 358786 106208
rect 289906 104864 289912 104916
rect 289964 104904 289970 104916
rect 289998 104904 290004 104916
rect 289964 104876 290004 104904
rect 289964 104864 289970 104876
rect 289998 104864 290004 104876
rect 290056 104864 290062 104916
rect 317782 104864 317788 104916
rect 317840 104904 317846 104916
rect 317966 104904 317972 104916
rect 317840 104876 317972 104904
rect 317840 104864 317846 104876
rect 317966 104864 317972 104876
rect 318024 104864 318030 104916
rect 325970 104904 325976 104916
rect 325931 104876 325976 104904
rect 325970 104864 325976 104876
rect 326028 104864 326034 104916
rect 327166 104904 327172 104916
rect 327127 104876 327172 104904
rect 327166 104864 327172 104876
rect 327224 104864 327230 104916
rect 339770 104864 339776 104916
rect 339828 104904 339834 104916
rect 339862 104904 339868 104916
rect 339828 104876 339868 104904
rect 339828 104864 339834 104876
rect 339862 104864 339868 104876
rect 339920 104864 339926 104916
rect 357526 104864 357532 104916
rect 357584 104904 357590 104916
rect 357710 104904 357716 104916
rect 357584 104876 357716 104904
rect 357584 104864 357590 104876
rect 357710 104864 357716 104876
rect 357768 104864 357774 104916
rect 232314 104836 232320 104848
rect 232275 104808 232320 104836
rect 232314 104796 232320 104808
rect 232372 104796 232378 104848
rect 324590 104796 324596 104848
rect 324648 104836 324654 104848
rect 324682 104836 324688 104848
rect 324648 104808 324688 104836
rect 324648 104796 324654 104808
rect 324682 104796 324688 104808
rect 324740 104796 324746 104848
rect 341150 104836 341156 104848
rect 341111 104808 341156 104836
rect 341150 104796 341156 104808
rect 341208 104796 341214 104848
rect 421190 104836 421196 104848
rect 421151 104808 421196 104836
rect 421190 104796 421196 104808
rect 421248 104796 421254 104848
rect 339770 104768 339776 104780
rect 339731 104740 339776 104768
rect 339770 104728 339776 104740
rect 339828 104728 339834 104780
rect 358722 104728 358728 104780
rect 358780 104768 358786 104780
rect 358998 104768 359004 104780
rect 358780 104740 359004 104768
rect 358780 104728 358786 104740
rect 358998 104728 359004 104740
rect 359056 104728 359062 104780
rect 291565 103615 291623 103621
rect 291565 103581 291577 103615
rect 291611 103612 291623 103615
rect 291654 103612 291660 103624
rect 291611 103584 291660 103612
rect 291611 103581 291623 103584
rect 291565 103575 291623 103581
rect 291654 103572 291660 103584
rect 291712 103572 291718 103624
rect 265250 103544 265256 103556
rect 265211 103516 265256 103544
rect 265250 103504 265256 103516
rect 265308 103504 265314 103556
rect 284662 103544 284668 103556
rect 284623 103516 284668 103544
rect 284662 103504 284668 103516
rect 284720 103504 284726 103556
rect 288802 103504 288808 103556
rect 288860 103544 288866 103556
rect 288894 103544 288900 103556
rect 288860 103516 288900 103544
rect 288860 103504 288866 103516
rect 288894 103504 288900 103516
rect 288952 103504 288958 103556
rect 296806 103544 296812 103556
rect 296767 103516 296812 103544
rect 296806 103504 296812 103516
rect 296864 103504 296870 103556
rect 262582 103436 262588 103488
rect 262640 103476 262646 103488
rect 262766 103476 262772 103488
rect 262640 103448 262772 103476
rect 262640 103436 262646 103448
rect 262766 103436 262772 103448
rect 262824 103436 262830 103488
rect 266814 103476 266820 103488
rect 266775 103448 266820 103476
rect 266814 103436 266820 103448
rect 266872 103436 266878 103488
rect 267918 103476 267924 103488
rect 267879 103448 267924 103476
rect 267918 103436 267924 103448
rect 267976 103436 267982 103488
rect 289998 103436 290004 103488
rect 290056 103436 290062 103488
rect 295610 103476 295616 103488
rect 295571 103448 295616 103476
rect 295610 103436 295616 103448
rect 295668 103436 295674 103488
rect 301133 103479 301191 103485
rect 301133 103445 301145 103479
rect 301179 103476 301191 103479
rect 301222 103476 301228 103488
rect 301179 103448 301228 103476
rect 301179 103445 301191 103448
rect 301133 103439 301191 103445
rect 301222 103436 301228 103448
rect 301280 103436 301286 103488
rect 306834 103476 306840 103488
rect 306795 103448 306840 103476
rect 306834 103436 306840 103448
rect 306892 103436 306898 103488
rect 324593 103479 324651 103485
rect 324593 103445 324605 103479
rect 324639 103476 324651 103479
rect 324682 103476 324688 103488
rect 324639 103448 324688 103476
rect 324639 103445 324651 103448
rect 324593 103439 324651 103445
rect 324682 103436 324688 103448
rect 324740 103436 324746 103488
rect 330110 103436 330116 103488
rect 330168 103476 330174 103488
rect 330202 103476 330208 103488
rect 330168 103448 330208 103476
rect 330168 103436 330174 103448
rect 330202 103436 330208 103448
rect 330260 103436 330266 103488
rect 290016 103408 290044 103436
rect 290090 103408 290096 103420
rect 290016 103380 290096 103408
rect 290090 103368 290096 103380
rect 290148 103368 290154 103420
rect 296898 103368 296904 103420
rect 296956 103408 296962 103420
rect 297082 103408 297088 103420
rect 296956 103380 297088 103408
rect 296956 103368 296962 103380
rect 297082 103368 297088 103380
rect 297140 103368 297146 103420
rect 294322 102184 294328 102196
rect 294283 102156 294328 102184
rect 294322 102144 294328 102156
rect 294380 102144 294386 102196
rect 262766 102116 262772 102128
rect 262727 102088 262772 102116
rect 262766 102076 262772 102088
rect 262824 102076 262830 102128
rect 291654 102116 291660 102128
rect 291615 102088 291660 102116
rect 291654 102076 291660 102088
rect 291712 102076 291718 102128
rect 330113 102119 330171 102125
rect 330113 102085 330125 102119
rect 330159 102116 330171 102119
rect 330202 102116 330208 102128
rect 330159 102088 330208 102116
rect 330159 102085 330171 102088
rect 330113 102079 330171 102085
rect 330202 102076 330208 102088
rect 330260 102076 330266 102128
rect 270678 101368 270684 101380
rect 270639 101340 270684 101368
rect 270678 101328 270684 101340
rect 270736 101328 270742 101380
rect 337102 99424 337108 99476
rect 337160 99424 337166 99476
rect 460106 99424 460112 99476
rect 460164 99424 460170 99476
rect 244366 99356 244372 99408
rect 244424 99396 244430 99408
rect 244424 99368 244504 99396
rect 244424 99356 244430 99368
rect 244476 99340 244504 99368
rect 337120 99340 337148 99424
rect 377030 99356 377036 99408
rect 377088 99396 377094 99408
rect 377088 99368 377168 99396
rect 377088 99356 377094 99368
rect 377140 99340 377168 99368
rect 460124 99340 460152 99424
rect 244458 99288 244464 99340
rect 244516 99288 244522 99340
rect 337102 99288 337108 99340
rect 337160 99288 337166 99340
rect 375558 99288 375564 99340
rect 375616 99328 375622 99340
rect 375742 99328 375748 99340
rect 375616 99300 375748 99328
rect 375616 99288 375622 99300
rect 375742 99288 375748 99300
rect 375800 99288 375806 99340
rect 377122 99288 377128 99340
rect 377180 99288 377186 99340
rect 386506 99328 386512 99340
rect 386467 99300 386512 99328
rect 386506 99288 386512 99300
rect 386564 99288 386570 99340
rect 460106 99288 460112 99340
rect 460164 99288 460170 99340
rect 463694 98948 463700 99000
rect 463752 98988 463758 99000
rect 463878 98988 463884 99000
rect 463752 98960 463884 98988
rect 463752 98948 463758 98960
rect 463878 98948 463884 98960
rect 463936 98948 463942 99000
rect 310882 96812 310888 96824
rect 310808 96784 310888 96812
rect 310808 96688 310836 96784
rect 310882 96772 310888 96784
rect 310940 96772 310946 96824
rect 247126 96636 247132 96688
rect 247184 96676 247190 96688
rect 247218 96676 247224 96688
rect 247184 96648 247224 96676
rect 247184 96636 247190 96648
rect 247218 96636 247224 96648
rect 247276 96636 247282 96688
rect 250070 96636 250076 96688
rect 250128 96676 250134 96688
rect 250162 96676 250168 96688
rect 250128 96648 250168 96676
rect 250128 96636 250134 96648
rect 250162 96636 250168 96648
rect 250220 96636 250226 96688
rect 251450 96676 251456 96688
rect 251411 96648 251456 96676
rect 251450 96636 251456 96648
rect 251508 96636 251514 96688
rect 310790 96636 310796 96688
rect 310848 96636 310854 96688
rect 270678 96568 270684 96620
rect 270736 96608 270742 96620
rect 270862 96608 270868 96620
rect 270736 96580 270868 96608
rect 270736 96568 270742 96580
rect 270862 96568 270868 96580
rect 270920 96568 270926 96620
rect 360286 96608 360292 96620
rect 360247 96580 360292 96608
rect 360286 96568 360292 96580
rect 360344 96568 360350 96620
rect 367002 96608 367008 96620
rect 366963 96580 367008 96608
rect 367002 96568 367008 96580
rect 367060 96568 367066 96620
rect 375374 96568 375380 96620
rect 375432 96608 375438 96620
rect 375558 96608 375564 96620
rect 375432 96580 375564 96608
rect 375432 96568 375438 96580
rect 375558 96568 375564 96580
rect 375616 96568 375622 96620
rect 470594 96608 470600 96620
rect 470555 96580 470600 96608
rect 470594 96568 470600 96580
rect 470652 96568 470658 96620
rect 266814 96472 266820 96484
rect 266775 96444 266820 96472
rect 266814 96432 266820 96444
rect 266872 96432 266878 96484
rect 273530 95276 273536 95328
rect 273588 95316 273594 95328
rect 273622 95316 273628 95328
rect 273588 95288 273628 95316
rect 273588 95276 273594 95288
rect 273622 95276 273628 95288
rect 273680 95276 273686 95328
rect 232314 95248 232320 95260
rect 232275 95220 232320 95248
rect 232314 95208 232320 95220
rect 232372 95208 232378 95260
rect 339773 95251 339831 95257
rect 339773 95217 339785 95251
rect 339819 95248 339831 95251
rect 339954 95248 339960 95260
rect 339819 95220 339960 95248
rect 339819 95217 339831 95220
rect 339773 95211 339831 95217
rect 339954 95208 339960 95220
rect 340012 95208 340018 95260
rect 341150 95248 341156 95260
rect 341111 95220 341156 95248
rect 341150 95208 341156 95220
rect 341208 95208 341214 95260
rect 247126 95180 247132 95192
rect 247087 95152 247132 95180
rect 247126 95140 247132 95152
rect 247184 95140 247190 95192
rect 284662 95140 284668 95192
rect 284720 95140 284726 95192
rect 310790 95180 310796 95192
rect 310751 95152 310796 95180
rect 310790 95140 310796 95152
rect 310848 95140 310854 95192
rect 284680 95112 284708 95140
rect 284754 95112 284760 95124
rect 284680 95084 284760 95112
rect 284754 95072 284760 95084
rect 284812 95072 284818 95124
rect 317966 93916 317972 93968
rect 318024 93916 318030 93968
rect 265158 93848 265164 93900
rect 265216 93888 265222 93900
rect 265250 93888 265256 93900
rect 265216 93860 265256 93888
rect 265216 93848 265222 93860
rect 265250 93848 265256 93860
rect 265308 93848 265314 93900
rect 267734 93848 267740 93900
rect 267792 93888 267798 93900
rect 267921 93891 267979 93897
rect 267921 93888 267933 93891
rect 267792 93860 267933 93888
rect 267792 93848 267798 93860
rect 267921 93857 267933 93860
rect 267967 93857 267979 93891
rect 295610 93888 295616 93900
rect 295571 93860 295616 93888
rect 267921 93851 267979 93857
rect 295610 93848 295616 93860
rect 295668 93848 295674 93900
rect 301130 93888 301136 93900
rect 301091 93860 301136 93888
rect 301130 93848 301136 93860
rect 301188 93848 301194 93900
rect 306834 93888 306840 93900
rect 306795 93860 306840 93888
rect 306834 93848 306840 93860
rect 306892 93848 306898 93900
rect 317690 93848 317696 93900
rect 317748 93888 317754 93900
rect 317984 93888 318012 93916
rect 324590 93888 324596 93900
rect 317748 93860 318012 93888
rect 324551 93860 324596 93888
rect 317748 93848 317754 93860
rect 324590 93848 324596 93860
rect 324648 93848 324654 93900
rect 262766 92528 262772 92540
rect 262727 92500 262772 92528
rect 262766 92488 262772 92500
rect 262824 92488 262830 92540
rect 291654 92528 291660 92540
rect 291615 92500 291660 92528
rect 291654 92488 291660 92500
rect 291712 92488 291718 92540
rect 341061 90423 341119 90429
rect 341061 90389 341073 90423
rect 341107 90420 341119 90423
rect 341150 90420 341156 90432
rect 341107 90392 341156 90420
rect 341107 90389 341119 90392
rect 341061 90383 341119 90389
rect 341150 90380 341156 90392
rect 341208 90380 341214 90432
rect 386414 89700 386420 89752
rect 386472 89740 386478 89752
rect 386598 89740 386604 89752
rect 386472 89712 386604 89740
rect 386472 89700 386478 89712
rect 386598 89700 386604 89712
rect 386656 89700 386662 89752
rect 360286 89672 360292 89684
rect 360247 89644 360292 89672
rect 360286 89632 360292 89644
rect 360344 89632 360350 89684
rect 262677 88995 262735 89001
rect 262677 88961 262689 88995
rect 262723 88992 262735 88995
rect 262766 88992 262772 89004
rect 262723 88964 262772 88992
rect 262723 88961 262735 88964
rect 262677 88955 262735 88961
rect 262766 88952 262772 88964
rect 262824 88952 262830 89004
rect 265158 88992 265164 89004
rect 265119 88964 265164 88992
rect 265158 88952 265164 88964
rect 265216 88952 265222 89004
rect 317690 88380 317696 88392
rect 317651 88352 317696 88380
rect 317690 88340 317696 88352
rect 317748 88340 317754 88392
rect 454034 87252 454040 87304
rect 454092 87292 454098 87304
rect 456978 87292 456984 87304
rect 454092 87264 456984 87292
rect 454092 87252 454098 87264
rect 456978 87252 456984 87264
rect 457036 87252 457042 87304
rect 437198 87116 437204 87168
rect 437256 87156 437262 87168
rect 437474 87156 437480 87168
rect 437256 87128 437480 87156
rect 437256 87116 437262 87128
rect 437474 87116 437480 87128
rect 437532 87116 437538 87168
rect 494606 87116 494612 87168
rect 494664 87156 494670 87168
rect 502242 87156 502248 87168
rect 494664 87128 502248 87156
rect 494664 87116 494670 87128
rect 502242 87116 502248 87128
rect 502300 87116 502306 87168
rect 251174 87048 251180 87100
rect 251232 87088 251238 87100
rect 260650 87088 260656 87100
rect 251232 87060 260656 87088
rect 251232 87048 251238 87060
rect 260650 87048 260656 87060
rect 260708 87048 260714 87100
rect 347774 86980 347780 87032
rect 347832 87020 347838 87032
rect 357342 87020 357348 87032
rect 347832 86992 357348 87020
rect 347832 86980 347838 86992
rect 357342 86980 357348 86992
rect 357400 86980 357406 87032
rect 367002 87020 367008 87032
rect 366963 86992 367008 87020
rect 367002 86980 367008 86992
rect 367060 86980 367066 87032
rect 421190 87020 421196 87032
rect 421151 86992 421196 87020
rect 421190 86980 421196 86992
rect 421248 86980 421254 87032
rect 470594 87020 470600 87032
rect 470555 86992 470600 87020
rect 470594 86980 470600 86992
rect 470652 86980 470658 87032
rect 236273 86955 236331 86961
rect 236273 86921 236285 86955
rect 236319 86952 236331 86955
rect 236454 86952 236460 86964
rect 236319 86924 236460 86952
rect 236319 86921 236331 86924
rect 236273 86915 236331 86921
rect 236454 86912 236460 86924
rect 236512 86912 236518 86964
rect 251450 86952 251456 86964
rect 251411 86924 251456 86952
rect 251450 86912 251456 86924
rect 251508 86912 251514 86964
rect 323302 86912 323308 86964
rect 323360 86952 323366 86964
rect 323394 86952 323400 86964
rect 323360 86924 323400 86952
rect 323360 86912 323366 86924
rect 323394 86912 323400 86924
rect 323452 86912 323458 86964
rect 324590 86912 324596 86964
rect 324648 86912 324654 86964
rect 325878 86912 325884 86964
rect 325936 86912 325942 86964
rect 327166 86912 327172 86964
rect 327224 86952 327230 86964
rect 327258 86952 327264 86964
rect 327224 86924 327264 86952
rect 327224 86912 327230 86924
rect 327258 86912 327264 86924
rect 327316 86912 327322 86964
rect 336918 86952 336924 86964
rect 336879 86924 336924 86952
rect 336918 86912 336924 86924
rect 336976 86912 336982 86964
rect 337194 86952 337200 86964
rect 337155 86924 337200 86952
rect 337194 86912 337200 86924
rect 337252 86912 337258 86964
rect 324608 86884 324636 86912
rect 324682 86884 324688 86896
rect 324608 86856 324688 86884
rect 324682 86844 324688 86856
rect 324740 86844 324746 86896
rect 325896 86884 325924 86912
rect 325970 86884 325976 86896
rect 325896 86856 325976 86884
rect 325970 86844 325976 86856
rect 326028 86844 326034 86896
rect 360194 86844 360200 86896
rect 360252 86884 360258 86896
rect 360378 86884 360384 86896
rect 360252 86856 360384 86884
rect 360252 86844 360258 86856
rect 360378 86844 360384 86856
rect 360436 86844 360442 86896
rect 375558 86844 375564 86896
rect 375616 86884 375622 86896
rect 375650 86884 375656 86896
rect 375616 86856 375656 86884
rect 375616 86844 375622 86856
rect 375650 86844 375656 86856
rect 375708 86844 375714 86896
rect 286226 85660 286232 85672
rect 285968 85632 286232 85660
rect 285968 85604 285996 85632
rect 286226 85620 286232 85632
rect 286284 85620 286290 85672
rect 247129 85595 247187 85601
rect 247129 85561 247141 85595
rect 247175 85592 247187 85595
rect 247218 85592 247224 85604
rect 247175 85564 247224 85592
rect 247175 85561 247187 85564
rect 247129 85555 247187 85561
rect 247218 85552 247224 85564
rect 247276 85552 247282 85604
rect 285950 85552 285956 85604
rect 286008 85552 286014 85604
rect 291565 85595 291623 85601
rect 291565 85561 291577 85595
rect 291611 85592 291623 85595
rect 291654 85592 291660 85604
rect 291611 85564 291660 85592
rect 291611 85561 291623 85564
rect 291565 85555 291623 85561
rect 291654 85552 291660 85564
rect 291712 85552 291718 85604
rect 294230 85552 294236 85604
rect 294288 85592 294294 85604
rect 294322 85592 294328 85604
rect 294288 85564 294328 85592
rect 294288 85552 294294 85564
rect 294322 85552 294328 85564
rect 294380 85552 294386 85604
rect 310790 85592 310796 85604
rect 310751 85564 310796 85592
rect 310790 85552 310796 85564
rect 310848 85552 310854 85604
rect 232314 85524 232320 85536
rect 232275 85496 232320 85524
rect 232314 85484 232320 85496
rect 232372 85484 232378 85536
rect 267734 85484 267740 85536
rect 267792 85524 267798 85536
rect 267826 85524 267832 85536
rect 267792 85496 267832 85524
rect 267792 85484 267798 85496
rect 267826 85484 267832 85496
rect 267884 85484 267890 85536
rect 273530 85484 273536 85536
rect 273588 85524 273594 85536
rect 273622 85524 273628 85536
rect 273588 85496 273628 85524
rect 273588 85484 273594 85496
rect 273622 85484 273628 85496
rect 273680 85484 273686 85536
rect 299842 85524 299848 85536
rect 299803 85496 299848 85524
rect 299842 85484 299848 85496
rect 299900 85484 299906 85536
rect 301038 85484 301044 85536
rect 301096 85524 301102 85536
rect 301222 85524 301228 85536
rect 301096 85496 301228 85524
rect 301096 85484 301102 85496
rect 301222 85484 301228 85496
rect 301280 85484 301286 85536
rect 306650 85484 306656 85536
rect 306708 85524 306714 85536
rect 306834 85524 306840 85536
rect 306708 85496 306840 85524
rect 306708 85484 306714 85496
rect 306834 85484 306840 85496
rect 306892 85484 306898 85536
rect 324682 85524 324688 85536
rect 324643 85496 324688 85524
rect 324682 85484 324688 85496
rect 324740 85484 324746 85536
rect 358722 85524 358728 85536
rect 358683 85496 358728 85524
rect 358722 85484 358728 85496
rect 358780 85484 358786 85536
rect 421190 85524 421196 85536
rect 421151 85496 421196 85524
rect 421190 85484 421196 85496
rect 421248 85484 421254 85536
rect 265161 84303 265219 84309
rect 265161 84269 265173 84303
rect 265207 84300 265219 84303
rect 265207 84272 265388 84300
rect 265207 84269 265219 84272
rect 265161 84263 265219 84269
rect 265360 84173 265388 84272
rect 296990 84260 296996 84312
rect 297048 84300 297054 84312
rect 297048 84272 297128 84300
rect 297048 84260 297054 84272
rect 297100 84244 297128 84272
rect 291562 84232 291568 84244
rect 291523 84204 291568 84232
rect 291562 84192 291568 84204
rect 291620 84192 291626 84244
rect 297082 84192 297088 84244
rect 297140 84192 297146 84244
rect 265345 84167 265403 84173
rect 265345 84133 265357 84167
rect 265391 84133 265403 84167
rect 265345 84127 265403 84133
rect 272245 84167 272303 84173
rect 272245 84133 272257 84167
rect 272291 84164 272303 84167
rect 272334 84164 272340 84176
rect 272291 84136 272340 84164
rect 272291 84133 272303 84136
rect 272245 84127 272303 84133
rect 272334 84124 272340 84136
rect 272392 84124 272398 84176
rect 284665 84167 284723 84173
rect 284665 84133 284677 84167
rect 284711 84164 284723 84167
rect 284754 84164 284760 84176
rect 284711 84136 284760 84164
rect 284711 84133 284723 84136
rect 284665 84127 284723 84133
rect 284754 84124 284760 84136
rect 284812 84124 284818 84176
rect 285950 84164 285956 84176
rect 285911 84136 285956 84164
rect 285950 84124 285956 84136
rect 286008 84124 286014 84176
rect 288710 82804 288716 82816
rect 288671 82776 288716 82804
rect 288710 82764 288716 82776
rect 288768 82764 288774 82816
rect 270770 80764 270776 80776
rect 270731 80736 270776 80764
rect 270770 80724 270776 80736
rect 270828 80724 270834 80776
rect 357710 80152 357716 80164
rect 357636 80124 357716 80152
rect 357636 80096 357664 80124
rect 357710 80112 357716 80124
rect 357768 80112 357774 80164
rect 359182 80152 359188 80164
rect 359108 80124 359188 80152
rect 359108 80096 359136 80124
rect 359182 80112 359188 80124
rect 359240 80112 359246 80164
rect 372798 80152 372804 80164
rect 372724 80124 372804 80152
rect 372724 80096 372752 80124
rect 372798 80112 372804 80124
rect 372856 80112 372862 80164
rect 303890 80044 303896 80096
rect 303948 80044 303954 80096
rect 357618 80044 357624 80096
rect 357676 80044 357682 80096
rect 359090 80044 359096 80096
rect 359148 80044 359154 80096
rect 372706 80044 372712 80096
rect 372764 80044 372770 80096
rect 303908 79960 303936 80044
rect 303890 79908 303896 79960
rect 303948 79908 303954 79960
rect 2774 79772 2780 79824
rect 2832 79812 2838 79824
rect 4890 79812 4896 79824
rect 2832 79784 4896 79812
rect 2832 79772 2838 79784
rect 4890 79772 4896 79784
rect 4948 79772 4954 79824
rect 236270 77432 236276 77444
rect 236231 77404 236276 77432
rect 236270 77392 236276 77404
rect 236328 77392 236334 77444
rect 358814 77324 358820 77376
rect 358872 77324 358878 77376
rect 358906 77324 358912 77376
rect 358964 77324 358970 77376
rect 251450 77296 251456 77308
rect 251411 77268 251456 77296
rect 251450 77256 251456 77268
rect 251508 77256 251514 77308
rect 330113 77299 330171 77305
rect 330113 77265 330125 77299
rect 330159 77296 330171 77299
rect 330202 77296 330208 77308
rect 330159 77268 330208 77296
rect 330159 77265 330171 77268
rect 330113 77259 330171 77265
rect 330202 77256 330208 77268
rect 330260 77256 330266 77308
rect 337194 77296 337200 77308
rect 337155 77268 337200 77296
rect 337194 77256 337200 77268
rect 337252 77256 337258 77308
rect 339770 77256 339776 77308
rect 339828 77296 339834 77308
rect 339954 77296 339960 77308
rect 339828 77268 339960 77296
rect 339828 77256 339834 77268
rect 339954 77256 339960 77268
rect 340012 77256 340018 77308
rect 341058 77296 341064 77308
rect 341019 77268 341064 77296
rect 341058 77256 341064 77268
rect 341116 77256 341122 77308
rect 358832 77240 358860 77324
rect 358924 77240 358952 77324
rect 303890 77188 303896 77240
rect 303948 77228 303954 77240
rect 303982 77228 303988 77240
rect 303948 77200 303988 77228
rect 303948 77188 303954 77200
rect 303982 77188 303988 77200
rect 304040 77188 304046 77240
rect 358814 77188 358820 77240
rect 358872 77188 358878 77240
rect 358906 77188 358912 77240
rect 358964 77188 358970 77240
rect 386601 77231 386659 77237
rect 386601 77197 386613 77231
rect 386647 77228 386659 77231
rect 386690 77228 386696 77240
rect 386647 77200 386696 77228
rect 386647 77197 386659 77200
rect 386601 77191 386659 77197
rect 386690 77188 386696 77200
rect 386748 77188 386754 77240
rect 470594 77228 470600 77240
rect 470555 77200 470600 77228
rect 470594 77188 470600 77200
rect 470652 77188 470658 77240
rect 310790 76100 310796 76152
rect 310848 76100 310854 76152
rect 328914 76100 328920 76152
rect 328972 76140 328978 76152
rect 338022 76140 338028 76152
rect 328972 76112 338028 76140
rect 328972 76100 328978 76112
rect 338022 76100 338028 76112
rect 338080 76100 338086 76152
rect 369854 76100 369860 76152
rect 369912 76140 369918 76152
rect 376662 76140 376668 76152
rect 369912 76112 376668 76140
rect 369912 76100 369918 76112
rect 376662 76100 376668 76112
rect 376720 76100 376726 76152
rect 310808 76016 310836 76100
rect 396074 76032 396080 76084
rect 396132 76072 396138 76084
rect 399386 76072 399392 76084
rect 396132 76044 399392 76072
rect 396132 76032 396138 76044
rect 399386 76032 399392 76044
rect 399444 76032 399450 76084
rect 414014 76032 414020 76084
rect 414072 76072 414078 76084
rect 423398 76072 423404 76084
rect 414072 76044 423404 76072
rect 414072 76032 414078 76044
rect 423398 76032 423404 76044
rect 423456 76032 423462 76084
rect 437198 76032 437204 76084
rect 437256 76072 437262 76084
rect 437474 76072 437480 76084
rect 437256 76044 437480 76072
rect 437256 76032 437262 76044
rect 437474 76032 437480 76044
rect 437532 76032 437538 76084
rect 310790 75964 310796 76016
rect 310848 75964 310854 76016
rect 324682 76004 324688 76016
rect 324643 75976 324688 76004
rect 324682 75964 324688 75976
rect 324740 75964 324746 76016
rect 232314 75936 232320 75948
rect 232275 75908 232320 75936
rect 232314 75896 232320 75908
rect 232372 75896 232378 75948
rect 262674 75936 262680 75948
rect 262635 75908 262680 75936
rect 262674 75896 262680 75908
rect 262732 75896 262738 75948
rect 289906 75896 289912 75948
rect 289964 75936 289970 75948
rect 290090 75936 290096 75948
rect 289964 75908 290096 75936
rect 289964 75896 289970 75908
rect 290090 75896 290096 75908
rect 290148 75896 290154 75948
rect 291378 75896 291384 75948
rect 291436 75936 291442 75948
rect 291562 75936 291568 75948
rect 291436 75908 291568 75936
rect 291436 75896 291442 75908
rect 291562 75896 291568 75908
rect 291620 75896 291626 75948
rect 295518 75896 295524 75948
rect 295576 75936 295582 75948
rect 295702 75936 295708 75948
rect 295576 75908 295708 75936
rect 295576 75896 295582 75908
rect 295702 75896 295708 75908
rect 295760 75896 295766 75948
rect 299842 75936 299848 75948
rect 299803 75908 299848 75936
rect 299842 75896 299848 75908
rect 299900 75896 299906 75948
rect 302510 75896 302516 75948
rect 302568 75936 302574 75948
rect 302602 75936 302608 75948
rect 302568 75908 302608 75936
rect 302568 75896 302574 75908
rect 302602 75896 302608 75908
rect 302660 75896 302666 75948
rect 317690 75936 317696 75948
rect 317651 75908 317696 75936
rect 317690 75896 317696 75908
rect 317748 75896 317754 75948
rect 336918 75936 336924 75948
rect 336879 75908 336924 75936
rect 336918 75896 336924 75908
rect 336976 75896 336982 75948
rect 358725 75939 358783 75945
rect 358725 75905 358737 75939
rect 358771 75936 358783 75939
rect 358998 75936 359004 75948
rect 358771 75908 359004 75936
rect 358771 75905 358783 75908
rect 358725 75899 358783 75905
rect 358998 75896 359004 75908
rect 359056 75896 359062 75948
rect 421190 75936 421196 75948
rect 421151 75908 421196 75936
rect 421190 75896 421196 75908
rect 421248 75896 421254 75948
rect 310790 75868 310796 75880
rect 310751 75840 310796 75868
rect 310790 75828 310796 75840
rect 310848 75828 310854 75880
rect 324593 75871 324651 75877
rect 324593 75837 324605 75871
rect 324639 75868 324651 75871
rect 324682 75868 324688 75880
rect 324639 75840 324688 75868
rect 324639 75837 324651 75840
rect 324593 75831 324651 75837
rect 324682 75828 324688 75840
rect 324740 75828 324746 75880
rect 296806 74604 296812 74656
rect 296864 74644 296870 74656
rect 297082 74644 297088 74656
rect 296864 74616 297088 74644
rect 296864 74604 296870 74616
rect 297082 74604 297088 74616
rect 297140 74604 297146 74656
rect 265345 74579 265403 74585
rect 265345 74545 265357 74579
rect 265391 74576 265403 74579
rect 265434 74576 265440 74588
rect 265391 74548 265440 74576
rect 265391 74545 265403 74548
rect 265345 74539 265403 74545
rect 265434 74536 265440 74548
rect 265492 74536 265498 74588
rect 272242 74576 272248 74588
rect 272203 74548 272248 74576
rect 272242 74536 272248 74548
rect 272300 74536 272306 74588
rect 239122 70496 239128 70508
rect 239083 70468 239128 70496
rect 239122 70456 239128 70468
rect 239180 70456 239186 70508
rect 244458 70496 244464 70508
rect 244419 70468 244464 70496
rect 244458 70456 244464 70468
rect 244516 70456 244522 70508
rect 377122 70496 377128 70508
rect 377083 70468 377128 70496
rect 377122 70456 377128 70468
rect 377180 70456 377186 70508
rect 367002 67736 367008 67788
rect 367060 67736 367066 67788
rect 272242 67708 272248 67720
rect 272203 67680 272248 67708
rect 272242 67668 272248 67680
rect 272300 67668 272306 67720
rect 323302 67668 323308 67720
rect 323360 67668 323366 67720
rect 239122 67640 239128 67652
rect 239083 67612 239128 67640
rect 239122 67600 239128 67612
rect 239180 67600 239186 67652
rect 244458 67640 244464 67652
rect 244419 67612 244464 67640
rect 244458 67600 244464 67612
rect 244516 67600 244522 67652
rect 270770 67640 270776 67652
rect 270731 67612 270776 67640
rect 270770 67600 270776 67612
rect 270828 67600 270834 67652
rect 299750 67600 299756 67652
rect 299808 67640 299814 67652
rect 299842 67640 299848 67652
rect 299808 67612 299848 67640
rect 299808 67600 299814 67612
rect 299842 67600 299848 67612
rect 299900 67600 299906 67652
rect 323320 67640 323348 67668
rect 367020 67652 367048 67736
rect 323394 67640 323400 67652
rect 323320 67612 323400 67640
rect 323394 67600 323400 67612
rect 323452 67600 323458 67652
rect 341058 67600 341064 67652
rect 341116 67640 341122 67652
rect 341150 67640 341156 67652
rect 341116 67612 341156 67640
rect 341116 67600 341122 67612
rect 341150 67600 341156 67612
rect 341208 67600 341214 67652
rect 358722 67600 358728 67652
rect 358780 67640 358786 67652
rect 358998 67640 359004 67652
rect 358780 67612 359004 67640
rect 358780 67600 358786 67612
rect 358998 67600 359004 67612
rect 359056 67600 359062 67652
rect 367002 67600 367008 67652
rect 367060 67600 367066 67652
rect 377122 67640 377128 67652
rect 377083 67612 377128 67640
rect 377122 67600 377128 67612
rect 377180 67600 377186 67652
rect 386598 67640 386604 67652
rect 386559 67612 386604 67640
rect 386598 67600 386604 67612
rect 386656 67600 386662 67652
rect 470594 67640 470600 67652
rect 470555 67612 470600 67640
rect 470594 67600 470600 67612
rect 470652 67600 470658 67652
rect 236270 67532 236276 67584
rect 236328 67572 236334 67584
rect 236362 67572 236368 67584
rect 236328 67544 236368 67572
rect 236328 67532 236334 67544
rect 236362 67532 236368 67544
rect 236420 67532 236426 67584
rect 250070 67572 250076 67584
rect 250031 67544 250076 67572
rect 250070 67532 250076 67544
rect 250128 67532 250134 67584
rect 375650 67572 375656 67584
rect 375611 67544 375656 67572
rect 375650 67532 375656 67544
rect 375708 67532 375714 67584
rect 459922 67532 459928 67584
rect 459980 67572 459986 67584
rect 460198 67572 460204 67584
rect 459980 67544 460204 67572
rect 459980 67532 459986 67544
rect 460198 67532 460204 67544
rect 460256 67532 460262 67584
rect 272242 67096 272248 67108
rect 272203 67068 272248 67096
rect 272242 67056 272248 67068
rect 272300 67056 272306 67108
rect 310790 66348 310796 66360
rect 310751 66320 310796 66348
rect 310790 66308 310796 66320
rect 310848 66308 310854 66360
rect 324590 66348 324596 66360
rect 324551 66320 324596 66348
rect 324590 66308 324596 66320
rect 324648 66308 324654 66360
rect 267734 66240 267740 66292
rect 267792 66280 267798 66292
rect 267826 66280 267832 66292
rect 267792 66252 267832 66280
rect 267792 66240 267798 66252
rect 267826 66240 267832 66252
rect 267884 66240 267890 66292
rect 284662 66280 284668 66292
rect 284623 66252 284668 66280
rect 284662 66240 284668 66252
rect 284720 66240 284726 66292
rect 285950 66280 285956 66292
rect 285911 66252 285956 66280
rect 285950 66240 285956 66252
rect 286008 66240 286014 66292
rect 296806 66240 296812 66292
rect 296864 66240 296870 66292
rect 327258 66240 327264 66292
rect 327316 66240 327322 66292
rect 232314 66212 232320 66224
rect 232275 66184 232320 66212
rect 232314 66172 232320 66184
rect 232372 66172 232378 66224
rect 236273 66215 236331 66221
rect 236273 66181 236285 66215
rect 236319 66212 236331 66215
rect 236362 66212 236368 66224
rect 236319 66184 236368 66212
rect 236319 66181 236331 66184
rect 236273 66175 236331 66181
rect 236362 66172 236368 66184
rect 236420 66172 236426 66224
rect 270770 66212 270776 66224
rect 270731 66184 270776 66212
rect 270770 66172 270776 66184
rect 270828 66172 270834 66224
rect 273438 66212 273444 66224
rect 273399 66184 273444 66212
rect 273438 66172 273444 66184
rect 273496 66172 273502 66224
rect 296824 66144 296852 66240
rect 310790 66212 310796 66224
rect 310751 66184 310796 66212
rect 310790 66172 310796 66184
rect 310848 66172 310854 66224
rect 323305 66215 323363 66221
rect 323305 66181 323317 66215
rect 323351 66212 323363 66215
rect 323394 66212 323400 66224
rect 323351 66184 323400 66212
rect 323351 66181 323363 66184
rect 323305 66175 323363 66181
rect 323394 66172 323400 66184
rect 323452 66172 323458 66224
rect 324590 66212 324596 66224
rect 324551 66184 324596 66212
rect 324590 66172 324596 66184
rect 324648 66172 324654 66224
rect 296898 66144 296904 66156
rect 296824 66116 296904 66144
rect 296898 66104 296904 66116
rect 296956 66104 296962 66156
rect 327276 66144 327304 66240
rect 330110 66212 330116 66224
rect 330071 66184 330116 66212
rect 330110 66172 330116 66184
rect 330168 66172 330174 66224
rect 336918 66212 336924 66224
rect 336879 66184 336924 66212
rect 336918 66172 336924 66184
rect 336976 66172 336982 66224
rect 358633 66215 358691 66221
rect 358633 66181 358645 66215
rect 358679 66212 358691 66215
rect 358722 66212 358728 66224
rect 358679 66184 358728 66212
rect 358679 66181 358691 66184
rect 358633 66175 358691 66181
rect 358722 66172 358728 66184
rect 358780 66172 358786 66224
rect 367002 66212 367008 66224
rect 366963 66184 367008 66212
rect 367002 66172 367008 66184
rect 367060 66172 367066 66224
rect 421190 66212 421196 66224
rect 421151 66184 421196 66212
rect 421190 66172 421196 66184
rect 421248 66172 421254 66224
rect 327350 66144 327356 66156
rect 327276 66116 327356 66144
rect 327350 66104 327356 66116
rect 327408 66104 327414 66156
rect 306650 65764 306656 65816
rect 306708 65804 306714 65816
rect 306834 65804 306840 65816
rect 306708 65776 306840 65804
rect 306708 65764 306714 65776
rect 306834 65764 306840 65776
rect 306892 65764 306898 65816
rect 288713 64923 288771 64929
rect 288713 64889 288725 64923
rect 288759 64920 288771 64923
rect 288894 64920 288900 64932
rect 288759 64892 288900 64920
rect 288759 64889 288771 64892
rect 288713 64883 288771 64889
rect 288894 64880 288900 64892
rect 288952 64880 288958 64932
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 24118 64852 24124 64864
rect 3384 64824 24124 64852
rect 3384 64812 3390 64824
rect 24118 64812 24124 64824
rect 24176 64812 24182 64864
rect 294230 64852 294236 64864
rect 294191 64824 294236 64852
rect 294230 64812 294236 64824
rect 294288 64812 294294 64864
rect 378502 63860 378508 63912
rect 378560 63900 378566 63912
rect 386322 63900 386328 63912
rect 378560 63872 386328 63900
rect 378560 63860 378566 63872
rect 386322 63860 386328 63872
rect 386380 63860 386386 63912
rect 367094 63724 367100 63776
rect 367152 63764 367158 63776
rect 376662 63764 376668 63776
rect 367152 63736 376668 63764
rect 367152 63724 367158 63736
rect 376662 63724 376668 63736
rect 376720 63724 376726 63776
rect 417878 63656 417884 63708
rect 417936 63696 417942 63708
rect 418154 63696 418160 63708
rect 417936 63668 418160 63696
rect 417936 63656 417942 63668
rect 418154 63656 418160 63668
rect 418212 63656 418218 63708
rect 437198 63656 437204 63708
rect 437256 63696 437262 63708
rect 437474 63696 437480 63708
rect 437256 63668 437480 63696
rect 437256 63656 437262 63668
rect 437474 63656 437480 63668
rect 437532 63656 437538 63708
rect 456518 63656 456524 63708
rect 456576 63696 456582 63708
rect 456886 63696 456892 63708
rect 456576 63668 456892 63696
rect 456576 63656 456582 63668
rect 456886 63656 456892 63668
rect 456944 63656 456950 63708
rect 262582 62772 262588 62824
rect 262640 62812 262646 62824
rect 262766 62812 262772 62824
rect 262640 62784 262772 62812
rect 262640 62772 262646 62784
rect 262766 62772 262772 62784
rect 262824 62772 262830 62824
rect 259730 62636 259736 62688
rect 259788 62636 259794 62688
rect 265161 62679 265219 62685
rect 265161 62645 265173 62679
rect 265207 62676 265219 62679
rect 265342 62676 265348 62688
rect 265207 62648 265348 62676
rect 265207 62645 265219 62648
rect 265161 62639 265219 62645
rect 265342 62636 265348 62648
rect 265400 62636 265406 62688
rect 259748 62608 259776 62636
rect 259914 62608 259920 62620
rect 259748 62580 259920 62608
rect 259914 62568 259920 62580
rect 259972 62568 259978 62620
rect 375650 61996 375656 62008
rect 375611 61968 375656 61996
rect 375650 61956 375656 61968
rect 375708 61956 375714 62008
rect 324593 61387 324651 61393
rect 324593 61353 324605 61387
rect 324639 61384 324651 61387
rect 324682 61384 324688 61396
rect 324639 61356 324688 61384
rect 324639 61353 324651 61356
rect 324593 61347 324651 61353
rect 324682 61344 324688 61356
rect 324740 61344 324746 61396
rect 339678 60664 339684 60716
rect 339736 60704 339742 60716
rect 339862 60704 339868 60716
rect 339736 60676 339868 60704
rect 339736 60664 339742 60676
rect 339862 60664 339868 60676
rect 339920 60664 339926 60716
rect 341150 60664 341156 60716
rect 341208 60704 341214 60716
rect 341334 60704 341340 60716
rect 341208 60676 341340 60704
rect 341208 60664 341214 60676
rect 341334 60664 341340 60676
rect 341392 60664 341398 60716
rect 360286 60664 360292 60716
rect 360344 60704 360350 60716
rect 360470 60704 360476 60716
rect 360344 60676 360476 60704
rect 360344 60664 360350 60676
rect 360470 60664 360476 60676
rect 360528 60664 360534 60716
rect 310793 60027 310851 60033
rect 310793 59993 310805 60027
rect 310839 60024 310851 60027
rect 310882 60024 310888 60036
rect 310839 59996 310888 60024
rect 310839 59993 310851 59996
rect 310793 59987 310851 59993
rect 310882 59984 310888 59996
rect 310940 59984 310946 60036
rect 239033 58055 239091 58061
rect 239033 58021 239045 58055
rect 239079 58052 239091 58055
rect 239122 58052 239128 58064
rect 239079 58024 239128 58052
rect 239079 58021 239091 58024
rect 239033 58015 239091 58021
rect 239122 58012 239128 58024
rect 239180 58012 239186 58064
rect 291470 58052 291476 58064
rect 291396 58024 291476 58052
rect 244458 57944 244464 57996
rect 244516 57944 244522 57996
rect 250073 57987 250131 57993
rect 250073 57953 250085 57987
rect 250119 57984 250131 57987
rect 250162 57984 250168 57996
rect 250119 57956 250168 57984
rect 250119 57953 250131 57956
rect 250073 57947 250131 57953
rect 250162 57944 250168 57956
rect 250220 57944 250226 57996
rect 266722 57944 266728 57996
rect 266780 57984 266786 57996
rect 266814 57984 266820 57996
rect 266780 57956 266820 57984
rect 266780 57944 266786 57956
rect 266814 57944 266820 57956
rect 266872 57944 266878 57996
rect 267734 57944 267740 57996
rect 267792 57984 267798 57996
rect 267826 57984 267832 57996
rect 267792 57956 267832 57984
rect 267792 57944 267798 57956
rect 267826 57944 267832 57956
rect 267884 57944 267890 57996
rect 284662 57944 284668 57996
rect 284720 57984 284726 57996
rect 284754 57984 284760 57996
rect 284720 57956 284760 57984
rect 284720 57944 284726 57956
rect 284754 57944 284760 57956
rect 284812 57944 284818 57996
rect 285950 57944 285956 57996
rect 286008 57984 286014 57996
rect 286042 57984 286048 57996
rect 286008 57956 286048 57984
rect 286008 57944 286014 57956
rect 286042 57944 286048 57956
rect 286100 57944 286106 57996
rect 244476 57848 244504 57944
rect 291396 57928 291424 58024
rect 291470 58012 291476 58024
rect 291528 58012 291534 58064
rect 303890 57944 303896 57996
rect 303948 57984 303954 57996
rect 303982 57984 303988 57996
rect 303948 57956 303988 57984
rect 303948 57944 303954 57956
rect 303982 57944 303988 57956
rect 304040 57944 304046 57996
rect 265158 57916 265164 57928
rect 265119 57888 265164 57916
rect 265158 57876 265164 57888
rect 265216 57876 265222 57928
rect 291378 57876 291384 57928
rect 291436 57876 291442 57928
rect 339773 57919 339831 57925
rect 339773 57885 339785 57919
rect 339819 57916 339831 57919
rect 339862 57916 339868 57928
rect 339819 57888 339868 57916
rect 339819 57885 339831 57888
rect 339773 57879 339831 57885
rect 339862 57876 339868 57888
rect 339920 57876 339926 57928
rect 460017 57919 460075 57925
rect 460017 57885 460029 57919
rect 460063 57916 460075 57919
rect 460106 57916 460112 57928
rect 460063 57888 460112 57916
rect 460063 57885 460075 57888
rect 460017 57879 460075 57885
rect 460106 57876 460112 57888
rect 460164 57876 460170 57928
rect 470594 57916 470600 57928
rect 470555 57888 470600 57916
rect 470594 57876 470600 57888
rect 470652 57876 470658 57928
rect 244550 57848 244556 57860
rect 244476 57820 244556 57848
rect 244550 57808 244556 57820
rect 244608 57808 244614 57860
rect 301038 56652 301044 56704
rect 301096 56692 301102 56704
rect 301222 56692 301228 56704
rect 301096 56664 301228 56692
rect 301096 56652 301102 56664
rect 301222 56652 301228 56664
rect 301280 56652 301286 56704
rect 232314 56624 232320 56636
rect 232275 56596 232320 56624
rect 232314 56584 232320 56596
rect 232372 56584 232378 56636
rect 236270 56624 236276 56636
rect 236231 56596 236276 56624
rect 236270 56584 236276 56596
rect 236328 56584 236334 56636
rect 239030 56624 239036 56636
rect 238991 56596 239036 56624
rect 239030 56584 239036 56596
rect 239088 56584 239094 56636
rect 270770 56624 270776 56636
rect 270731 56596 270776 56624
rect 270770 56584 270776 56596
rect 270828 56584 270834 56636
rect 330113 56627 330171 56633
rect 330113 56593 330125 56627
rect 330159 56624 330171 56627
rect 330202 56624 330208 56636
rect 330159 56596 330208 56624
rect 330159 56593 330171 56596
rect 330113 56587 330171 56593
rect 330202 56584 330208 56596
rect 330260 56584 330266 56636
rect 336918 56624 336924 56636
rect 336879 56596 336924 56624
rect 336918 56584 336924 56596
rect 336976 56584 336982 56636
rect 357526 56584 357532 56636
rect 357584 56624 357590 56636
rect 357710 56624 357716 56636
rect 357584 56596 357716 56624
rect 357584 56584 357590 56596
rect 357710 56584 357716 56596
rect 357768 56584 357774 56636
rect 358630 56624 358636 56636
rect 358591 56596 358636 56624
rect 358630 56584 358636 56596
rect 358688 56584 358694 56636
rect 421190 56624 421196 56636
rect 421151 56596 421196 56624
rect 421190 56584 421196 56596
rect 421248 56584 421254 56636
rect 244550 56556 244556 56568
rect 244511 56528 244556 56556
rect 244550 56516 244556 56528
rect 244608 56516 244614 56568
rect 299658 56556 299664 56568
rect 299619 56528 299664 56556
rect 299658 56516 299664 56528
rect 299716 56516 299722 56568
rect 301038 56556 301044 56568
rect 300999 56528 301044 56556
rect 301038 56516 301044 56528
rect 301096 56516 301102 56568
rect 324774 56556 324780 56568
rect 324735 56528 324780 56556
rect 324774 56516 324780 56528
rect 324832 56516 324838 56568
rect 337286 56556 337292 56568
rect 337247 56528 337292 56556
rect 337286 56516 337292 56528
rect 337344 56516 337350 56568
rect 357526 56488 357532 56500
rect 357487 56460 357532 56488
rect 357526 56448 357532 56460
rect 357584 56448 357590 56500
rect 288710 55292 288716 55344
rect 288768 55332 288774 55344
rect 288768 55304 288940 55332
rect 288768 55292 288774 55304
rect 288912 55276 288940 55304
rect 288894 55224 288900 55276
rect 288952 55224 288958 55276
rect 317506 55224 317512 55276
rect 317564 55264 317570 55276
rect 317690 55264 317696 55276
rect 317564 55236 317696 55264
rect 317564 55224 317570 55236
rect 317690 55224 317696 55236
rect 317748 55224 317754 55276
rect 310882 55156 310888 55208
rect 310940 55196 310946 55208
rect 311066 55196 311072 55208
rect 310940 55168 311072 55196
rect 310940 55156 310946 55168
rect 311066 55156 311072 55168
rect 311124 55156 311130 55208
rect 239030 53184 239036 53236
rect 239088 53224 239094 53236
rect 239125 53227 239183 53233
rect 239125 53224 239137 53227
rect 239088 53196 239137 53224
rect 239088 53184 239094 53196
rect 239125 53193 239137 53196
rect 239171 53193 239183 53227
rect 239125 53187 239183 53193
rect 265158 53116 265164 53168
rect 265216 53156 265222 53168
rect 265342 53156 265348 53168
rect 265216 53128 265348 53156
rect 265216 53116 265222 53128
rect 265342 53116 265348 53128
rect 265400 53116 265406 53168
rect 247218 51116 247224 51128
rect 247144 51088 247224 51116
rect 247144 51060 247172 51088
rect 247218 51076 247224 51088
rect 247276 51076 247282 51128
rect 247126 51008 247132 51060
rect 247184 51008 247190 51060
rect 386414 51008 386420 51060
rect 386472 51048 386478 51060
rect 386598 51048 386604 51060
rect 386472 51020 386604 51048
rect 386472 51008 386478 51020
rect 386598 51008 386604 51020
rect 386656 51008 386662 51060
rect 273441 50983 273499 50989
rect 273441 50949 273453 50983
rect 273487 50980 273499 50983
rect 273530 50980 273536 50992
rect 273487 50952 273536 50980
rect 273487 50949 273499 50952
rect 273441 50943 273499 50949
rect 273530 50940 273536 50952
rect 273588 50940 273594 50992
rect 2774 50464 2780 50516
rect 2832 50504 2838 50516
rect 4798 50504 4804 50516
rect 2832 50476 4804 50504
rect 2832 50464 2838 50476
rect 4798 50464 4804 50476
rect 4856 50464 4862 50516
rect 286042 48396 286048 48408
rect 285968 48368 286048 48396
rect 285968 48340 285996 48368
rect 286042 48356 286048 48368
rect 286100 48356 286106 48408
rect 360470 48396 360476 48408
rect 360396 48368 360476 48396
rect 360396 48340 360424 48368
rect 360470 48356 360476 48368
rect 360528 48356 360534 48408
rect 239122 48328 239128 48340
rect 239083 48300 239128 48328
rect 239122 48288 239128 48300
rect 239180 48288 239186 48340
rect 267826 48288 267832 48340
rect 267884 48328 267890 48340
rect 267884 48300 267964 48328
rect 267884 48288 267890 48300
rect 236270 48260 236276 48272
rect 236231 48232 236276 48260
rect 236270 48220 236276 48232
rect 236328 48220 236334 48272
rect 250162 48220 250168 48272
rect 250220 48260 250226 48272
rect 250254 48260 250260 48272
rect 250220 48232 250260 48260
rect 250220 48220 250226 48232
rect 250254 48220 250260 48232
rect 250312 48220 250318 48272
rect 267936 48204 267964 48300
rect 284662 48288 284668 48340
rect 284720 48328 284726 48340
rect 284754 48328 284760 48340
rect 284720 48300 284760 48328
rect 284720 48288 284726 48300
rect 284754 48288 284760 48300
rect 284812 48288 284818 48340
rect 285950 48288 285956 48340
rect 286008 48288 286014 48340
rect 323302 48328 323308 48340
rect 323263 48300 323308 48328
rect 323302 48288 323308 48300
rect 323360 48288 323366 48340
rect 339770 48328 339776 48340
rect 339731 48300 339776 48328
rect 339770 48288 339776 48300
rect 339828 48288 339834 48340
rect 341242 48288 341248 48340
rect 341300 48328 341306 48340
rect 341426 48328 341432 48340
rect 341300 48300 341432 48328
rect 341300 48288 341306 48300
rect 341426 48288 341432 48300
rect 341484 48288 341490 48340
rect 358630 48288 358636 48340
rect 358688 48328 358694 48340
rect 358722 48328 358728 48340
rect 358688 48300 358728 48328
rect 358688 48288 358694 48300
rect 358722 48288 358728 48300
rect 358780 48288 358786 48340
rect 360378 48288 360384 48340
rect 360436 48288 360442 48340
rect 367002 48328 367008 48340
rect 366963 48300 367008 48328
rect 367002 48288 367008 48300
rect 367060 48288 367066 48340
rect 460014 48328 460020 48340
rect 459975 48300 460020 48328
rect 460014 48288 460020 48300
rect 460072 48288 460078 48340
rect 470594 48328 470600 48340
rect 470555 48300 470600 48328
rect 470594 48288 470600 48300
rect 470652 48288 470658 48340
rect 273530 48260 273536 48272
rect 273491 48232 273536 48260
rect 273530 48220 273536 48232
rect 273588 48220 273594 48272
rect 244550 48192 244556 48204
rect 244511 48164 244556 48192
rect 244550 48152 244556 48164
rect 244608 48152 244614 48204
rect 267918 48152 267924 48204
rect 267976 48152 267982 48204
rect 460014 48192 460020 48204
rect 459975 48164 460020 48192
rect 460014 48152 460020 48164
rect 460072 48152 460078 48204
rect 291378 46996 291384 47048
rect 291436 46996 291442 47048
rect 337194 46996 337200 47048
rect 337252 47036 337258 47048
rect 337289 47039 337347 47045
rect 337289 47036 337301 47039
rect 337252 47008 337301 47036
rect 337252 46996 337258 47008
rect 337289 47005 337301 47008
rect 337335 47005 337347 47039
rect 337289 46999 337347 47005
rect 266538 46928 266544 46980
rect 266596 46968 266602 46980
rect 266722 46968 266728 46980
rect 266596 46940 266728 46968
rect 266596 46928 266602 46940
rect 266722 46928 266728 46940
rect 266780 46928 266786 46980
rect 288710 46928 288716 46980
rect 288768 46968 288774 46980
rect 288894 46968 288900 46980
rect 288768 46940 288900 46968
rect 288768 46928 288774 46940
rect 288894 46928 288900 46940
rect 288952 46928 288958 46980
rect 291396 46968 291424 46996
rect 291470 46968 291476 46980
rect 291396 46940 291476 46968
rect 291470 46928 291476 46940
rect 291528 46928 291534 46980
rect 294230 46968 294236 46980
rect 294191 46940 294236 46968
rect 294230 46928 294236 46940
rect 294288 46928 294294 46980
rect 301038 46968 301044 46980
rect 300999 46940 301044 46968
rect 301038 46928 301044 46940
rect 301096 46928 301102 46980
rect 303798 46928 303804 46980
rect 303856 46968 303862 46980
rect 303890 46968 303896 46980
rect 303856 46940 303896 46968
rect 303856 46928 303862 46940
rect 303890 46928 303896 46940
rect 303948 46928 303954 46980
rect 306742 46928 306748 46980
rect 306800 46968 306806 46980
rect 306834 46968 306840 46980
rect 306800 46940 306840 46968
rect 306800 46928 306806 46940
rect 306834 46928 306840 46940
rect 306892 46928 306898 46980
rect 324590 46928 324596 46980
rect 324648 46968 324654 46980
rect 324777 46971 324835 46977
rect 324777 46968 324789 46971
rect 324648 46940 324789 46968
rect 324648 46928 324654 46940
rect 324777 46937 324789 46940
rect 324823 46937 324835 46971
rect 324777 46931 324835 46937
rect 357529 46971 357587 46977
rect 357529 46937 357541 46971
rect 357575 46968 357587 46971
rect 357618 46968 357624 46980
rect 357575 46940 357624 46968
rect 357575 46937 357587 46940
rect 357529 46931 357587 46937
rect 357618 46928 357624 46940
rect 357676 46928 357682 46980
rect 377214 46928 377220 46980
rect 377272 46968 377278 46980
rect 377306 46968 377312 46980
rect 377272 46940 377312 46968
rect 377272 46928 377278 46940
rect 377306 46928 377312 46940
rect 377364 46928 377370 46980
rect 244550 46900 244556 46912
rect 244511 46872 244556 46900
rect 244550 46860 244556 46872
rect 244608 46860 244614 46912
rect 262582 46860 262588 46912
rect 262640 46900 262646 46912
rect 262766 46900 262772 46912
rect 262640 46872 262772 46900
rect 262640 46860 262646 46872
rect 262766 46860 262772 46872
rect 262824 46860 262830 46912
rect 323302 46900 323308 46912
rect 323263 46872 323308 46900
rect 323302 46860 323308 46872
rect 323360 46860 323366 46912
rect 327258 46900 327264 46912
rect 327219 46872 327264 46900
rect 327258 46860 327264 46872
rect 327316 46860 327322 46912
rect 330110 46900 330116 46912
rect 330071 46872 330116 46900
rect 330110 46860 330116 46872
rect 330168 46860 330174 46912
rect 336918 46900 336924 46912
rect 336879 46872 336924 46900
rect 336918 46860 336924 46872
rect 336976 46860 336982 46912
rect 337194 46900 337200 46912
rect 337155 46872 337200 46900
rect 337194 46860 337200 46872
rect 337252 46860 337258 46912
rect 341245 46903 341303 46909
rect 341245 46869 341257 46903
rect 341291 46900 341303 46903
rect 341426 46900 341432 46912
rect 341291 46872 341432 46900
rect 341291 46869 341303 46872
rect 341245 46863 341303 46869
rect 341426 46860 341432 46872
rect 341484 46860 341490 46912
rect 358633 46903 358691 46909
rect 358633 46869 358645 46903
rect 358679 46900 358691 46903
rect 358722 46900 358728 46912
rect 358679 46872 358728 46900
rect 358679 46869 358691 46872
rect 358633 46863 358691 46869
rect 358722 46860 358728 46872
rect 358780 46860 358786 46912
rect 359001 46903 359059 46909
rect 359001 46869 359013 46903
rect 359047 46900 359059 46903
rect 359090 46900 359096 46912
rect 359047 46872 359096 46900
rect 359047 46869 359059 46872
rect 359001 46863 359059 46869
rect 359090 46860 359096 46872
rect 359148 46860 359154 46912
rect 367002 46900 367008 46912
rect 366963 46872 367008 46900
rect 367002 46860 367008 46872
rect 367060 46860 367066 46912
rect 421190 46900 421196 46912
rect 421151 46872 421196 46900
rect 421190 46860 421196 46872
rect 421248 46860 421254 46912
rect 357618 46832 357624 46844
rect 357579 46804 357624 46832
rect 357618 46792 357624 46804
rect 357676 46792 357682 46844
rect 299661 45611 299719 45617
rect 299661 45577 299673 45611
rect 299707 45608 299719 45611
rect 299750 45608 299756 45620
rect 299707 45580 299756 45608
rect 299707 45577 299719 45580
rect 299661 45571 299719 45577
rect 299750 45568 299756 45580
rect 299808 45568 299814 45620
rect 262766 45540 262772 45552
rect 262727 45512 262772 45540
rect 262766 45500 262772 45512
rect 262824 45500 262830 45552
rect 294230 45540 294236 45552
rect 294191 45512 294236 45540
rect 294230 45500 294236 45512
rect 294288 45500 294294 45552
rect 310882 45500 310888 45552
rect 310940 45540 310946 45552
rect 311066 45540 311072 45552
rect 310940 45512 311072 45540
rect 310940 45500 310946 45512
rect 311066 45500 311072 45512
rect 311124 45500 311130 45552
rect 317506 45500 317512 45552
rect 317564 45540 317570 45552
rect 317690 45540 317696 45552
rect 317564 45512 317696 45540
rect 317564 45500 317570 45512
rect 317690 45500 317696 45512
rect 317748 45500 317754 45552
rect 299750 45432 299756 45484
rect 299808 45472 299814 45484
rect 299842 45472 299848 45484
rect 299808 45444 299848 45472
rect 299808 45432 299814 45444
rect 299842 45432 299848 45444
rect 299900 45432 299906 45484
rect 284662 44684 284668 44736
rect 284720 44724 284726 44736
rect 284757 44727 284815 44733
rect 284757 44724 284769 44727
rect 284720 44696 284769 44724
rect 284720 44684 284726 44696
rect 284757 44693 284769 44696
rect 284803 44693 284815 44727
rect 284757 44687 284815 44693
rect 239033 42075 239091 42081
rect 239033 42041 239045 42075
rect 239079 42072 239091 42075
rect 239122 42072 239128 42084
rect 239079 42044 239128 42072
rect 239079 42041 239091 42044
rect 239033 42035 239091 42041
rect 239122 42032 239128 42044
rect 239180 42032 239186 42084
rect 360286 41352 360292 41404
rect 360344 41392 360350 41404
rect 360470 41392 360476 41404
rect 360344 41364 360476 41392
rect 360344 41352 360350 41364
rect 360470 41352 360476 41364
rect 360528 41352 360534 41404
rect 460017 41395 460075 41401
rect 460017 41361 460029 41395
rect 460063 41392 460075 41395
rect 460198 41392 460204 41404
rect 460063 41364 460204 41392
rect 460063 41361 460075 41364
rect 460017 41355 460075 41361
rect 460198 41352 460204 41364
rect 460256 41352 460262 41404
rect 367094 40196 367100 40248
rect 367152 40236 367158 40248
rect 376662 40236 376668 40248
rect 367152 40208 376668 40236
rect 367152 40196 367158 40208
rect 376662 40196 376668 40208
rect 376720 40196 376726 40248
rect 417878 40196 417884 40248
rect 417936 40236 417942 40248
rect 420362 40236 420368 40248
rect 417936 40208 420368 40236
rect 417936 40196 417942 40208
rect 420362 40196 420368 40208
rect 420420 40196 420426 40248
rect 437198 40196 437204 40248
rect 437256 40236 437262 40248
rect 437474 40236 437480 40248
rect 437256 40208 437480 40236
rect 437256 40196 437262 40208
rect 437474 40196 437480 40208
rect 437532 40196 437538 40248
rect 456518 40196 456524 40248
rect 456576 40236 456582 40248
rect 456886 40236 456892 40248
rect 456576 40208 456892 40236
rect 456576 40196 456582 40208
rect 456886 40196 456892 40208
rect 456944 40196 456950 40248
rect 306374 40128 306380 40180
rect 306432 40168 306438 40180
rect 315942 40168 315948 40180
rect 306432 40140 315948 40168
rect 306432 40128 306438 40140
rect 315942 40128 315948 40140
rect 316000 40128 316006 40180
rect 232314 38632 232320 38684
rect 232372 38672 232378 38684
rect 236270 38672 236276 38684
rect 232372 38644 232544 38672
rect 236231 38644 236276 38672
rect 232372 38632 232378 38644
rect 232516 38548 232544 38644
rect 236270 38632 236276 38644
rect 236328 38632 236334 38684
rect 247126 38632 247132 38684
rect 247184 38672 247190 38684
rect 247218 38672 247224 38684
rect 247184 38644 247224 38672
rect 247184 38632 247190 38644
rect 247218 38632 247224 38644
rect 247276 38632 247282 38684
rect 270770 38632 270776 38684
rect 270828 38672 270834 38684
rect 270862 38672 270868 38684
rect 270828 38644 270868 38672
rect 270828 38632 270834 38644
rect 270862 38632 270868 38644
rect 270920 38632 270926 38684
rect 272150 38632 272156 38684
rect 272208 38672 272214 38684
rect 272242 38672 272248 38684
rect 272208 38644 272248 38672
rect 272208 38632 272214 38644
rect 272242 38632 272248 38644
rect 272300 38632 272306 38684
rect 273530 38672 273536 38684
rect 273491 38644 273536 38672
rect 273530 38632 273536 38644
rect 273588 38632 273594 38684
rect 296806 38632 296812 38684
rect 296864 38632 296870 38684
rect 301038 38632 301044 38684
rect 301096 38632 301102 38684
rect 302510 38632 302516 38684
rect 302568 38672 302574 38684
rect 302602 38672 302608 38684
rect 302568 38644 302608 38672
rect 302568 38632 302574 38644
rect 302602 38632 302608 38644
rect 302660 38632 302666 38684
rect 232498 38496 232504 38548
rect 232556 38496 232562 38548
rect 236270 38536 236276 38548
rect 236231 38508 236276 38536
rect 236270 38496 236276 38508
rect 236328 38496 236334 38548
rect 296824 38536 296852 38632
rect 301056 38604 301084 38632
rect 301314 38604 301320 38616
rect 301056 38576 301320 38604
rect 301314 38564 301320 38576
rect 301372 38564 301378 38616
rect 303798 38604 303804 38616
rect 303759 38576 303804 38604
rect 303798 38564 303804 38576
rect 303856 38564 303862 38616
rect 306742 38564 306748 38616
rect 306800 38604 306806 38616
rect 306834 38604 306840 38616
rect 306800 38576 306840 38604
rect 306800 38564 306806 38576
rect 306834 38564 306840 38576
rect 306892 38564 306898 38616
rect 377122 38564 377128 38616
rect 377180 38604 377186 38616
rect 377306 38604 377312 38616
rect 377180 38576 377312 38604
rect 377180 38564 377186 38576
rect 377306 38564 377312 38576
rect 377364 38564 377370 38616
rect 296898 38536 296904 38548
rect 296824 38508 296904 38536
rect 296898 38496 296904 38508
rect 296956 38496 296962 38548
rect 250254 38156 250260 38208
rect 250312 38156 250318 38208
rect 250272 38072 250300 38156
rect 250254 38020 250260 38072
rect 250312 38020 250318 38072
rect 337194 37380 337200 37392
rect 337155 37352 337200 37380
rect 337194 37340 337200 37352
rect 337252 37340 337258 37392
rect 244550 37312 244556 37324
rect 244511 37284 244556 37312
rect 244550 37272 244556 37284
rect 244608 37272 244614 37324
rect 266538 37272 266544 37324
rect 266596 37312 266602 37324
rect 266630 37312 266636 37324
rect 266596 37284 266636 37312
rect 266596 37272 266602 37284
rect 266630 37272 266636 37284
rect 266688 37272 266694 37324
rect 323305 37315 323363 37321
rect 323305 37281 323317 37315
rect 323351 37312 323363 37315
rect 323394 37312 323400 37324
rect 323351 37284 323400 37312
rect 323351 37281 323363 37284
rect 323305 37275 323363 37281
rect 323394 37272 323400 37284
rect 323452 37272 323458 37324
rect 327258 37312 327264 37324
rect 327219 37284 327264 37312
rect 327258 37272 327264 37284
rect 327316 37272 327322 37324
rect 330110 37312 330116 37324
rect 330071 37284 330116 37312
rect 330110 37272 330116 37284
rect 330168 37272 330174 37324
rect 336918 37312 336924 37324
rect 336879 37284 336924 37312
rect 336918 37272 336924 37284
rect 336976 37272 336982 37324
rect 341242 37312 341248 37324
rect 341203 37284 341248 37312
rect 341242 37272 341248 37284
rect 341300 37272 341306 37324
rect 357618 37312 357624 37324
rect 357579 37284 357624 37312
rect 357618 37272 357624 37284
rect 357676 37272 357682 37324
rect 358630 37312 358636 37324
rect 358591 37284 358636 37312
rect 358630 37272 358636 37284
rect 358688 37272 358694 37324
rect 358998 37312 359004 37324
rect 358959 37284 359004 37312
rect 358998 37272 359004 37284
rect 359056 37272 359062 37324
rect 367002 37312 367008 37324
rect 366963 37284 367008 37312
rect 367002 37272 367008 37284
rect 367060 37272 367066 37324
rect 421190 37312 421196 37324
rect 421151 37284 421196 37312
rect 421190 37272 421196 37284
rect 421248 37272 421254 37324
rect 251174 37204 251180 37256
rect 251232 37244 251238 37256
rect 251450 37244 251456 37256
rect 251232 37216 251456 37244
rect 251232 37204 251238 37216
rect 251450 37204 251456 37216
rect 251508 37204 251514 37256
rect 259730 37244 259736 37256
rect 259691 37216 259736 37244
rect 259730 37204 259736 37216
rect 259788 37204 259794 37256
rect 267829 37247 267887 37253
rect 267829 37213 267841 37247
rect 267875 37244 267887 37247
rect 267918 37244 267924 37256
rect 267875 37216 267924 37244
rect 267875 37213 267887 37216
rect 267829 37207 267887 37213
rect 267918 37204 267924 37216
rect 267976 37204 267982 37256
rect 272242 37204 272248 37256
rect 272300 37244 272306 37256
rect 272334 37244 272340 37256
rect 272300 37216 272340 37244
rect 272300 37204 272306 37216
rect 272334 37204 272340 37216
rect 272392 37204 272398 37256
rect 288710 37204 288716 37256
rect 288768 37204 288774 37256
rect 337194 37204 337200 37256
rect 337252 37244 337258 37256
rect 337286 37244 337292 37256
rect 337252 37216 337292 37244
rect 337252 37204 337258 37216
rect 337286 37204 337292 37216
rect 337344 37204 337350 37256
rect 288728 37176 288756 37204
rect 288802 37176 288808 37188
rect 288728 37148 288808 37176
rect 288802 37136 288808 37148
rect 288860 37136 288866 37188
rect 262766 35952 262772 35964
rect 262727 35924 262772 35952
rect 262766 35912 262772 35924
rect 262824 35912 262830 35964
rect 3142 35844 3148 35896
rect 3200 35884 3206 35896
rect 6178 35884 6184 35896
rect 3200 35856 6184 35884
rect 3200 35844 3206 35856
rect 6178 35844 6184 35856
rect 6236 35844 6242 35896
rect 272245 35887 272303 35893
rect 272245 35853 272257 35887
rect 272291 35884 272303 35887
rect 272334 35884 272340 35896
rect 272291 35856 272340 35884
rect 272291 35853 272303 35856
rect 272245 35847 272303 35853
rect 272334 35844 272340 35856
rect 272392 35844 272398 35896
rect 301133 35887 301191 35893
rect 301133 35853 301145 35887
rect 301179 35884 301191 35887
rect 301314 35884 301320 35896
rect 301179 35856 301320 35884
rect 301179 35853 301191 35856
rect 301133 35847 301191 35853
rect 301314 35844 301320 35856
rect 301372 35844 301378 35896
rect 310885 35887 310943 35893
rect 310885 35853 310897 35887
rect 310931 35884 310943 35887
rect 311066 35884 311072 35896
rect 310931 35856 311072 35884
rect 310931 35853 310943 35856
rect 310885 35847 310943 35853
rect 311066 35844 311072 35856
rect 311124 35844 311130 35896
rect 358998 34076 359004 34128
rect 359056 34076 359062 34128
rect 359016 34048 359044 34076
rect 359090 34048 359096 34060
rect 359016 34020 359096 34048
rect 359090 34008 359096 34020
rect 359148 34008 359154 34060
rect 336734 33804 336740 33856
rect 336792 33844 336798 33856
rect 336918 33844 336924 33856
rect 336792 33816 336924 33844
rect 336792 33804 336798 33816
rect 336918 33804 336924 33816
rect 336976 33804 336982 33856
rect 303801 32419 303859 32425
rect 303801 32385 303813 32419
rect 303847 32416 303859 32419
rect 303890 32416 303896 32428
rect 303847 32388 303896 32416
rect 303847 32385 303859 32388
rect 303801 32379 303859 32385
rect 303890 32376 303896 32388
rect 303948 32376 303954 32428
rect 357618 32376 357624 32428
rect 357676 32416 357682 32428
rect 357802 32416 357808 32428
rect 357676 32388 357808 32416
rect 357676 32376 357682 32388
rect 357802 32376 357808 32388
rect 357860 32376 357866 32428
rect 341242 32280 341248 32292
rect 341203 32252 341248 32280
rect 341242 32240 341248 32252
rect 341300 32240 341306 32292
rect 317506 31764 317512 31816
rect 317564 31804 317570 31816
rect 317690 31804 317696 31816
rect 317564 31776 317696 31804
rect 317564 31764 317570 31776
rect 317690 31764 317696 31776
rect 317748 31764 317754 31816
rect 327258 31764 327264 31816
rect 327316 31764 327322 31816
rect 377122 31764 377128 31816
rect 377180 31764 377186 31816
rect 386506 31764 386512 31816
rect 386564 31764 386570 31816
rect 236273 31671 236331 31677
rect 236273 31637 236285 31671
rect 236319 31668 236331 31671
rect 236362 31668 236368 31680
rect 236319 31640 236368 31668
rect 236319 31637 236331 31640
rect 236273 31631 236331 31637
rect 236362 31628 236368 31640
rect 236420 31628 236426 31680
rect 327276 31612 327304 31764
rect 377140 31680 377168 31764
rect 377122 31628 377128 31680
rect 377180 31628 377186 31680
rect 386524 31668 386552 31764
rect 386598 31668 386604 31680
rect 386524 31640 386604 31668
rect 386598 31628 386604 31640
rect 386656 31628 386662 31680
rect 327258 31560 327264 31612
rect 327316 31560 327322 31612
rect 278774 29248 278780 29300
rect 278832 29288 278838 29300
rect 281258 29288 281264 29300
rect 278832 29260 281264 29288
rect 278832 29248 278838 29260
rect 281258 29248 281264 29260
rect 281316 29248 281322 29300
rect 367094 29180 367100 29232
rect 367152 29220 367158 29232
rect 376662 29220 376668 29232
rect 367152 29192 376668 29220
rect 367152 29180 367158 29192
rect 376662 29180 376668 29192
rect 376720 29180 376726 29232
rect 240134 29112 240140 29164
rect 240192 29152 240198 29164
rect 249702 29152 249708 29164
rect 240192 29124 249708 29152
rect 240192 29112 240198 29124
rect 249702 29112 249708 29124
rect 249760 29112 249766 29164
rect 367002 29112 367008 29164
rect 367060 29112 367066 29164
rect 437198 29112 437204 29164
rect 437256 29152 437262 29164
rect 437474 29152 437480 29164
rect 437256 29124 437480 29152
rect 437256 29112 437262 29124
rect 437474 29112 437480 29124
rect 437532 29112 437538 29164
rect 456518 29112 456524 29164
rect 456576 29152 456582 29164
rect 456794 29152 456800 29164
rect 456576 29124 456800 29152
rect 456576 29112 456582 29124
rect 456794 29112 456800 29124
rect 456852 29112 456858 29164
rect 302510 29044 302516 29096
rect 302568 29044 302574 29096
rect 341242 29084 341248 29096
rect 341203 29056 341248 29084
rect 341242 29044 341248 29056
rect 341300 29044 341306 29096
rect 347774 29044 347780 29096
rect 347832 29084 347838 29096
rect 357342 29084 357348 29096
rect 347832 29056 357348 29084
rect 347832 29044 347838 29056
rect 357342 29044 357348 29056
rect 357400 29044 357406 29096
rect 239030 29016 239036 29028
rect 238991 28988 239036 29016
rect 239030 28976 239036 28988
rect 239088 28976 239094 29028
rect 284754 29016 284760 29028
rect 284715 28988 284760 29016
rect 284754 28976 284760 28988
rect 284812 28976 284818 29028
rect 285950 28976 285956 29028
rect 286008 29016 286014 29028
rect 286042 29016 286048 29028
rect 286008 28988 286048 29016
rect 286008 28976 286014 28988
rect 286042 28976 286048 28988
rect 286100 28976 286106 29028
rect 302528 28960 302556 29044
rect 367020 29028 367048 29112
rect 492766 29044 492772 29096
rect 492824 29084 492830 29096
rect 502242 29084 502248 29096
rect 492824 29056 502248 29084
rect 492824 29044 492830 29056
rect 502242 29044 502248 29056
rect 502300 29044 502306 29096
rect 325970 28976 325976 29028
rect 326028 29016 326034 29028
rect 326062 29016 326068 29028
rect 326028 28988 326068 29016
rect 326028 28976 326034 28988
rect 326062 28976 326068 28988
rect 326120 28976 326126 29028
rect 358630 28976 358636 29028
rect 358688 29016 358694 29028
rect 358722 29016 358728 29028
rect 358688 28988 358728 29016
rect 358688 28976 358694 28988
rect 358722 28976 358728 28988
rect 358780 28976 358786 29028
rect 367002 28976 367008 29028
rect 367060 28976 367066 29028
rect 232222 28908 232228 28960
rect 232280 28948 232286 28960
rect 232406 28948 232412 28960
rect 232280 28920 232412 28948
rect 232280 28908 232286 28920
rect 232406 28908 232412 28920
rect 232464 28908 232470 28960
rect 236362 28948 236368 28960
rect 236323 28920 236368 28948
rect 236362 28908 236368 28920
rect 236420 28908 236426 28960
rect 291470 28908 291476 28960
rect 291528 28948 291534 28960
rect 291654 28948 291660 28960
rect 291528 28920 291660 28948
rect 291528 28908 291534 28920
rect 291654 28908 291660 28920
rect 291712 28908 291718 28960
rect 295518 28908 295524 28960
rect 295576 28948 295582 28960
rect 295610 28948 295616 28960
rect 295576 28920 295616 28948
rect 295576 28908 295582 28920
rect 295610 28908 295616 28920
rect 295668 28908 295674 28960
rect 302510 28908 302516 28960
rect 302568 28908 302574 28960
rect 323302 28908 323308 28960
rect 323360 28948 323366 28960
rect 323394 28948 323400 28960
rect 323360 28920 323400 28948
rect 323360 28908 323366 28920
rect 323394 28908 323400 28920
rect 323452 28908 323458 28960
rect 324590 28908 324596 28960
rect 324648 28948 324654 28960
rect 324682 28948 324688 28960
rect 324648 28920 324688 28948
rect 324648 28908 324654 28920
rect 324682 28908 324688 28920
rect 324740 28908 324746 28960
rect 306374 28840 306380 28892
rect 306432 28880 306438 28892
rect 315942 28880 315948 28892
rect 306432 28852 315948 28880
rect 306432 28840 306438 28852
rect 315942 28840 315948 28852
rect 316000 28840 316006 28892
rect 267826 28608 267832 28620
rect 267787 28580 267832 28608
rect 267826 28568 267832 28580
rect 267884 28568 267890 28620
rect 259730 27656 259736 27668
rect 259691 27628 259736 27656
rect 259730 27616 259736 27628
rect 259788 27616 259794 27668
rect 247126 27588 247132 27600
rect 247087 27560 247132 27588
rect 247126 27548 247132 27560
rect 247184 27548 247190 27600
rect 249981 27591 250039 27597
rect 249981 27557 249993 27591
rect 250027 27588 250039 27591
rect 250162 27588 250168 27600
rect 250027 27560 250168 27588
rect 250027 27557 250039 27560
rect 249981 27551 250039 27557
rect 250162 27548 250168 27560
rect 250220 27548 250226 27600
rect 251358 27588 251364 27600
rect 251319 27560 251364 27588
rect 251358 27548 251364 27560
rect 251416 27548 251422 27600
rect 262582 27548 262588 27600
rect 262640 27588 262646 27600
rect 262674 27588 262680 27600
rect 262640 27560 262680 27588
rect 262640 27548 262646 27560
rect 262674 27548 262680 27560
rect 262732 27548 262738 27600
rect 265161 27591 265219 27597
rect 265161 27557 265173 27591
rect 265207 27588 265219 27591
rect 265250 27588 265256 27600
rect 265207 27560 265256 27588
rect 265207 27557 265219 27560
rect 265161 27551 265219 27557
rect 265250 27548 265256 27560
rect 265308 27548 265314 27600
rect 284754 27588 284760 27600
rect 284715 27560 284760 27588
rect 284754 27548 284760 27560
rect 284812 27548 284818 27600
rect 285953 27591 286011 27597
rect 285953 27557 285965 27591
rect 285999 27588 286011 27591
rect 286042 27588 286048 27600
rect 285999 27560 286048 27588
rect 285999 27557 286011 27560
rect 285953 27551 286011 27557
rect 286042 27548 286048 27560
rect 286100 27548 286106 27600
rect 341150 27548 341156 27600
rect 341208 27588 341214 27600
rect 341245 27591 341303 27597
rect 341245 27588 341257 27591
rect 341208 27560 341257 27588
rect 341208 27548 341214 27560
rect 341245 27557 341257 27560
rect 341291 27557 341303 27591
rect 357618 27588 357624 27600
rect 357579 27560 357624 27588
rect 341245 27551 341303 27557
rect 357618 27548 357624 27560
rect 357676 27548 357682 27600
rect 358541 27591 358599 27597
rect 358541 27557 358553 27591
rect 358587 27588 358599 27591
rect 358722 27588 358728 27600
rect 358587 27560 358728 27588
rect 358587 27557 358599 27560
rect 358541 27551 358599 27557
rect 358722 27548 358728 27560
rect 358780 27548 358786 27600
rect 359090 27548 359096 27600
rect 359148 27588 359154 27600
rect 359182 27588 359188 27600
rect 359148 27560 359188 27588
rect 359148 27548 359154 27560
rect 359182 27548 359188 27560
rect 359240 27548 359246 27600
rect 366821 27591 366879 27597
rect 366821 27557 366833 27591
rect 366867 27588 366879 27591
rect 367002 27588 367008 27600
rect 366867 27560 367008 27588
rect 366867 27557 366879 27560
rect 366821 27551 366879 27557
rect 367002 27548 367008 27560
rect 367060 27548 367066 27600
rect 421190 27588 421196 27600
rect 421151 27560 421196 27588
rect 421190 27548 421196 27560
rect 421248 27548 421254 27600
rect 272242 26296 272248 26308
rect 272203 26268 272248 26296
rect 272242 26256 272248 26268
rect 272300 26256 272306 26308
rect 294233 26299 294291 26305
rect 294233 26265 294245 26299
rect 294279 26296 294291 26299
rect 294414 26296 294420 26308
rect 294279 26268 294420 26296
rect 294279 26265 294291 26268
rect 294233 26259 294291 26265
rect 294414 26256 294420 26268
rect 294472 26256 294478 26308
rect 301130 26296 301136 26308
rect 301091 26268 301136 26296
rect 301130 26256 301136 26268
rect 301188 26256 301194 26308
rect 310882 26296 310888 26308
rect 310843 26268 310888 26296
rect 310882 26256 310888 26268
rect 310940 26256 310946 26308
rect 386233 26231 386291 26237
rect 386233 26197 386245 26231
rect 386279 26228 386291 26231
rect 386598 26228 386604 26240
rect 386279 26200 386604 26228
rect 386279 26197 386291 26200
rect 386233 26191 386291 26197
rect 386598 26188 386604 26200
rect 386656 26188 386662 26240
rect 271874 26120 271880 26172
rect 271932 26160 271938 26172
rect 272242 26160 272248 26172
rect 271932 26132 272248 26160
rect 271932 26120 271938 26132
rect 272242 26120 272248 26132
rect 272300 26120 272306 26172
rect 236365 22763 236423 22769
rect 236365 22729 236377 22763
rect 236411 22760 236423 22763
rect 236454 22760 236460 22772
rect 236411 22732 236460 22760
rect 236411 22729 236423 22732
rect 236365 22723 236423 22729
rect 236454 22720 236460 22732
rect 236512 22720 236518 22772
rect 270497 22151 270555 22157
rect 270497 22117 270509 22151
rect 270543 22148 270555 22151
rect 270770 22148 270776 22160
rect 270543 22120 270776 22148
rect 270543 22117 270555 22120
rect 270497 22111 270555 22117
rect 270770 22108 270776 22120
rect 270828 22108 270834 22160
rect 310790 22108 310796 22160
rect 310848 22148 310854 22160
rect 310885 22151 310943 22157
rect 310885 22148 310897 22151
rect 310848 22120 310897 22148
rect 310848 22108 310854 22120
rect 310885 22117 310897 22120
rect 310931 22117 310943 22151
rect 377122 22148 377128 22160
rect 310885 22111 310943 22117
rect 377048 22120 377128 22148
rect 377048 22092 377076 22120
rect 377122 22108 377128 22120
rect 377180 22108 377186 22160
rect 377030 22040 377036 22092
rect 377088 22040 377094 22092
rect 291562 19932 291568 19984
rect 291620 19932 291626 19984
rect 291580 19848 291608 19932
rect 291562 19796 291568 19848
rect 291620 19796 291626 19848
rect 306742 19320 306748 19372
rect 306800 19360 306806 19372
rect 306834 19360 306840 19372
rect 306800 19332 306840 19360
rect 306800 19320 306806 19332
rect 306834 19320 306840 19332
rect 306892 19320 306898 19372
rect 336734 19320 336740 19372
rect 336792 19360 336798 19372
rect 336918 19360 336924 19372
rect 336792 19332 336924 19360
rect 336792 19320 336798 19332
rect 336918 19320 336924 19332
rect 336976 19320 336982 19372
rect 251358 19292 251364 19304
rect 251319 19264 251364 19292
rect 251358 19252 251364 19264
rect 251416 19252 251422 19304
rect 325970 19252 325976 19304
rect 326028 19252 326034 19304
rect 327258 19252 327264 19304
rect 327316 19252 327322 19304
rect 470594 19292 470600 19304
rect 470555 19264 470600 19292
rect 470594 19252 470600 19264
rect 470652 19252 470658 19304
rect 325988 19168 326016 19252
rect 327276 19168 327304 19252
rect 325970 19116 325976 19168
rect 326028 19116 326034 19168
rect 327258 19116 327264 19168
rect 327316 19116 327322 19168
rect 337105 18479 337163 18485
rect 337105 18445 337117 18479
rect 337151 18476 337163 18479
rect 337286 18476 337292 18488
rect 337151 18448 337292 18476
rect 337151 18445 337163 18448
rect 337105 18439 337163 18445
rect 337286 18436 337292 18448
rect 337344 18436 337350 18488
rect 247126 18000 247132 18012
rect 247087 17972 247132 18000
rect 247126 17960 247132 17972
rect 247184 17960 247190 18012
rect 249978 18000 249984 18012
rect 249939 17972 249984 18000
rect 249978 17960 249984 17972
rect 250036 17960 250042 18012
rect 265158 18000 265164 18012
rect 265119 17972 265164 18000
rect 265158 17960 265164 17972
rect 265216 17960 265222 18012
rect 270586 17960 270592 18012
rect 270644 17960 270650 18012
rect 271966 17960 271972 18012
rect 272024 17960 272030 18012
rect 284754 18000 284760 18012
rect 284715 17972 284760 18000
rect 284754 17960 284760 17972
rect 284812 17960 284818 18012
rect 285950 18000 285956 18012
rect 285911 17972 285956 18000
rect 285950 17960 285956 17972
rect 286008 17960 286014 18012
rect 337102 18000 337108 18012
rect 337063 17972 337108 18000
rect 337102 17960 337108 17972
rect 337160 17960 337166 18012
rect 357621 18003 357679 18009
rect 357621 17969 357633 18003
rect 357667 18000 357679 18003
rect 357710 18000 357716 18012
rect 357667 17972 357716 18000
rect 357667 17969 357679 17972
rect 357621 17963 357679 17969
rect 357710 17960 357716 17972
rect 357768 17960 357774 18012
rect 236273 17935 236331 17941
rect 236273 17901 236285 17935
rect 236319 17932 236331 17935
rect 236454 17932 236460 17944
rect 236319 17904 236460 17932
rect 236319 17901 236331 17904
rect 236273 17895 236331 17901
rect 236454 17892 236460 17904
rect 236512 17892 236518 17944
rect 244369 17935 244427 17941
rect 244369 17901 244381 17935
rect 244415 17932 244427 17935
rect 244550 17932 244556 17944
rect 244415 17904 244556 17932
rect 244415 17901 244427 17904
rect 244369 17895 244427 17901
rect 244550 17892 244556 17904
rect 244608 17892 244614 17944
rect 270494 17932 270500 17944
rect 270455 17904 270500 17932
rect 270494 17892 270500 17904
rect 270552 17892 270558 17944
rect 270604 17876 270632 17960
rect 271984 17876 272012 17960
rect 273438 17932 273444 17944
rect 273399 17904 273444 17932
rect 273438 17892 273444 17904
rect 273496 17892 273502 17944
rect 270586 17824 270592 17876
rect 270644 17824 270650 17876
rect 271966 17824 271972 17876
rect 272024 17824 272030 17876
rect 347774 16872 347780 16924
rect 347832 16912 347838 16924
rect 352650 16912 352656 16924
rect 347832 16884 352656 16912
rect 347832 16872 347838 16884
rect 352650 16872 352656 16884
rect 352708 16872 352714 16924
rect 456518 16872 456524 16924
rect 456576 16912 456582 16924
rect 457438 16912 457444 16924
rect 456576 16884 457444 16912
rect 456576 16872 456582 16884
rect 457438 16872 457444 16884
rect 457496 16872 457502 16924
rect 369670 16804 369676 16856
rect 369728 16844 369734 16856
rect 376662 16844 376668 16856
rect 369728 16816 376668 16844
rect 369728 16804 369734 16816
rect 376662 16804 376668 16816
rect 376720 16804 376726 16856
rect 475562 16804 475568 16856
rect 475620 16844 475626 16856
rect 482922 16844 482928 16856
rect 475620 16816 482928 16844
rect 475620 16804 475626 16816
rect 482922 16804 482928 16816
rect 482980 16804 482986 16856
rect 437198 16736 437204 16788
rect 437256 16776 437262 16788
rect 437474 16776 437480 16788
rect 437256 16748 437480 16776
rect 437256 16736 437262 16748
rect 437474 16736 437480 16748
rect 437532 16736 437538 16788
rect 320818 16668 320824 16720
rect 320876 16708 320882 16720
rect 325602 16708 325608 16720
rect 320876 16680 325608 16708
rect 320876 16668 320882 16680
rect 325602 16668 325608 16680
rect 325660 16668 325666 16720
rect 386230 16640 386236 16652
rect 386191 16612 386236 16640
rect 386230 16600 386236 16612
rect 386288 16600 386294 16652
rect 278774 16532 278780 16584
rect 278832 16572 278838 16584
rect 290550 16572 290556 16584
rect 278832 16544 290556 16572
rect 278832 16532 278838 16544
rect 290550 16532 290556 16544
rect 290608 16532 290614 16584
rect 310882 15212 310888 15224
rect 310843 15184 310888 15212
rect 310882 15172 310888 15184
rect 310940 15172 310946 15224
rect 110322 15104 110328 15156
rect 110380 15144 110386 15156
rect 274726 15144 274732 15156
rect 110380 15116 274732 15144
rect 110380 15104 110386 15116
rect 274726 15104 274732 15116
rect 274784 15104 274790 15156
rect 107470 15036 107476 15088
rect 107528 15076 107534 15088
rect 273346 15076 273352 15088
rect 107528 15048 273352 15076
rect 107528 15036 107534 15048
rect 273346 15036 273352 15048
rect 273404 15036 273410 15088
rect 103422 14968 103428 15020
rect 103480 15008 103486 15020
rect 271966 15008 271972 15020
rect 103480 14980 271972 15008
rect 103480 14968 103486 14980
rect 271966 14968 271972 14980
rect 272024 14968 272030 15020
rect 99282 14900 99288 14952
rect 99340 14940 99346 14952
rect 270586 14940 270592 14952
rect 99340 14912 270592 14940
rect 99340 14900 99346 14912
rect 270586 14900 270592 14912
rect 270644 14900 270650 14952
rect 96522 14832 96528 14884
rect 96580 14872 96586 14884
rect 269206 14872 269212 14884
rect 96580 14844 269212 14872
rect 96580 14832 96586 14844
rect 269206 14832 269212 14844
rect 269264 14832 269270 14884
rect 92382 14764 92388 14816
rect 92440 14804 92446 14816
rect 266446 14804 266452 14816
rect 92440 14776 266452 14804
rect 92440 14764 92446 14776
rect 266446 14764 266452 14776
rect 266504 14764 266510 14816
rect 89622 14696 89628 14748
rect 89680 14736 89686 14748
rect 265066 14736 265072 14748
rect 89680 14708 265072 14736
rect 89680 14696 89686 14708
rect 265066 14696 265072 14708
rect 265124 14696 265130 14748
rect 85482 14628 85488 14680
rect 85540 14668 85546 14680
rect 263686 14668 263692 14680
rect 85540 14640 263692 14668
rect 85540 14628 85546 14640
rect 263686 14628 263692 14640
rect 263744 14628 263750 14680
rect 82722 14560 82728 14612
rect 82780 14600 82786 14612
rect 262582 14600 262588 14612
rect 82780 14572 262588 14600
rect 82780 14560 82786 14572
rect 262582 14560 262588 14572
rect 262640 14560 262646 14612
rect 78582 14492 78588 14544
rect 78640 14532 78646 14544
rect 260926 14532 260932 14544
rect 78640 14504 260932 14532
rect 78640 14492 78646 14504
rect 260926 14492 260932 14504
rect 260984 14492 260990 14544
rect 74442 14424 74448 14476
rect 74500 14464 74506 14476
rect 259638 14464 259644 14476
rect 74500 14436 259644 14464
rect 74500 14424 74506 14436
rect 259638 14424 259644 14436
rect 259696 14424 259702 14476
rect 114462 14356 114468 14408
rect 114520 14396 114526 14408
rect 276106 14396 276112 14408
rect 114520 14368 276112 14396
rect 114520 14356 114526 14368
rect 276106 14356 276112 14368
rect 276164 14356 276170 14408
rect 117222 14288 117228 14340
rect 117280 14328 117286 14340
rect 277670 14328 277676 14340
rect 117280 14300 277676 14328
rect 117280 14288 117286 14300
rect 277670 14288 277676 14300
rect 277728 14288 277734 14340
rect 121362 14220 121368 14272
rect 121420 14260 121426 14272
rect 278866 14260 278872 14272
rect 121420 14232 278872 14260
rect 121420 14220 121426 14232
rect 278866 14220 278872 14232
rect 278924 14220 278930 14272
rect 125410 14152 125416 14204
rect 125468 14192 125474 14204
rect 280246 14192 280252 14204
rect 125468 14164 280252 14192
rect 125468 14152 125474 14164
rect 280246 14152 280252 14164
rect 280304 14152 280310 14204
rect 186222 13744 186228 13796
rect 186280 13784 186286 13796
rect 306558 13784 306564 13796
rect 186280 13756 306564 13784
rect 186280 13744 186286 13756
rect 306558 13744 306564 13756
rect 306616 13744 306622 13796
rect 183462 13676 183468 13728
rect 183520 13716 183526 13728
rect 303890 13716 303896 13728
rect 183520 13688 303896 13716
rect 183520 13676 183526 13688
rect 303890 13676 303896 13688
rect 303948 13676 303954 13728
rect 179322 13608 179328 13660
rect 179380 13648 179386 13660
rect 302602 13648 302608 13660
rect 179380 13620 302608 13648
rect 179380 13608 179386 13620
rect 302602 13608 302608 13620
rect 302660 13608 302666 13660
rect 176562 13540 176568 13592
rect 176620 13580 176626 13592
rect 301130 13580 301136 13592
rect 176620 13552 301136 13580
rect 176620 13540 176626 13552
rect 301130 13540 301136 13552
rect 301188 13540 301194 13592
rect 172422 13472 172428 13524
rect 172480 13512 172486 13524
rect 299750 13512 299756 13524
rect 172480 13484 299756 13512
rect 172480 13472 172486 13484
rect 299750 13472 299756 13484
rect 299808 13472 299814 13524
rect 168282 13404 168288 13456
rect 168340 13444 168346 13456
rect 298278 13444 298284 13456
rect 168340 13416 298284 13444
rect 168340 13404 168346 13416
rect 298278 13404 298284 13416
rect 298336 13404 298342 13456
rect 165522 13336 165528 13388
rect 165580 13376 165586 13388
rect 296898 13376 296904 13388
rect 165580 13348 296904 13376
rect 165580 13336 165586 13348
rect 296898 13336 296904 13348
rect 296956 13336 296962 13388
rect 160002 13268 160008 13320
rect 160060 13308 160066 13320
rect 294322 13308 294328 13320
rect 160060 13280 294328 13308
rect 160060 13268 160066 13280
rect 294322 13268 294328 13280
rect 294380 13268 294386 13320
rect 155862 13200 155868 13252
rect 155920 13240 155926 13252
rect 292758 13240 292764 13252
rect 155920 13212 292764 13240
rect 155920 13200 155926 13212
rect 292758 13200 292764 13212
rect 292816 13200 292822 13252
rect 71682 13132 71688 13184
rect 71740 13172 71746 13184
rect 258166 13172 258172 13184
rect 71740 13144 258172 13172
rect 71740 13132 71746 13144
rect 258166 13132 258172 13144
rect 258224 13132 258230 13184
rect 31662 13064 31668 13116
rect 31720 13104 31726 13116
rect 241606 13104 241612 13116
rect 31720 13076 241612 13104
rect 31720 13064 31726 13076
rect 241606 13064 241612 13076
rect 241664 13064 241670 13116
rect 190362 12996 190368 13048
rect 190420 13036 190426 13048
rect 307938 13036 307944 13048
rect 190420 13008 307944 13036
rect 190420 12996 190426 13008
rect 307938 12996 307944 13008
rect 307996 12996 308002 13048
rect 206922 12928 206928 12980
rect 206980 12968 206986 12980
rect 314838 12968 314844 12980
rect 206980 12940 314844 12968
rect 206980 12928 206986 12940
rect 314838 12928 314844 12940
rect 314896 12928 314902 12980
rect 211062 12860 211068 12912
rect 211120 12900 211126 12912
rect 316218 12900 316224 12912
rect 211120 12872 316224 12900
rect 211120 12860 211126 12872
rect 316218 12860 316224 12872
rect 316276 12860 316282 12912
rect 213822 12792 213828 12844
rect 213880 12832 213886 12844
rect 317598 12832 317604 12844
rect 213880 12804 317604 12832
rect 213880 12792 213886 12804
rect 317598 12792 317604 12804
rect 317656 12792 317662 12844
rect 217962 12724 217968 12776
rect 218020 12764 218026 12776
rect 318978 12764 318984 12776
rect 218020 12736 318984 12764
rect 218020 12724 218026 12736
rect 318978 12724 318984 12736
rect 319036 12724 319042 12776
rect 220722 12656 220728 12708
rect 220780 12696 220786 12708
rect 320266 12696 320272 12708
rect 220780 12668 320272 12696
rect 220780 12656 220786 12668
rect 320266 12656 320272 12668
rect 320324 12656 320330 12708
rect 224862 12588 224868 12640
rect 224920 12628 224926 12640
rect 321738 12628 321744 12640
rect 224920 12600 321744 12628
rect 224920 12588 224926 12600
rect 321738 12588 321744 12600
rect 321796 12588 321802 12640
rect 229002 12520 229008 12572
rect 229060 12560 229066 12572
rect 323118 12560 323124 12572
rect 229060 12532 323124 12560
rect 229060 12520 229066 12532
rect 323118 12520 323124 12532
rect 323176 12520 323182 12572
rect 295610 12492 295616 12504
rect 295571 12464 295616 12492
rect 295610 12452 295616 12464
rect 295668 12452 295674 12504
rect 366910 12452 366916 12504
rect 366968 12452 366974 12504
rect 173802 12384 173808 12436
rect 173860 12424 173866 12436
rect 300946 12424 300952 12436
rect 173860 12396 300952 12424
rect 173860 12384 173866 12396
rect 300946 12384 300952 12396
rect 301004 12384 301010 12436
rect 366928 12368 366956 12452
rect 426434 12384 426440 12436
rect 426492 12424 426498 12436
rect 427538 12424 427544 12436
rect 426492 12396 427544 12424
rect 426492 12384 426498 12396
rect 427538 12384 427544 12396
rect 427596 12384 427602 12436
rect 169662 12316 169668 12368
rect 169720 12356 169726 12368
rect 299566 12356 299572 12368
rect 169720 12328 299572 12356
rect 169720 12316 169726 12328
rect 299566 12316 299572 12328
rect 299624 12316 299630 12368
rect 366910 12316 366916 12368
rect 366968 12316 366974 12368
rect 386230 12316 386236 12368
rect 386288 12356 386294 12368
rect 386598 12356 386604 12368
rect 386288 12328 386604 12356
rect 386288 12316 386294 12328
rect 386598 12316 386604 12328
rect 386656 12316 386662 12368
rect 166902 12248 166908 12300
rect 166960 12288 166966 12300
rect 298186 12288 298192 12300
rect 166960 12260 298192 12288
rect 166960 12248 166966 12260
rect 298186 12248 298192 12260
rect 298244 12248 298250 12300
rect 162762 12180 162768 12232
rect 162820 12220 162826 12232
rect 295613 12223 295671 12229
rect 295613 12220 295625 12223
rect 162820 12192 295625 12220
rect 162820 12180 162826 12192
rect 295613 12189 295625 12192
rect 295659 12189 295671 12223
rect 295613 12183 295671 12189
rect 151722 12112 151728 12164
rect 151780 12152 151786 12164
rect 291562 12152 291568 12164
rect 151780 12124 291568 12152
rect 151780 12112 151786 12124
rect 291562 12112 291568 12124
rect 291620 12112 291626 12164
rect 148962 12044 148968 12096
rect 149020 12084 149026 12096
rect 289998 12084 290004 12096
rect 149020 12056 290004 12084
rect 149020 12044 149026 12056
rect 289998 12044 290004 12056
rect 290056 12044 290062 12096
rect 144822 11976 144828 12028
rect 144880 12016 144886 12028
rect 288802 12016 288808 12028
rect 144880 11988 288808 12016
rect 144880 11976 144886 11988
rect 288802 11976 288808 11988
rect 288860 11976 288866 12028
rect 142062 11908 142068 11960
rect 142120 11948 142126 11960
rect 287330 11948 287336 11960
rect 142120 11920 287336 11948
rect 142120 11908 142126 11920
rect 287330 11908 287336 11920
rect 287388 11908 287394 11960
rect 128262 11840 128268 11892
rect 128320 11880 128326 11892
rect 281534 11880 281540 11892
rect 128320 11852 281540 11880
rect 128320 11840 128326 11852
rect 281534 11840 281540 11852
rect 281592 11840 281598 11892
rect 284570 11840 284576 11892
rect 284628 11880 284634 11892
rect 284754 11880 284760 11892
rect 284628 11852 284760 11880
rect 284628 11840 284634 11852
rect 284754 11840 284760 11852
rect 284812 11840 284818 11892
rect 126882 11772 126888 11824
rect 126940 11812 126946 11824
rect 281626 11812 281632 11824
rect 126940 11784 281632 11812
rect 126940 11772 126946 11784
rect 281626 11772 281632 11784
rect 281684 11772 281690 11824
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 238938 11744 238944 11756
rect 23440 11716 238944 11744
rect 23440 11704 23446 11716
rect 238938 11704 238944 11716
rect 238996 11704 239002 11756
rect 176470 11636 176476 11688
rect 176528 11676 176534 11688
rect 302326 11676 302332 11688
rect 176528 11648 302332 11676
rect 176528 11636 176534 11648
rect 302326 11636 302332 11648
rect 302384 11636 302390 11688
rect 180702 11568 180708 11620
rect 180760 11608 180766 11620
rect 303706 11608 303712 11620
rect 180760 11580 303712 11608
rect 180760 11568 180766 11580
rect 303706 11568 303712 11580
rect 303764 11568 303770 11620
rect 184842 11500 184848 11552
rect 184900 11540 184906 11552
rect 305086 11540 305092 11552
rect 184900 11512 305092 11540
rect 184900 11500 184906 11512
rect 305086 11500 305092 11512
rect 305144 11500 305150 11552
rect 187602 11432 187608 11484
rect 187660 11472 187666 11484
rect 306466 11472 306472 11484
rect 187660 11444 306472 11472
rect 187660 11432 187666 11444
rect 306466 11432 306472 11444
rect 306524 11432 306530 11484
rect 191742 11364 191748 11416
rect 191800 11404 191806 11416
rect 308030 11404 308036 11416
rect 191800 11376 308036 11404
rect 191800 11364 191806 11376
rect 308030 11364 308036 11376
rect 308088 11364 308094 11416
rect 194502 11296 194508 11348
rect 194560 11336 194566 11348
rect 309410 11336 309416 11348
rect 194560 11308 309416 11336
rect 194560 11296 194566 11308
rect 309410 11296 309416 11308
rect 309468 11296 309474 11348
rect 198642 11228 198648 11280
rect 198700 11268 198706 11280
rect 310882 11268 310888 11280
rect 198700 11240 310888 11268
rect 198700 11228 198706 11240
rect 310882 11228 310888 11240
rect 310940 11228 310946 11280
rect 113082 10956 113088 11008
rect 113140 10996 113146 11008
rect 276014 10996 276020 11008
rect 113140 10968 276020 10996
rect 113140 10956 113146 10968
rect 276014 10956 276020 10968
rect 276072 10956 276078 11008
rect 108942 10888 108948 10940
rect 109000 10928 109006 10940
rect 273441 10931 273499 10937
rect 273441 10928 273453 10931
rect 109000 10900 273453 10928
rect 109000 10888 109006 10900
rect 273441 10897 273453 10900
rect 273487 10897 273499 10931
rect 273441 10891 273499 10897
rect 106182 10820 106188 10872
rect 106240 10860 106246 10872
rect 271874 10860 271880 10872
rect 106240 10832 271880 10860
rect 106240 10820 106246 10832
rect 271874 10820 271880 10832
rect 271932 10820 271938 10872
rect 102042 10752 102048 10804
rect 102100 10792 102106 10804
rect 270494 10792 270500 10804
rect 102100 10764 270500 10792
rect 102100 10752 102106 10764
rect 270494 10752 270500 10764
rect 270552 10752 270558 10804
rect 99190 10684 99196 10736
rect 99248 10724 99254 10736
rect 269298 10724 269304 10736
rect 99248 10696 269304 10724
rect 99248 10684 99254 10696
rect 269298 10684 269304 10696
rect 269356 10684 269362 10736
rect 95142 10616 95148 10668
rect 95200 10656 95206 10668
rect 267734 10656 267740 10668
rect 95200 10628 267740 10656
rect 95200 10616 95206 10628
rect 267734 10616 267740 10628
rect 267792 10616 267798 10668
rect 91002 10548 91008 10600
rect 91060 10588 91066 10600
rect 266538 10588 266544 10600
rect 91060 10560 266544 10588
rect 91060 10548 91066 10560
rect 266538 10548 266544 10560
rect 266596 10548 266602 10600
rect 64782 10480 64788 10532
rect 64840 10520 64846 10532
rect 255590 10520 255596 10532
rect 64840 10492 255596 10520
rect 64840 10480 64846 10492
rect 255590 10480 255596 10492
rect 255648 10480 255654 10532
rect 60642 10412 60648 10464
rect 60700 10452 60706 10464
rect 254026 10452 254032 10464
rect 60700 10424 254032 10452
rect 60700 10412 60706 10424
rect 254026 10412 254032 10424
rect 254084 10412 254090 10464
rect 56502 10344 56508 10396
rect 56560 10384 56566 10396
rect 252646 10384 252652 10396
rect 56560 10356 252652 10384
rect 56560 10344 56566 10356
rect 252646 10344 252652 10356
rect 252704 10344 252710 10396
rect 53742 10276 53748 10328
rect 53800 10316 53806 10328
rect 251266 10316 251272 10328
rect 53800 10288 251272 10316
rect 53800 10276 53806 10288
rect 251266 10276 251272 10288
rect 251324 10276 251330 10328
rect 117130 10208 117136 10260
rect 117188 10248 117194 10260
rect 277578 10248 277584 10260
rect 117188 10220 277584 10248
rect 117188 10208 117194 10220
rect 277578 10208 277584 10220
rect 277636 10208 277642 10260
rect 119982 10140 119988 10192
rect 120040 10180 120046 10192
rect 278958 10180 278964 10192
rect 120040 10152 278964 10180
rect 120040 10140 120046 10152
rect 278958 10140 278964 10152
rect 279016 10140 279022 10192
rect 124122 10072 124128 10124
rect 124180 10112 124186 10124
rect 280338 10112 280344 10124
rect 124180 10084 280344 10112
rect 124180 10072 124186 10084
rect 280338 10072 280344 10084
rect 280396 10072 280402 10124
rect 143442 10004 143448 10056
rect 143500 10044 143506 10056
rect 288526 10044 288532 10056
rect 143500 10016 288532 10044
rect 143500 10004 143506 10016
rect 288526 10004 288532 10016
rect 288584 10004 288590 10056
rect 147582 9936 147588 9988
rect 147640 9976 147646 9988
rect 289814 9976 289820 9988
rect 147640 9948 289820 9976
rect 147640 9936 147646 9948
rect 289814 9936 289820 9948
rect 289872 9936 289878 9988
rect 151630 9868 151636 9920
rect 151688 9908 151694 9920
rect 291286 9908 291292 9920
rect 151688 9880 291292 9908
rect 151688 9868 151694 9880
rect 291286 9868 291292 9880
rect 291344 9868 291350 9920
rect 154482 9800 154488 9852
rect 154540 9840 154546 9852
rect 292850 9840 292856 9852
rect 154540 9812 292856 9840
rect 154540 9800 154546 9812
rect 292850 9800 292856 9812
rect 292908 9800 292914 9852
rect 158622 9732 158628 9784
rect 158680 9772 158686 9784
rect 294046 9772 294052 9784
rect 158680 9744 294052 9772
rect 158680 9732 158686 9744
rect 294046 9732 294052 9744
rect 294104 9732 294110 9784
rect 306742 9772 306748 9784
rect 306668 9744 306748 9772
rect 306668 9716 306696 9744
rect 306742 9732 306748 9744
rect 306800 9732 306806 9784
rect 161382 9664 161388 9716
rect 161440 9704 161446 9716
rect 295426 9704 295432 9716
rect 161440 9676 295432 9704
rect 161440 9664 161446 9676
rect 295426 9664 295432 9676
rect 295484 9664 295490 9716
rect 306650 9664 306656 9716
rect 306708 9664 306714 9716
rect 341242 9704 341248 9716
rect 341203 9676 341248 9704
rect 341242 9664 341248 9676
rect 341300 9664 341306 9716
rect 358538 9704 358544 9716
rect 358499 9676 358544 9704
rect 358538 9664 358544 9676
rect 358596 9664 358602 9716
rect 366818 9704 366824 9716
rect 366779 9676 366824 9704
rect 366818 9664 366824 9676
rect 366876 9664 366882 9716
rect 421193 9707 421251 9713
rect 421193 9673 421205 9707
rect 421239 9704 421251 9707
rect 421374 9704 421380 9716
rect 421239 9676 421380 9704
rect 421239 9673 421251 9676
rect 421193 9667 421251 9673
rect 421374 9664 421380 9676
rect 421432 9664 421438 9716
rect 470594 9704 470600 9716
rect 470555 9676 470600 9704
rect 470594 9664 470600 9676
rect 470652 9664 470658 9716
rect 203886 9596 203892 9648
rect 203944 9636 203950 9648
rect 313366 9636 313372 9648
rect 203944 9608 313372 9636
rect 203944 9596 203950 9608
rect 313366 9596 313372 9608
rect 313424 9596 313430 9648
rect 200390 9528 200396 9580
rect 200448 9568 200454 9580
rect 311986 9568 311992 9580
rect 200448 9540 311992 9568
rect 200448 9528 200454 9540
rect 311986 9528 311992 9540
rect 312044 9528 312050 9580
rect 196802 9460 196808 9512
rect 196860 9500 196866 9512
rect 310606 9500 310612 9512
rect 196860 9472 310612 9500
rect 196860 9460 196866 9472
rect 310606 9460 310612 9472
rect 310664 9460 310670 9512
rect 193214 9392 193220 9444
rect 193272 9432 193278 9444
rect 309226 9432 309232 9444
rect 193272 9404 309232 9432
rect 193272 9392 193278 9404
rect 309226 9392 309232 9404
rect 309284 9392 309290 9444
rect 139670 9324 139676 9376
rect 139728 9364 139734 9376
rect 287146 9364 287152 9376
rect 139728 9336 287152 9364
rect 139728 9324 139734 9336
rect 287146 9324 287152 9336
rect 287204 9324 287210 9376
rect 136082 9256 136088 9308
rect 136140 9296 136146 9308
rect 285858 9296 285864 9308
rect 136140 9268 285864 9296
rect 136140 9256 136146 9268
rect 285858 9256 285864 9268
rect 285916 9256 285922 9308
rect 49326 9188 49332 9240
rect 49384 9228 49390 9240
rect 249886 9228 249892 9240
rect 49384 9200 249892 9228
rect 49384 9188 49390 9200
rect 249886 9188 249892 9200
rect 249944 9188 249950 9240
rect 253842 9188 253848 9240
rect 253900 9228 253906 9240
rect 334158 9228 334164 9240
rect 253900 9200 334164 9228
rect 253900 9188 253906 9200
rect 334158 9188 334164 9200
rect 334216 9188 334222 9240
rect 44542 9120 44548 9172
rect 44600 9160 44606 9172
rect 247126 9160 247132 9172
rect 44600 9132 247132 9160
rect 44600 9120 44606 9132
rect 247126 9120 247132 9132
rect 247184 9120 247190 9172
rect 250346 9120 250352 9172
rect 250404 9160 250410 9172
rect 332778 9160 332784 9172
rect 250404 9132 332784 9160
rect 250404 9120 250410 9132
rect 332778 9120 332784 9132
rect 332836 9120 332842 9172
rect 27890 9052 27896 9104
rect 27948 9092 27954 9104
rect 233878 9092 233884 9104
rect 27948 9064 233884 9092
rect 27948 9052 27954 9064
rect 233878 9052 233884 9064
rect 233936 9052 233942 9104
rect 243170 9052 243176 9104
rect 243228 9092 243234 9104
rect 330018 9092 330024 9104
rect 243228 9064 330024 9092
rect 243228 9052 243234 9064
rect 330018 9052 330024 9064
rect 330076 9052 330082 9104
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 236178 9024 236184 9036
rect 18380 8996 236184 9024
rect 18380 8984 18386 8996
rect 236178 8984 236184 8996
rect 236236 8984 236242 9036
rect 239582 8984 239588 9036
rect 239640 9024 239646 9036
rect 328638 9024 328644 9036
rect 239640 8996 328644 9024
rect 239640 8984 239646 8996
rect 328638 8984 328644 8996
rect 328696 8984 328702 9036
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 234798 8956 234804 8968
rect 13688 8928 234804 8956
rect 13688 8916 13694 8928
rect 234798 8916 234804 8928
rect 234856 8916 234862 8968
rect 235994 8916 236000 8968
rect 236052 8956 236058 8968
rect 325970 8956 325976 8968
rect 236052 8928 325976 8956
rect 236052 8916 236058 8928
rect 325970 8916 325976 8928
rect 326028 8916 326034 8968
rect 207474 8848 207480 8900
rect 207532 8888 207538 8900
rect 314930 8888 314936 8900
rect 207532 8860 314936 8888
rect 207532 8848 207538 8860
rect 314930 8848 314936 8860
rect 314988 8848 314994 8900
rect 210970 8780 210976 8832
rect 211028 8820 211034 8832
rect 316126 8820 316132 8832
rect 211028 8792 316132 8820
rect 211028 8780 211034 8792
rect 316126 8780 316132 8792
rect 316184 8780 316190 8832
rect 214650 8712 214656 8764
rect 214708 8752 214714 8764
rect 317506 8752 317512 8764
rect 214708 8724 317512 8752
rect 214708 8712 214714 8724
rect 317506 8712 317512 8724
rect 317564 8712 317570 8764
rect 218146 8644 218152 8696
rect 218204 8684 218210 8696
rect 318886 8684 318892 8696
rect 218204 8656 318892 8684
rect 218204 8644 218210 8656
rect 318886 8644 318892 8656
rect 318944 8644 318950 8696
rect 221734 8576 221740 8628
rect 221792 8616 221798 8628
rect 320174 8616 320180 8628
rect 221792 8588 320180 8616
rect 221792 8576 221798 8588
rect 320174 8576 320180 8588
rect 320232 8576 320238 8628
rect 225322 8508 225328 8560
rect 225380 8548 225386 8560
rect 321646 8548 321652 8560
rect 225380 8520 321652 8548
rect 225380 8508 225386 8520
rect 321646 8508 321652 8520
rect 321704 8508 321710 8560
rect 228910 8440 228916 8492
rect 228968 8480 228974 8492
rect 323302 8480 323308 8492
rect 228968 8452 323308 8480
rect 228968 8440 228974 8452
rect 323302 8440 323308 8452
rect 323360 8440 323366 8492
rect 232498 8372 232504 8424
rect 232556 8412 232562 8424
rect 324590 8412 324596 8424
rect 232556 8384 324596 8412
rect 232556 8372 232562 8384
rect 324590 8372 324596 8384
rect 324648 8372 324654 8424
rect 236270 8344 236276 8356
rect 236231 8316 236276 8344
rect 236270 8304 236276 8316
rect 236328 8304 236334 8356
rect 238938 8304 238944 8356
rect 238996 8344 239002 8356
rect 239030 8344 239036 8356
rect 238996 8316 239036 8344
rect 238996 8304 239002 8316
rect 239030 8304 239036 8316
rect 239088 8304 239094 8356
rect 244366 8344 244372 8356
rect 244327 8316 244372 8344
rect 244366 8304 244372 8316
rect 244424 8304 244430 8356
rect 246758 8304 246764 8356
rect 246816 8344 246822 8356
rect 331398 8344 331404 8356
rect 246816 8316 331404 8344
rect 246816 8304 246822 8316
rect 331398 8304 331404 8316
rect 331456 8304 331462 8356
rect 468754 8304 468760 8356
rect 468812 8344 468818 8356
rect 469030 8344 469036 8356
rect 468812 8316 469036 8344
rect 468812 8304 468818 8316
rect 469030 8304 469036 8316
rect 469088 8304 469094 8356
rect 87322 8236 87328 8288
rect 87380 8276 87386 8288
rect 265158 8276 265164 8288
rect 87380 8248 265164 8276
rect 87380 8236 87386 8248
rect 265158 8236 265164 8248
rect 265216 8236 265222 8288
rect 270494 8236 270500 8288
rect 270552 8276 270558 8288
rect 340966 8276 340972 8288
rect 270552 8248 340972 8276
rect 270552 8236 270558 8248
rect 340966 8236 340972 8248
rect 341024 8236 341030 8288
rect 445478 8236 445484 8288
rect 445536 8276 445542 8288
rect 523862 8276 523868 8288
rect 445536 8248 523868 8276
rect 445536 8236 445542 8248
rect 523862 8236 523868 8248
rect 523920 8236 523926 8288
rect 83826 8168 83832 8220
rect 83884 8208 83890 8220
rect 263870 8208 263876 8220
rect 83884 8180 263876 8208
rect 83884 8168 83890 8180
rect 263870 8168 263876 8180
rect 263928 8168 263934 8220
rect 266998 8168 267004 8220
rect 267056 8208 267062 8220
rect 339586 8208 339592 8220
rect 267056 8180 339592 8208
rect 267056 8168 267062 8180
rect 339586 8168 339592 8180
rect 339644 8168 339650 8220
rect 446950 8168 446956 8220
rect 447008 8208 447014 8220
rect 527450 8208 527456 8220
rect 447008 8180 527456 8208
rect 447008 8168 447014 8180
rect 527450 8168 527456 8180
rect 527508 8168 527514 8220
rect 80238 8100 80244 8152
rect 80296 8140 80302 8152
rect 262398 8140 262404 8152
rect 80296 8112 262404 8140
rect 80296 8100 80302 8112
rect 262398 8100 262404 8112
rect 262456 8100 262462 8152
rect 263410 8100 263416 8152
rect 263468 8140 263474 8152
rect 338298 8140 338304 8152
rect 263468 8112 338304 8140
rect 263468 8100 263474 8112
rect 338298 8100 338304 8112
rect 338356 8100 338362 8152
rect 448238 8100 448244 8152
rect 448296 8140 448302 8152
rect 531038 8140 531044 8152
rect 448296 8112 531044 8140
rect 448296 8100 448302 8112
rect 531038 8100 531044 8112
rect 531096 8100 531102 8152
rect 40954 8032 40960 8084
rect 41012 8072 41018 8084
rect 245838 8072 245844 8084
rect 41012 8044 245844 8072
rect 41012 8032 41018 8044
rect 245838 8032 245844 8044
rect 245896 8032 245902 8084
rect 259822 8032 259828 8084
rect 259880 8072 259886 8084
rect 336918 8072 336924 8084
rect 259880 8044 336924 8072
rect 259880 8032 259886 8044
rect 336918 8032 336924 8044
rect 336976 8032 336982 8084
rect 450998 8032 451004 8084
rect 451056 8072 451062 8084
rect 534534 8072 534540 8084
rect 451056 8044 534540 8072
rect 451056 8032 451062 8044
rect 534534 8032 534540 8044
rect 534592 8032 534598 8084
rect 37366 7964 37372 8016
rect 37424 8004 37430 8016
rect 244366 8004 244372 8016
rect 37424 7976 244372 8004
rect 37424 7964 37430 7976
rect 244366 7964 244372 7976
rect 244424 7964 244430 8016
rect 256234 7964 256240 8016
rect 256292 8004 256298 8016
rect 334066 8004 334072 8016
rect 256292 7976 334072 8004
rect 256292 7964 256298 7976
rect 334066 7964 334072 7976
rect 334124 7964 334130 8016
rect 452470 7964 452476 8016
rect 452528 8004 452534 8016
rect 538122 8004 538128 8016
rect 452528 7976 538128 8004
rect 452528 7964 452534 7976
rect 538122 7964 538128 7976
rect 538180 7964 538186 8016
rect 33870 7896 33876 7948
rect 33928 7936 33934 7948
rect 242986 7936 242992 7948
rect 33928 7908 242992 7936
rect 33928 7896 33934 7908
rect 242986 7896 242992 7908
rect 243044 7896 243050 7948
rect 252646 7896 252652 7948
rect 252704 7936 252710 7948
rect 332686 7936 332692 7948
rect 252704 7908 332692 7936
rect 252704 7896 252710 7908
rect 332686 7896 332692 7908
rect 332744 7896 332750 7948
rect 453758 7896 453764 7948
rect 453816 7936 453822 7948
rect 541710 7936 541716 7948
rect 453816 7908 541716 7936
rect 453816 7896 453822 7908
rect 541710 7896 541716 7908
rect 541768 7896 541774 7948
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 241790 7868 241796 7880
rect 30340 7840 241796 7868
rect 30340 7828 30346 7840
rect 241790 7828 241796 7840
rect 241848 7828 241854 7880
rect 249150 7828 249156 7880
rect 249208 7868 249214 7880
rect 331306 7868 331312 7880
rect 249208 7840 331312 7868
rect 249208 7828 249214 7840
rect 331306 7828 331312 7840
rect 331364 7828 331370 7880
rect 455230 7828 455236 7880
rect 455288 7868 455294 7880
rect 545298 7868 545304 7880
rect 455288 7840 545304 7868
rect 455288 7828 455294 7840
rect 545298 7828 545304 7840
rect 545356 7828 545362 7880
rect 26694 7760 26700 7812
rect 26752 7800 26758 7812
rect 240410 7800 240416 7812
rect 26752 7772 240416 7800
rect 26752 7760 26758 7772
rect 240410 7760 240416 7772
rect 240468 7760 240474 7812
rect 245562 7760 245568 7812
rect 245620 7800 245626 7812
rect 330202 7800 330208 7812
rect 245620 7772 330208 7800
rect 245620 7760 245626 7772
rect 330202 7760 330208 7772
rect 330260 7760 330266 7812
rect 456610 7760 456616 7812
rect 456668 7800 456674 7812
rect 548886 7800 548892 7812
rect 456668 7772 548892 7800
rect 456668 7760 456674 7772
rect 548886 7760 548892 7772
rect 548944 7760 548950 7812
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 238846 7732 238852 7744
rect 21968 7704 238852 7732
rect 21968 7692 21974 7704
rect 238846 7692 238852 7704
rect 238904 7692 238910 7744
rect 241974 7692 241980 7744
rect 242032 7732 242038 7744
rect 328546 7732 328552 7744
rect 242032 7704 328552 7732
rect 242032 7692 242038 7704
rect 328546 7692 328552 7704
rect 328604 7692 328610 7744
rect 457990 7692 457996 7744
rect 458048 7732 458054 7744
rect 552382 7732 552388 7744
rect 458048 7704 552388 7732
rect 458048 7692 458054 7704
rect 552382 7692 552388 7704
rect 552440 7692 552446 7744
rect 8846 7624 8852 7676
rect 8904 7664 8910 7676
rect 227533 7667 227591 7673
rect 227533 7664 227545 7667
rect 8904 7636 227545 7664
rect 8904 7624 8910 7636
rect 227533 7633 227545 7636
rect 227579 7633 227591 7667
rect 230658 7664 230664 7676
rect 227533 7627 227591 7633
rect 227640 7636 230664 7664
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 227640 7596 227668 7636
rect 230658 7624 230664 7636
rect 230716 7624 230722 7676
rect 234798 7624 234804 7676
rect 234856 7664 234862 7676
rect 325786 7664 325792 7676
rect 234856 7636 325792 7664
rect 234856 7624 234862 7636
rect 325786 7624 325792 7636
rect 325844 7624 325850 7676
rect 459370 7624 459376 7676
rect 459428 7664 459434 7676
rect 555970 7664 555976 7676
rect 459428 7636 555976 7664
rect 459428 7624 459434 7636
rect 555970 7624 555976 7636
rect 556028 7624 556034 7676
rect 4120 7568 227668 7596
rect 4120 7556 4126 7568
rect 227714 7556 227720 7608
rect 227772 7596 227778 7608
rect 229002 7596 229008 7608
rect 227772 7568 229008 7596
rect 227772 7556 227778 7568
rect 229002 7556 229008 7568
rect 229060 7556 229066 7608
rect 231302 7556 231308 7608
rect 231360 7596 231366 7608
rect 324406 7596 324412 7608
rect 231360 7568 324412 7596
rect 231360 7556 231366 7568
rect 324406 7556 324412 7568
rect 324464 7556 324470 7608
rect 460750 7556 460756 7608
rect 460808 7596 460814 7608
rect 559558 7596 559564 7608
rect 460808 7568 559564 7596
rect 460808 7556 460814 7568
rect 559558 7556 559564 7568
rect 559616 7556 559622 7608
rect 134886 7488 134892 7540
rect 134944 7528 134950 7540
rect 284570 7528 284576 7540
rect 134944 7500 284576 7528
rect 134944 7488 134950 7500
rect 284570 7488 284576 7500
rect 284628 7488 284634 7540
rect 444190 7488 444196 7540
rect 444248 7528 444254 7540
rect 520274 7528 520280 7540
rect 444248 7500 520280 7528
rect 444248 7488 444254 7500
rect 520274 7488 520280 7500
rect 520332 7488 520338 7540
rect 138474 7420 138480 7472
rect 138532 7460 138538 7472
rect 285950 7460 285956 7472
rect 138532 7432 285956 7460
rect 138532 7420 138538 7432
rect 285950 7420 285956 7432
rect 286008 7420 286014 7472
rect 442810 7420 442816 7472
rect 442868 7460 442874 7472
rect 516778 7460 516784 7472
rect 442868 7432 516784 7460
rect 442868 7420 442874 7432
rect 516778 7420 516784 7432
rect 516836 7420 516842 7472
rect 141970 7352 141976 7404
rect 142028 7392 142034 7404
rect 287054 7392 287060 7404
rect 142028 7364 287060 7392
rect 142028 7352 142034 7364
rect 287054 7352 287060 7364
rect 287112 7352 287118 7404
rect 441430 7352 441436 7404
rect 441488 7392 441494 7404
rect 513190 7392 513196 7404
rect 441488 7364 513196 7392
rect 441488 7352 441494 7364
rect 513190 7352 513196 7364
rect 513248 7352 513254 7404
rect 145650 7284 145656 7336
rect 145708 7324 145714 7336
rect 288434 7324 288440 7336
rect 145708 7296 288440 7324
rect 145708 7284 145714 7296
rect 288434 7284 288440 7296
rect 288492 7284 288498 7336
rect 440050 7284 440056 7336
rect 440108 7324 440114 7336
rect 509602 7324 509608 7336
rect 440108 7296 509608 7324
rect 440108 7284 440114 7296
rect 509602 7284 509608 7296
rect 509660 7284 509666 7336
rect 149238 7216 149244 7268
rect 149296 7256 149302 7268
rect 291194 7256 291200 7268
rect 149296 7228 291200 7256
rect 149296 7216 149302 7228
rect 291194 7216 291200 7228
rect 291252 7216 291258 7268
rect 152734 7148 152740 7200
rect 152792 7188 152798 7200
rect 292574 7188 292580 7200
rect 152792 7160 292580 7188
rect 152792 7148 152798 7160
rect 292574 7148 292580 7160
rect 292632 7148 292638 7200
rect 156322 7080 156328 7132
rect 156380 7120 156386 7132
rect 293954 7120 293960 7132
rect 156380 7092 293960 7120
rect 156380 7080 156386 7092
rect 293954 7080 293960 7092
rect 294012 7080 294018 7132
rect 159910 7012 159916 7064
rect 159968 7052 159974 7064
rect 295334 7052 295340 7064
rect 159968 7024 295340 7052
rect 159968 7012 159974 7024
rect 295334 7012 295340 7024
rect 295392 7012 295398 7064
rect 227533 6987 227591 6993
rect 227533 6953 227545 6987
rect 227579 6984 227591 6987
rect 233418 6984 233424 6996
rect 227579 6956 233424 6984
rect 227579 6953 227591 6956
rect 227533 6947 227591 6953
rect 233418 6944 233424 6956
rect 233476 6944 233482 6996
rect 238386 6944 238392 6996
rect 238444 6984 238450 6996
rect 327258 6984 327264 6996
rect 238444 6956 327264 6984
rect 238444 6944 238450 6956
rect 327258 6944 327264 6956
rect 327316 6944 327322 6996
rect 516686 6876 516692 6928
rect 516744 6916 516750 6928
rect 516870 6916 516876 6928
rect 516744 6888 516876 6916
rect 516744 6876 516750 6888
rect 516870 6876 516876 6888
rect 516928 6876 516934 6928
rect 170582 6808 170588 6860
rect 170640 6848 170646 6860
rect 299474 6848 299480 6860
rect 170640 6820 299480 6848
rect 170640 6808 170646 6820
rect 299474 6808 299480 6820
rect 299532 6808 299538 6860
rect 431770 6808 431776 6860
rect 431828 6848 431834 6860
rect 490558 6848 490564 6860
rect 431828 6820 490564 6848
rect 431828 6808 431834 6820
rect 490558 6808 490564 6820
rect 490616 6808 490622 6860
rect 167086 6740 167092 6792
rect 167144 6780 167150 6792
rect 298370 6780 298376 6792
rect 167144 6752 298376 6780
rect 167144 6740 167150 6752
rect 298370 6740 298376 6752
rect 298428 6740 298434 6792
rect 433150 6740 433156 6792
rect 433208 6780 433214 6792
rect 491754 6780 491760 6792
rect 433208 6752 491760 6780
rect 433208 6740 433214 6752
rect 491754 6740 491760 6752
rect 491812 6740 491818 6792
rect 163498 6672 163504 6724
rect 163556 6712 163562 6724
rect 296714 6712 296720 6724
rect 163556 6684 296720 6712
rect 163556 6672 163562 6684
rect 296714 6672 296720 6684
rect 296772 6672 296778 6724
rect 298094 6672 298100 6724
rect 298152 6712 298158 6724
rect 338390 6712 338396 6724
rect 298152 6684 338396 6712
rect 298152 6672 298158 6684
rect 338390 6672 338396 6684
rect 338448 6672 338454 6724
rect 434622 6672 434628 6724
rect 434680 6712 434686 6724
rect 495342 6712 495348 6724
rect 434680 6684 495348 6712
rect 434680 6672 434686 6684
rect 495342 6672 495348 6684
rect 495400 6672 495406 6724
rect 131390 6604 131396 6656
rect 131448 6644 131454 6656
rect 283006 6644 283012 6656
rect 131448 6616 283012 6644
rect 131448 6604 131454 6616
rect 283006 6604 283012 6616
rect 283064 6604 283070 6656
rect 297358 6604 297364 6656
rect 297416 6644 297422 6656
rect 336826 6644 336832 6656
rect 297416 6616 336832 6644
rect 297416 6604 297422 6616
rect 336826 6604 336832 6616
rect 336884 6604 336890 6656
rect 436002 6604 436008 6656
rect 436060 6644 436066 6656
rect 497734 6644 497740 6656
rect 436060 6616 497740 6644
rect 436060 6604 436066 6616
rect 497734 6604 497740 6616
rect 497792 6604 497798 6656
rect 76650 6536 76656 6588
rect 76708 6576 76714 6588
rect 261018 6576 261024 6588
rect 76708 6548 261024 6576
rect 76708 6536 76714 6548
rect 261018 6536 261024 6548
rect 261076 6536 261082 6588
rect 295886 6536 295892 6588
rect 295944 6576 295950 6588
rect 335446 6576 335452 6588
rect 295944 6548 335452 6576
rect 295944 6536 295950 6548
rect 335446 6536 335452 6548
rect 335504 6536 335510 6588
rect 433242 6536 433248 6588
rect 433300 6576 433306 6588
rect 494146 6576 494152 6588
rect 433300 6548 494152 6576
rect 433300 6536 433306 6548
rect 494146 6536 494152 6548
rect 494204 6536 494210 6588
rect 73062 6468 73068 6520
rect 73120 6508 73126 6520
rect 259454 6508 259460 6520
rect 73120 6480 259460 6508
rect 73120 6468 73126 6480
rect 259454 6468 259460 6480
rect 259512 6468 259518 6520
rect 289814 6468 289820 6520
rect 289872 6508 289878 6520
rect 339678 6508 339684 6520
rect 289872 6480 339684 6508
rect 289872 6468 289878 6480
rect 339678 6468 339684 6480
rect 339736 6468 339742 6520
rect 433518 6468 433524 6520
rect 433576 6508 433582 6520
rect 434622 6508 434628 6520
rect 433576 6480 434628 6508
rect 433576 6468 433582 6480
rect 434622 6468 434628 6480
rect 434680 6468 434686 6520
rect 435910 6468 435916 6520
rect 435968 6508 435974 6520
rect 498930 6508 498936 6520
rect 435968 6480 498936 6508
rect 435968 6468 435974 6480
rect 498930 6468 498936 6480
rect 498988 6468 498994 6520
rect 69474 6400 69480 6452
rect 69532 6440 69538 6452
rect 258258 6440 258264 6452
rect 69532 6412 258264 6440
rect 69532 6400 69538 6412
rect 258258 6400 258264 6412
rect 258316 6400 258322 6452
rect 288434 6400 288440 6452
rect 288492 6440 288498 6452
rect 341242 6440 341248 6452
rect 288492 6412 341248 6440
rect 288492 6400 288498 6412
rect 341242 6400 341248 6412
rect 341300 6400 341306 6452
rect 437290 6400 437296 6452
rect 437348 6440 437354 6452
rect 501230 6440 501236 6452
rect 437348 6412 501236 6440
rect 437348 6400 437354 6412
rect 501230 6400 501236 6412
rect 501288 6400 501294 6452
rect 65978 6332 65984 6384
rect 66036 6372 66042 6384
rect 256786 6372 256792 6384
rect 66036 6344 256792 6372
rect 66036 6332 66042 6344
rect 256786 6332 256792 6344
rect 256844 6332 256850 6384
rect 288526 6332 288532 6384
rect 288584 6372 288590 6384
rect 343634 6372 343640 6384
rect 288584 6344 343640 6372
rect 288584 6332 288590 6344
rect 343634 6332 343640 6344
rect 343692 6332 343698 6384
rect 437382 6332 437388 6384
rect 437440 6372 437446 6384
rect 502426 6372 502432 6384
rect 437440 6344 502432 6372
rect 437440 6332 437446 6344
rect 502426 6332 502432 6344
rect 502484 6332 502490 6384
rect 62390 6264 62396 6316
rect 62448 6304 62454 6316
rect 255498 6304 255504 6316
rect 62448 6276 255504 6304
rect 62448 6264 62454 6276
rect 255498 6264 255504 6276
rect 255556 6264 255562 6316
rect 294322 6264 294328 6316
rect 294380 6304 294386 6316
rect 350626 6304 350632 6316
rect 294380 6276 350632 6304
rect 294380 6264 294386 6276
rect 350626 6264 350632 6276
rect 350684 6264 350690 6316
rect 438670 6264 438676 6316
rect 438728 6304 438734 6316
rect 504818 6304 504824 6316
rect 438728 6276 504824 6304
rect 438728 6264 438734 6276
rect 504818 6264 504824 6276
rect 504876 6264 504882 6316
rect 58802 6196 58808 6248
rect 58860 6236 58866 6248
rect 253934 6236 253940 6248
rect 58860 6208 253940 6236
rect 58860 6196 58866 6208
rect 253934 6196 253940 6208
rect 253992 6196 253998 6248
rect 280062 6196 280068 6248
rect 280120 6236 280126 6248
rect 345198 6236 345204 6248
rect 280120 6208 345204 6236
rect 280120 6196 280126 6208
rect 345198 6196 345204 6208
rect 345256 6196 345262 6248
rect 438762 6196 438768 6248
rect 438820 6236 438826 6248
rect 506014 6236 506020 6248
rect 438820 6208 506020 6236
rect 438820 6196 438826 6208
rect 506014 6196 506020 6208
rect 506072 6196 506078 6248
rect 55214 6128 55220 6180
rect 55272 6168 55278 6180
rect 251358 6168 251364 6180
rect 55272 6140 251364 6168
rect 55272 6128 55278 6140
rect 251358 6128 251364 6140
rect 251416 6128 251422 6180
rect 274082 6128 274088 6180
rect 274140 6168 274146 6180
rect 342346 6168 342352 6180
rect 274140 6140 342352 6168
rect 274140 6128 274146 6140
rect 342346 6128 342352 6140
rect 342404 6128 342410 6180
rect 440142 6128 440148 6180
rect 440200 6168 440206 6180
rect 508406 6168 508412 6180
rect 440200 6140 508412 6168
rect 440200 6128 440206 6140
rect 508406 6128 508412 6140
rect 508464 6128 508470 6180
rect 174170 6060 174176 6112
rect 174228 6100 174234 6112
rect 300854 6100 300860 6112
rect 174228 6072 300860 6100
rect 174228 6060 174234 6072
rect 300854 6060 300860 6072
rect 300912 6060 300918 6112
rect 337102 6100 337108 6112
rect 337063 6072 337108 6100
rect 337102 6060 337108 6072
rect 337160 6060 337166 6112
rect 430390 6060 430396 6112
rect 430448 6100 430454 6112
rect 486970 6100 486976 6112
rect 430448 6072 486976 6100
rect 430448 6060 430454 6072
rect 486970 6060 486976 6072
rect 487028 6060 487034 6112
rect 177758 5992 177764 6044
rect 177816 6032 177822 6044
rect 302234 6032 302240 6044
rect 177816 6004 302240 6032
rect 177816 5992 177822 6004
rect 302234 5992 302240 6004
rect 302292 5992 302298 6044
rect 431862 5992 431868 6044
rect 431920 6032 431926 6044
rect 488166 6032 488172 6044
rect 431920 6004 488172 6032
rect 431920 5992 431926 6004
rect 488166 5992 488172 6004
rect 488224 5992 488230 6044
rect 181346 5924 181352 5976
rect 181404 5964 181410 5976
rect 303614 5964 303620 5976
rect 181404 5936 303620 5964
rect 181404 5924 181410 5936
rect 303614 5924 303620 5936
rect 303672 5924 303678 5976
rect 429102 5924 429108 5976
rect 429160 5964 429166 5976
rect 483474 5964 483480 5976
rect 429160 5936 483480 5964
rect 429160 5924 429166 5936
rect 483474 5924 483480 5936
rect 483532 5924 483538 5976
rect 184842 5856 184848 5908
rect 184900 5896 184906 5908
rect 304994 5896 305000 5908
rect 184900 5868 305000 5896
rect 184900 5856 184906 5868
rect 304994 5856 305000 5868
rect 305052 5856 305058 5908
rect 430482 5856 430488 5908
rect 430540 5896 430546 5908
rect 484578 5896 484584 5908
rect 430540 5868 484584 5896
rect 430540 5856 430546 5868
rect 484578 5856 484584 5868
rect 484636 5856 484642 5908
rect 188430 5788 188436 5840
rect 188488 5828 188494 5840
rect 306650 5828 306656 5840
rect 188488 5800 306656 5828
rect 188488 5788 188494 5800
rect 306650 5788 306656 5800
rect 306708 5788 306714 5840
rect 427722 5788 427728 5840
rect 427780 5828 427786 5840
rect 479886 5828 479892 5840
rect 427780 5800 479892 5828
rect 427780 5788 427786 5800
rect 479886 5788 479892 5800
rect 479944 5788 479950 5840
rect 192018 5720 192024 5772
rect 192076 5760 192082 5772
rect 307754 5760 307760 5772
rect 192076 5732 307760 5760
rect 192076 5720 192082 5732
rect 307754 5720 307760 5732
rect 307812 5720 307818 5772
rect 426342 5720 426348 5772
rect 426400 5760 426406 5772
rect 476298 5760 476304 5772
rect 426400 5732 476304 5760
rect 426400 5720 426406 5732
rect 476298 5720 476304 5732
rect 476356 5720 476362 5772
rect 195606 5652 195612 5704
rect 195664 5692 195670 5704
rect 309134 5692 309140 5704
rect 195664 5664 309140 5692
rect 195664 5652 195670 5664
rect 309134 5652 309140 5664
rect 309192 5652 309198 5704
rect 199194 5584 199200 5636
rect 199252 5624 199258 5636
rect 310514 5624 310520 5636
rect 199252 5596 310520 5624
rect 199252 5584 199258 5596
rect 310514 5584 310520 5596
rect 310572 5584 310578 5636
rect 470594 5584 470600 5636
rect 470652 5624 470658 5636
rect 471517 5627 471575 5633
rect 471517 5624 471529 5627
rect 470652 5596 471529 5624
rect 470652 5584 470658 5596
rect 471517 5593 471529 5596
rect 471563 5593 471575 5627
rect 471517 5587 471575 5593
rect 202690 5516 202696 5568
rect 202748 5556 202754 5568
rect 313274 5556 313280 5568
rect 202748 5528 313280 5556
rect 202748 5516 202754 5528
rect 313274 5516 313280 5528
rect 313332 5516 313338 5568
rect 468938 5516 468944 5568
rect 468996 5556 469002 5568
rect 471425 5559 471483 5565
rect 471425 5556 471437 5559
rect 468996 5528 471437 5556
rect 468996 5516 469002 5528
rect 471425 5525 471437 5528
rect 471471 5525 471483 5559
rect 471425 5519 471483 5525
rect 137278 5448 137284 5500
rect 137336 5488 137342 5500
rect 285674 5488 285680 5500
rect 137336 5460 285680 5488
rect 137336 5448 137342 5460
rect 285674 5448 285680 5460
rect 285732 5448 285738 5500
rect 287701 5491 287759 5497
rect 287701 5457 287713 5491
rect 287747 5488 287759 5491
rect 297085 5491 297143 5497
rect 297085 5488 297097 5491
rect 287747 5460 297097 5488
rect 287747 5457 287759 5460
rect 287701 5451 287759 5457
rect 297085 5457 297097 5460
rect 297131 5457 297143 5491
rect 297085 5451 297143 5457
rect 297818 5448 297824 5500
rect 297876 5488 297882 5500
rect 352098 5488 352104 5500
rect 297876 5460 352104 5488
rect 297876 5448 297882 5460
rect 352098 5448 352104 5460
rect 352156 5448 352162 5500
rect 452562 5448 452568 5500
rect 452620 5488 452626 5500
rect 540514 5488 540520 5500
rect 452620 5460 540520 5488
rect 452620 5448 452626 5460
rect 540514 5448 540520 5460
rect 540572 5448 540578 5500
rect 133782 5380 133788 5432
rect 133840 5420 133846 5432
rect 284294 5420 284300 5432
rect 133840 5392 284300 5420
rect 133840 5380 133846 5392
rect 284294 5380 284300 5392
rect 284352 5380 284358 5432
rect 290734 5380 290740 5432
rect 290792 5420 290798 5432
rect 349338 5420 349344 5432
rect 290792 5392 349344 5420
rect 290792 5380 290798 5392
rect 349338 5380 349344 5392
rect 349396 5380 349402 5432
rect 408402 5380 408408 5432
rect 408460 5420 408466 5432
rect 433518 5420 433524 5432
rect 408460 5392 433524 5420
rect 408460 5380 408466 5392
rect 433518 5380 433524 5392
rect 433576 5380 433582 5432
rect 453850 5380 453856 5432
rect 453908 5420 453914 5432
rect 544102 5420 544108 5432
rect 453908 5392 544108 5420
rect 453908 5380 453914 5392
rect 544102 5380 544108 5392
rect 544160 5380 544166 5432
rect 130194 5312 130200 5364
rect 130252 5352 130258 5364
rect 283190 5352 283196 5364
rect 130252 5324 283196 5352
rect 130252 5312 130258 5324
rect 283190 5312 283196 5324
rect 283248 5312 283254 5364
rect 287146 5312 287152 5364
rect 287204 5352 287210 5364
rect 347958 5352 347964 5364
rect 287204 5324 347964 5352
rect 287204 5312 287210 5324
rect 347958 5312 347964 5324
rect 348016 5312 348022 5364
rect 412358 5312 412364 5364
rect 412416 5352 412422 5364
rect 440602 5352 440608 5364
rect 412416 5324 440608 5352
rect 412416 5312 412422 5324
rect 440602 5312 440608 5324
rect 440660 5312 440666 5364
rect 455322 5312 455328 5364
rect 455380 5352 455386 5364
rect 547690 5352 547696 5364
rect 455380 5324 547696 5352
rect 455380 5312 455386 5324
rect 547690 5312 547696 5324
rect 547748 5312 547754 5364
rect 67174 5244 67180 5296
rect 67232 5284 67238 5296
rect 256970 5284 256976 5296
rect 67232 5256 256976 5284
rect 67232 5244 67238 5256
rect 256970 5244 256976 5256
rect 257028 5244 257034 5296
rect 268381 5287 268439 5293
rect 268381 5253 268393 5287
rect 268427 5284 268439 5287
rect 278041 5287 278099 5293
rect 278041 5284 278053 5287
rect 268427 5256 278053 5284
rect 268427 5253 268439 5256
rect 268381 5247 268439 5253
rect 278041 5253 278053 5256
rect 278087 5253 278099 5287
rect 278041 5247 278099 5253
rect 283650 5244 283656 5296
rect 283708 5284 283714 5296
rect 346578 5284 346584 5296
rect 283708 5256 346584 5284
rect 283708 5244 283714 5256
rect 346578 5244 346584 5256
rect 346636 5244 346642 5296
rect 413830 5244 413836 5296
rect 413888 5284 413894 5296
rect 444190 5284 444196 5296
rect 413888 5256 444196 5284
rect 413888 5244 413894 5256
rect 444190 5244 444196 5256
rect 444248 5244 444254 5296
rect 459462 5244 459468 5296
rect 459520 5284 459526 5296
rect 466089 5287 466147 5293
rect 459520 5256 466040 5284
rect 459520 5244 459526 5256
rect 48130 5176 48136 5228
rect 48188 5216 48194 5228
rect 248506 5216 248512 5228
rect 48188 5188 248512 5216
rect 48188 5176 48194 5188
rect 248506 5176 248512 5188
rect 248564 5176 248570 5228
rect 251450 5176 251456 5228
rect 251508 5216 251514 5228
rect 332594 5216 332600 5228
rect 251508 5188 332600 5216
rect 251508 5176 251514 5188
rect 332594 5176 332600 5188
rect 332652 5176 332658 5228
rect 415302 5176 415308 5228
rect 415360 5216 415366 5228
rect 447778 5216 447784 5228
rect 415360 5188 447784 5216
rect 415360 5176 415366 5188
rect 447778 5176 447784 5188
rect 447836 5176 447842 5228
rect 460842 5176 460848 5228
rect 460900 5216 460906 5228
rect 466012 5216 466040 5256
rect 466089 5253 466101 5287
rect 466135 5284 466147 5287
rect 551186 5284 551192 5296
rect 466135 5256 551192 5284
rect 466135 5253 466147 5256
rect 466089 5247 466147 5253
rect 551186 5244 551192 5256
rect 551244 5244 551250 5296
rect 554774 5216 554780 5228
rect 460900 5188 465948 5216
rect 466012 5188 554780 5216
rect 460900 5176 460906 5188
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 236086 5148 236092 5160
rect 17276 5120 236092 5148
rect 17276 5108 17282 5120
rect 236086 5108 236092 5120
rect 236144 5108 236150 5160
rect 247954 5108 247960 5160
rect 248012 5148 248018 5160
rect 331214 5148 331220 5160
rect 248012 5120 331220 5148
rect 248012 5108 248018 5120
rect 331214 5108 331220 5120
rect 331272 5108 331278 5160
rect 416498 5108 416504 5160
rect 416556 5148 416562 5160
rect 451274 5148 451280 5160
rect 416556 5120 451280 5148
rect 416556 5108 416562 5120
rect 451274 5108 451280 5120
rect 451332 5108 451338 5160
rect 461213 5151 461271 5157
rect 461213 5117 461225 5151
rect 461259 5148 461271 5151
rect 461259 5120 462268 5148
rect 461259 5117 461271 5120
rect 461213 5111 461271 5117
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 234706 5080 234712 5092
rect 12492 5052 234712 5080
rect 12492 5040 12498 5052
rect 234706 5040 234712 5052
rect 234764 5040 234770 5092
rect 244366 5040 244372 5092
rect 244424 5080 244430 5092
rect 322661 5083 322719 5089
rect 322661 5080 322673 5083
rect 244424 5052 322673 5080
rect 244424 5040 244430 5052
rect 322661 5049 322673 5052
rect 322707 5049 322719 5083
rect 322661 5043 322719 5049
rect 322753 5083 322811 5089
rect 322753 5049 322765 5083
rect 322799 5080 322811 5083
rect 327074 5080 327080 5092
rect 322799 5052 327080 5080
rect 322799 5049 322811 5052
rect 322753 5043 322811 5049
rect 327074 5040 327080 5052
rect 327132 5040 327138 5092
rect 327169 5083 327227 5089
rect 327169 5049 327181 5083
rect 327215 5080 327227 5083
rect 329834 5080 329840 5092
rect 327215 5052 329840 5080
rect 327215 5049 327227 5052
rect 327169 5043 327227 5049
rect 329834 5040 329840 5052
rect 329892 5040 329898 5092
rect 337102 5040 337108 5092
rect 337160 5080 337166 5092
rect 368566 5080 368572 5092
rect 337160 5052 368572 5080
rect 337160 5040 337166 5052
rect 368566 5040 368572 5052
rect 368624 5040 368630 5092
rect 417970 5040 417976 5092
rect 418028 5080 418034 5092
rect 454862 5080 454868 5092
rect 418028 5052 454868 5080
rect 418028 5040 418034 5052
rect 454862 5040 454868 5052
rect 454920 5040 454926 5092
rect 458082 5040 458088 5092
rect 458140 5080 458146 5092
rect 458140 5052 462176 5080
rect 458140 5040 458146 5052
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 232130 5012 232136 5024
rect 7708 4984 232136 5012
rect 7708 4972 7714 4984
rect 232130 4972 232136 4984
rect 232188 4972 232194 5024
rect 240778 4972 240784 5024
rect 240836 5012 240842 5024
rect 249061 5015 249119 5021
rect 249061 5012 249073 5015
rect 240836 4984 249073 5012
rect 240836 4972 240842 4984
rect 249061 4981 249073 4984
rect 249107 4981 249119 5015
rect 249061 4975 249119 4981
rect 257985 5015 258043 5021
rect 257985 4981 257997 5015
rect 258031 5012 258043 5015
rect 268381 5015 268439 5021
rect 268381 5012 268393 5015
rect 258031 4984 268393 5012
rect 258031 4981 258043 4984
rect 257985 4975 258043 4981
rect 268381 4981 268393 4984
rect 268427 4981 268439 5015
rect 268381 4975 268439 4981
rect 278041 5015 278099 5021
rect 278041 4981 278053 5015
rect 278087 5012 278099 5015
rect 287701 5015 287759 5021
rect 287701 5012 287713 5015
rect 278087 4984 287713 5012
rect 278087 4981 278099 4984
rect 278041 4975 278099 4981
rect 287701 4981 287713 4984
rect 287747 4981 287759 5015
rect 287701 4975 287759 4981
rect 297085 5015 297143 5021
rect 297085 4981 297097 5015
rect 297131 5012 297143 5015
rect 307021 5015 307079 5021
rect 307021 5012 307033 5015
rect 297131 4984 307033 5012
rect 297131 4981 297143 4984
rect 297085 4975 297143 4981
rect 307021 4981 307033 4984
rect 307067 4981 307079 5015
rect 307021 4975 307079 4981
rect 315942 4972 315948 5024
rect 316000 5012 316006 5024
rect 325145 5015 325203 5021
rect 325145 5012 325157 5015
rect 316000 4984 325157 5012
rect 316000 4972 316006 4984
rect 325145 4981 325157 4984
rect 325191 4981 325203 5015
rect 325145 4975 325203 4981
rect 325602 4972 325608 5024
rect 325660 5012 325666 5024
rect 338114 5012 338120 5024
rect 325660 4984 338120 5012
rect 325660 4972 325666 4984
rect 338114 4972 338120 4984
rect 338172 4972 338178 5024
rect 419442 4972 419448 5024
rect 419500 5012 419506 5024
rect 458450 5012 458456 5024
rect 419500 4984 458456 5012
rect 419500 4972 419506 4984
rect 458450 4972 458456 4984
rect 458508 4972 458514 5024
rect 462038 5012 462044 5024
rect 459388 4984 462044 5012
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 224221 4947 224279 4953
rect 224221 4944 224233 4947
rect 2924 4916 224233 4944
rect 2924 4904 2930 4916
rect 224221 4913 224233 4916
rect 224267 4913 224279 4947
rect 229094 4944 229100 4956
rect 224221 4907 224279 4913
rect 224328 4916 229100 4944
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 224328 4876 224356 4916
rect 229094 4904 229100 4916
rect 229152 4904 229158 4956
rect 237190 4904 237196 4956
rect 237248 4944 237254 4956
rect 237248 4916 317460 4944
rect 237248 4904 237254 4916
rect 624 4848 224356 4876
rect 624 4836 630 4848
rect 230106 4836 230112 4888
rect 230164 4876 230170 4888
rect 317325 4879 317383 4885
rect 317325 4876 317337 4879
rect 230164 4848 317337 4876
rect 230164 4836 230170 4848
rect 317325 4845 317337 4848
rect 317371 4845 317383 4879
rect 317432 4876 317460 4916
rect 318702 4904 318708 4956
rect 318760 4944 318766 4956
rect 326157 4947 326215 4953
rect 326157 4944 326169 4947
rect 318760 4916 326169 4944
rect 318760 4904 318766 4916
rect 326157 4913 326169 4916
rect 326203 4913 326215 4947
rect 328730 4944 328736 4956
rect 326157 4907 326215 4913
rect 326264 4916 328736 4944
rect 322753 4879 322811 4885
rect 322753 4876 322765 4879
rect 317432 4848 322765 4876
rect 317325 4839 317383 4845
rect 322753 4845 322765 4848
rect 322799 4845 322811 4879
rect 325694 4876 325700 4888
rect 322753 4839 322811 4845
rect 322860 4848 325700 4876
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 224129 4811 224187 4817
rect 224129 4808 224141 4811
rect 1728 4780 224141 4808
rect 1728 4768 1734 4780
rect 224129 4777 224141 4780
rect 224175 4777 224187 4811
rect 224129 4771 224187 4777
rect 224221 4811 224279 4817
rect 224221 4777 224233 4811
rect 224267 4808 224279 4811
rect 230750 4808 230756 4820
rect 224267 4780 230756 4808
rect 224267 4777 224279 4780
rect 224221 4771 224279 4777
rect 230750 4768 230756 4780
rect 230808 4768 230814 4820
rect 233694 4768 233700 4820
rect 233752 4808 233758 4820
rect 322860 4808 322888 4848
rect 325694 4836 325700 4848
rect 325752 4836 325758 4888
rect 324314 4808 324320 4820
rect 233752 4780 322888 4808
rect 322952 4780 324320 4808
rect 233752 4768 233758 4780
rect 212258 4700 212264 4752
rect 212316 4740 212322 4752
rect 316034 4740 316040 4752
rect 212316 4712 316040 4740
rect 212316 4700 212322 4712
rect 316034 4700 316040 4712
rect 316092 4700 316098 4752
rect 317325 4743 317383 4749
rect 317325 4709 317337 4743
rect 317371 4740 317383 4743
rect 322952 4740 322980 4780
rect 324314 4768 324320 4780
rect 324372 4768 324378 4820
rect 325145 4811 325203 4817
rect 325145 4777 325157 4811
rect 325191 4808 325203 4811
rect 326264 4808 326292 4916
rect 328730 4904 328736 4916
rect 328788 4904 328794 4956
rect 333606 4904 333612 4956
rect 333664 4944 333670 4956
rect 367186 4944 367192 4956
rect 333664 4916 367192 4944
rect 333664 4904 333670 4916
rect 367186 4904 367192 4916
rect 367244 4904 367250 4956
rect 420730 4904 420736 4956
rect 420788 4944 420794 4956
rect 459388 4944 459416 4984
rect 462038 4972 462044 4984
rect 462096 4972 462102 5024
rect 420788 4916 459416 4944
rect 462148 4944 462176 5052
rect 462240 5012 462268 5120
rect 463510 5108 463516 5160
rect 463568 5148 463574 5160
rect 465920 5148 465948 5188
rect 554774 5176 554780 5188
rect 554832 5176 554838 5228
rect 558362 5148 558368 5160
rect 463568 5120 465856 5148
rect 465920 5120 558368 5148
rect 463568 5108 463574 5120
rect 464982 5040 464988 5092
rect 465040 5080 465046 5092
rect 465828 5080 465856 5120
rect 558362 5108 558368 5120
rect 558420 5108 558426 5160
rect 471333 5083 471391 5089
rect 465040 5052 465764 5080
rect 465828 5052 471284 5080
rect 465040 5040 465046 5052
rect 465626 5012 465632 5024
rect 462240 4984 465632 5012
rect 465626 4972 465632 4984
rect 465684 4972 465690 5024
rect 465736 5012 465764 5052
rect 471256 5012 471284 5052
rect 471333 5049 471345 5083
rect 471379 5080 471391 5083
rect 561950 5080 561956 5092
rect 471379 5052 561956 5080
rect 471379 5049 471391 5052
rect 471333 5043 471391 5049
rect 561950 5040 561956 5052
rect 562008 5040 562014 5092
rect 565538 5012 565544 5024
rect 465736 4984 471192 5012
rect 471256 4984 565544 5012
rect 466089 4947 466147 4953
rect 466089 4944 466101 4947
rect 462148 4916 466101 4944
rect 420788 4904 420794 4916
rect 466089 4913 466101 4916
rect 466135 4913 466147 4947
rect 466089 4907 466147 4913
rect 466178 4904 466184 4956
rect 466236 4944 466242 4956
rect 471164 4944 471192 4984
rect 565538 4972 565544 4984
rect 565596 4972 565602 5024
rect 569034 4944 569040 4956
rect 466236 4916 471100 4944
rect 471164 4916 569040 4944
rect 466236 4904 466242 4916
rect 327074 4836 327080 4888
rect 327132 4876 327138 4888
rect 361666 4876 361672 4888
rect 327132 4848 361672 4876
rect 327132 4836 327138 4848
rect 361666 4836 361672 4848
rect 361724 4836 361730 4888
rect 422202 4836 422208 4888
rect 422260 4876 422266 4888
rect 461213 4879 461271 4885
rect 461213 4876 461225 4879
rect 422260 4848 461225 4876
rect 422260 4836 422266 4848
rect 461213 4845 461225 4848
rect 461259 4845 461271 4879
rect 469122 4876 469128 4888
rect 461213 4839 461271 4845
rect 461596 4848 469128 4876
rect 325191 4780 326292 4808
rect 326617 4811 326675 4817
rect 325191 4777 325203 4780
rect 325145 4771 325203 4777
rect 326617 4777 326629 4811
rect 326663 4808 326675 4811
rect 327169 4811 327227 4817
rect 327169 4808 327181 4811
rect 326663 4780 327181 4808
rect 326663 4777 326675 4780
rect 326617 4771 326675 4777
rect 327169 4777 327181 4780
rect 327215 4777 327227 4811
rect 327169 4771 327227 4777
rect 328454 4768 328460 4820
rect 328512 4808 328518 4820
rect 363046 4808 363052 4820
rect 328512 4780 363052 4808
rect 328512 4768 328518 4780
rect 363046 4768 363052 4780
rect 363104 4768 363110 4820
rect 376757 4811 376815 4817
rect 376757 4777 376769 4811
rect 376803 4808 376815 4811
rect 381538 4808 381544 4820
rect 376803 4780 381544 4808
rect 376803 4777 376815 4780
rect 376757 4771 376815 4777
rect 381538 4768 381544 4780
rect 381596 4768 381602 4820
rect 423582 4768 423588 4820
rect 423640 4808 423646 4820
rect 461596 4808 461624 4848
rect 469122 4836 469128 4848
rect 469180 4836 469186 4888
rect 471072 4876 471100 4916
rect 569034 4904 569040 4916
rect 569092 4904 569098 4956
rect 572622 4876 572628 4888
rect 471072 4848 572628 4876
rect 572622 4836 572628 4848
rect 572680 4836 572686 4888
rect 423640 4780 461624 4808
rect 423640 4768 423646 4780
rect 462130 4768 462136 4820
rect 462188 4808 462194 4820
rect 471333 4811 471391 4817
rect 471333 4808 471345 4811
rect 462188 4780 471345 4808
rect 462188 4768 462194 4780
rect 471333 4777 471345 4780
rect 471379 4777 471391 4811
rect 471333 4771 471391 4777
rect 471425 4811 471483 4817
rect 471425 4777 471437 4811
rect 471471 4808 471483 4811
rect 579798 4808 579804 4820
rect 471471 4780 579804 4808
rect 471471 4777 471483 4780
rect 471425 4771 471483 4777
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 317371 4712 322980 4740
rect 317371 4709 317383 4712
rect 317325 4703 317383 4709
rect 324222 4700 324228 4752
rect 324280 4740 324286 4752
rect 359182 4740 359188 4752
rect 324280 4712 359188 4740
rect 324280 4700 324286 4712
rect 359182 4700 359188 4712
rect 359240 4700 359246 4752
rect 451090 4700 451096 4752
rect 451148 4740 451154 4752
rect 536926 4740 536932 4752
rect 451148 4712 536932 4740
rect 451148 4700 451154 4712
rect 536926 4700 536932 4712
rect 536984 4700 536990 4752
rect 215846 4632 215852 4684
rect 215904 4672 215910 4684
rect 317414 4672 317420 4684
rect 215904 4644 317420 4672
rect 215904 4632 215910 4644
rect 317414 4632 317420 4644
rect 317472 4632 317478 4684
rect 319441 4675 319499 4681
rect 319441 4641 319453 4675
rect 319487 4672 319499 4675
rect 322934 4672 322940 4684
rect 319487 4644 322940 4672
rect 319487 4641 319499 4644
rect 319441 4635 319499 4641
rect 322934 4632 322940 4644
rect 322992 4632 322998 4684
rect 326157 4675 326215 4681
rect 326157 4641 326169 4675
rect 326203 4672 326215 4675
rect 326203 4644 326384 4672
rect 326203 4641 326215 4644
rect 326157 4635 326215 4641
rect 219342 4564 219348 4616
rect 219400 4604 219406 4616
rect 318794 4604 318800 4616
rect 219400 4576 318800 4604
rect 219400 4564 219406 4576
rect 318794 4564 318800 4576
rect 318852 4564 318858 4616
rect 321554 4604 321560 4616
rect 318904 4576 321560 4604
rect 222930 4496 222936 4548
rect 222988 4536 222994 4548
rect 318904 4536 318932 4576
rect 321554 4564 321560 4576
rect 321612 4564 321618 4616
rect 322661 4607 322719 4613
rect 322661 4573 322673 4607
rect 322707 4604 322719 4607
rect 326249 4607 326307 4613
rect 326249 4604 326261 4607
rect 322707 4576 326261 4604
rect 322707 4573 322719 4576
rect 322661 4567 322719 4573
rect 326249 4573 326261 4576
rect 326295 4573 326307 4607
rect 326356 4604 326384 4644
rect 326522 4632 326528 4684
rect 326580 4672 326586 4684
rect 360286 4672 360292 4684
rect 326580 4644 360292 4672
rect 326580 4632 326586 4644
rect 360286 4632 360292 4644
rect 360344 4632 360350 4684
rect 449802 4632 449808 4684
rect 449860 4672 449866 4684
rect 533430 4672 533436 4684
rect 449860 4644 533436 4672
rect 449860 4632 449866 4644
rect 533430 4632 533436 4644
rect 533488 4632 533494 4684
rect 333974 4604 333980 4616
rect 326356 4576 333980 4604
rect 326249 4567 326307 4573
rect 333974 4564 333980 4576
rect 334032 4564 334038 4616
rect 448330 4564 448336 4616
rect 448388 4604 448394 4616
rect 529842 4604 529848 4616
rect 448388 4576 529848 4604
rect 448388 4564 448394 4576
rect 529842 4564 529848 4576
rect 529900 4564 529906 4616
rect 222988 4508 318932 4536
rect 222988 4496 222994 4508
rect 320358 4496 320364 4548
rect 320416 4536 320422 4548
rect 335354 4536 335360 4548
rect 320416 4508 335360 4536
rect 320416 4496 320422 4508
rect 335354 4496 335360 4508
rect 335412 4496 335418 4548
rect 447042 4496 447048 4548
rect 447100 4536 447106 4548
rect 526254 4536 526260 4548
rect 447100 4508 526260 4536
rect 447100 4496 447106 4508
rect 526254 4496 526260 4508
rect 526312 4496 526318 4548
rect 226518 4428 226524 4480
rect 226576 4468 226582 4480
rect 319441 4471 319499 4477
rect 319441 4468 319453 4471
rect 226576 4440 319453 4468
rect 226576 4428 226582 4440
rect 319441 4437 319453 4440
rect 319487 4437 319499 4471
rect 319441 4431 319499 4437
rect 322566 4428 322572 4480
rect 322624 4468 322630 4480
rect 337105 4471 337163 4477
rect 337105 4468 337117 4471
rect 322624 4440 337117 4468
rect 322624 4428 322630 4440
rect 337105 4437 337117 4440
rect 337151 4437 337163 4471
rect 337105 4431 337163 4437
rect 445570 4428 445576 4480
rect 445628 4468 445634 4480
rect 522666 4468 522672 4480
rect 445628 4440 522672 4468
rect 445628 4428 445634 4440
rect 522666 4428 522672 4440
rect 522724 4428 522730 4480
rect 201494 4360 201500 4412
rect 201552 4400 201558 4412
rect 271138 4400 271144 4412
rect 201552 4372 271144 4400
rect 201552 4360 201558 4372
rect 271138 4360 271144 4372
rect 271196 4360 271202 4412
rect 301406 4360 301412 4412
rect 301464 4400 301470 4412
rect 353478 4400 353484 4412
rect 301464 4372 353484 4400
rect 301464 4360 301470 4372
rect 353478 4360 353484 4372
rect 353536 4360 353542 4412
rect 376849 4403 376907 4409
rect 376849 4369 376861 4403
rect 376895 4400 376907 4403
rect 380158 4400 380164 4412
rect 376895 4372 380164 4400
rect 376895 4369 376907 4372
rect 376849 4363 376907 4369
rect 380158 4360 380164 4372
rect 380216 4360 380222 4412
rect 444282 4360 444288 4412
rect 444340 4400 444346 4412
rect 519078 4400 519084 4412
rect 444340 4372 519084 4400
rect 444340 4360 444346 4372
rect 519078 4360 519084 4372
rect 519136 4360 519142 4412
rect 205082 4292 205088 4344
rect 205140 4332 205146 4344
rect 272518 4332 272524 4344
rect 205140 4304 272524 4332
rect 205140 4292 205146 4304
rect 272518 4292 272524 4304
rect 272576 4292 272582 4344
rect 304994 4292 305000 4344
rect 305052 4332 305058 4344
rect 354950 4332 354956 4344
rect 305052 4304 354956 4332
rect 305052 4292 305058 4304
rect 354950 4292 354956 4304
rect 355008 4292 355014 4344
rect 442902 4292 442908 4344
rect 442960 4332 442966 4344
rect 515582 4332 515588 4344
rect 442960 4304 515588 4332
rect 442960 4292 442966 4304
rect 515582 4292 515588 4304
rect 515640 4292 515646 4344
rect 224129 4267 224187 4273
rect 224129 4233 224141 4267
rect 224175 4264 224187 4267
rect 230566 4264 230572 4276
rect 224175 4236 230572 4264
rect 224175 4233 224187 4236
rect 224129 4227 224187 4233
rect 230566 4224 230572 4236
rect 230624 4224 230630 4276
rect 249061 4267 249119 4273
rect 249061 4233 249073 4267
rect 249107 4264 249119 4267
rect 257985 4267 258043 4273
rect 257985 4264 257997 4267
rect 249107 4236 257997 4264
rect 249107 4233 249119 4236
rect 249061 4227 249119 4233
rect 257985 4233 257997 4236
rect 258031 4233 258043 4267
rect 257985 4227 258043 4233
rect 308582 4224 308588 4276
rect 308640 4264 308646 4276
rect 356146 4264 356152 4276
rect 308640 4236 356152 4264
rect 308640 4224 308646 4236
rect 356146 4224 356152 4236
rect 356204 4224 356210 4276
rect 437477 4267 437535 4273
rect 437477 4233 437489 4267
rect 437523 4264 437535 4267
rect 437523 4236 438348 4264
rect 437523 4233 437535 4236
rect 437477 4227 437535 4233
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 140866 4156 140872 4208
rect 140924 4196 140930 4208
rect 142062 4196 142068 4208
rect 140924 4168 142068 4196
rect 140924 4156 140930 4168
rect 142062 4156 142068 4168
rect 142120 4156 142126 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 160002 4196 160008 4208
rect 158772 4168 160008 4196
rect 158772 4156 158778 4168
rect 160002 4156 160008 4168
rect 160060 4156 160066 4208
rect 175366 4156 175372 4208
rect 175424 4196 175430 4208
rect 176562 4196 176568 4208
rect 175424 4168 176568 4196
rect 175424 4156 175430 4168
rect 176562 4156 176568 4168
rect 176620 4156 176626 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 307021 4199 307079 4205
rect 307021 4165 307033 4199
rect 307067 4196 307079 4199
rect 312078 4196 312084 4208
rect 307067 4168 312084 4196
rect 307067 4165 307079 4168
rect 307021 4159 307079 4165
rect 312078 4156 312084 4168
rect 312136 4156 312142 4208
rect 312170 4156 312176 4208
rect 312228 4196 312234 4208
rect 357710 4196 357716 4208
rect 312228 4168 357716 4196
rect 312228 4156 312234 4168
rect 357710 4156 357716 4168
rect 357768 4156 357774 4208
rect 417344 4168 418200 4196
rect 34974 4088 34980 4140
rect 35032 4128 35038 4140
rect 50338 4128 50344 4140
rect 35032 4100 50344 4128
rect 35032 4088 35038 4100
rect 50338 4088 50344 4100
rect 50396 4088 50402 4140
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 250438 4128 250444 4140
rect 57664 4100 250444 4128
rect 57664 4088 57670 4100
rect 250438 4088 250444 4100
rect 250496 4088 250502 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269022 4128 269028 4140
rect 268160 4100 269028 4128
rect 268160 4088 268166 4100
rect 269022 4088 269028 4100
rect 269080 4088 269086 4140
rect 269117 4131 269175 4137
rect 269117 4097 269129 4131
rect 269163 4128 269175 4131
rect 283101 4131 283159 4137
rect 283101 4128 283113 4131
rect 269163 4100 283113 4128
rect 269163 4097 269175 4100
rect 269117 4091 269175 4097
rect 283101 4097 283113 4100
rect 283147 4097 283159 4131
rect 283101 4091 283159 4097
rect 283193 4131 283251 4137
rect 283193 4097 283205 4131
rect 283239 4128 283251 4131
rect 295886 4128 295892 4140
rect 283239 4100 295892 4128
rect 283239 4097 283251 4100
rect 283193 4091 283251 4097
rect 295886 4088 295892 4100
rect 295944 4088 295950 4140
rect 296714 4088 296720 4140
rect 296772 4128 296778 4140
rect 297910 4128 297916 4140
rect 296772 4100 297916 4128
rect 296772 4088 296778 4100
rect 297910 4088 297916 4100
rect 297968 4088 297974 4140
rect 300302 4088 300308 4140
rect 300360 4128 300366 4140
rect 332321 4131 332379 4137
rect 332321 4128 332333 4131
rect 300360 4100 332333 4128
rect 300360 4088 300366 4100
rect 332321 4097 332333 4100
rect 332367 4097 332379 4131
rect 332321 4091 332379 4097
rect 332410 4088 332416 4140
rect 332468 4128 332474 4140
rect 333238 4128 333244 4140
rect 332468 4100 333244 4128
rect 332468 4088 332474 4100
rect 333238 4088 333244 4100
rect 333296 4088 333302 4140
rect 334710 4088 334716 4140
rect 334768 4128 334774 4140
rect 335262 4128 335268 4140
rect 334768 4100 335268 4128
rect 334768 4088 334774 4100
rect 335262 4088 335268 4100
rect 335320 4088 335326 4140
rect 335357 4131 335415 4137
rect 335357 4097 335369 4131
rect 335403 4128 335415 4131
rect 338758 4128 338764 4140
rect 335403 4100 338764 4128
rect 335403 4097 335415 4100
rect 335357 4091 335415 4097
rect 338758 4088 338764 4100
rect 338816 4088 338822 4140
rect 339494 4088 339500 4140
rect 339552 4128 339558 4140
rect 340782 4128 340788 4140
rect 339552 4100 340788 4128
rect 339552 4088 339558 4100
rect 340782 4088 340788 4100
rect 340840 4088 340846 4140
rect 340877 4131 340935 4137
rect 340877 4097 340889 4131
rect 340923 4128 340935 4131
rect 345658 4128 345664 4140
rect 340923 4100 345664 4128
rect 340923 4097 340935 4100
rect 340877 4091 340935 4097
rect 345658 4088 345664 4100
rect 345716 4088 345722 4140
rect 347866 4088 347872 4140
rect 347924 4128 347930 4140
rect 349062 4128 349068 4140
rect 347924 4100 349068 4128
rect 347924 4088 347930 4100
rect 349062 4088 349068 4100
rect 349120 4088 349126 4140
rect 349157 4131 349215 4137
rect 349157 4097 349169 4131
rect 349203 4128 349215 4131
rect 351178 4128 351184 4140
rect 349203 4100 351184 4128
rect 349203 4097 349215 4100
rect 349157 4091 349215 4097
rect 351178 4088 351184 4100
rect 351236 4088 351242 4140
rect 351362 4088 351368 4140
rect 351420 4128 351426 4140
rect 351822 4128 351828 4140
rect 351420 4100 351828 4128
rect 351420 4088 351426 4100
rect 351822 4088 351828 4100
rect 351880 4088 351886 4140
rect 351914 4088 351920 4140
rect 351972 4128 351978 4140
rect 352558 4128 352564 4140
rect 351972 4100 352564 4128
rect 351972 4088 351978 4100
rect 352558 4088 352564 4100
rect 352616 4088 352622 4140
rect 352653 4131 352711 4137
rect 352653 4097 352665 4131
rect 352699 4128 352711 4131
rect 355229 4131 355287 4137
rect 355229 4128 355241 4131
rect 352699 4100 355241 4128
rect 352699 4097 352711 4100
rect 352653 4091 352711 4097
rect 355229 4097 355241 4100
rect 355275 4097 355287 4131
rect 355229 4091 355287 4097
rect 355321 4131 355379 4137
rect 355321 4097 355333 4131
rect 355367 4128 355379 4131
rect 355367 4100 370360 4128
rect 355367 4097 355379 4100
rect 355321 4091 355379 4097
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 28258 4060 28264 4072
rect 20772 4032 28264 4060
rect 20772 4020 20778 4032
rect 28258 4020 28264 4032
rect 28316 4020 28322 4072
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 249058 4060 249064 4072
rect 50580 4032 249064 4060
rect 50580 4020 50586 4032
rect 249058 4020 249064 4032
rect 249116 4020 249122 4072
rect 261018 4020 261024 4072
rect 261076 4060 261082 4072
rect 297358 4060 297364 4072
rect 261076 4032 297364 4060
rect 261076 4020 261082 4032
rect 297358 4020 297364 4032
rect 297416 4020 297422 4072
rect 302602 4020 302608 4072
rect 302660 4060 302666 4072
rect 309778 4060 309784 4072
rect 302660 4032 309784 4060
rect 302660 4020 302666 4032
rect 309778 4020 309784 4032
rect 309836 4020 309842 4072
rect 314562 4020 314568 4072
rect 314620 4060 314626 4072
rect 358906 4060 358912 4072
rect 314620 4032 358912 4060
rect 314620 4020 314626 4032
rect 358906 4020 358912 4032
rect 358964 4020 358970 4072
rect 365714 4020 365720 4072
rect 365772 4060 365778 4072
rect 366910 4060 366916 4072
rect 365772 4032 366916 4060
rect 365772 4020 365778 4032
rect 366910 4020 366916 4032
rect 366968 4020 366974 4072
rect 369210 4020 369216 4072
rect 369268 4060 369274 4072
rect 369762 4060 369768 4072
rect 369268 4032 369768 4060
rect 369268 4020 369274 4032
rect 369762 4020 369768 4032
rect 369820 4020 369826 4072
rect 370332 4060 370360 4100
rect 370406 4088 370412 4140
rect 370464 4128 370470 4140
rect 371142 4128 371148 4140
rect 370464 4100 371148 4128
rect 370464 4088 370470 4100
rect 371142 4088 371148 4100
rect 371200 4088 371206 4140
rect 377582 4088 377588 4140
rect 377640 4128 377646 4140
rect 378042 4128 378048 4140
rect 377640 4100 378048 4128
rect 377640 4088 377646 4100
rect 378042 4088 378048 4100
rect 378100 4088 378106 4140
rect 378778 4088 378784 4140
rect 378836 4128 378842 4140
rect 378836 4100 379928 4128
rect 378836 4088 378842 4100
rect 372614 4060 372620 4072
rect 370332 4032 372620 4060
rect 372614 4020 372620 4032
rect 372672 4020 372678 4072
rect 376754 4020 376760 4072
rect 376812 4020 376818 4072
rect 46934 3952 46940 4004
rect 46992 3992 46998 4004
rect 248690 3992 248696 4004
rect 46992 3964 248696 3992
rect 46992 3952 46998 3964
rect 248690 3952 248696 3964
rect 248748 3952 248754 4004
rect 257430 3952 257436 4004
rect 257488 3992 257494 4004
rect 283193 3995 283251 4001
rect 283193 3992 283205 3995
rect 257488 3964 283205 3992
rect 257488 3952 257494 3964
rect 283193 3961 283205 3964
rect 283239 3961 283251 3995
rect 283193 3955 283251 3961
rect 283285 3995 283343 4001
rect 283285 3961 283297 3995
rect 283331 3992 283343 3995
rect 298094 3992 298100 4004
rect 283331 3964 298100 3992
rect 283331 3961 283343 3964
rect 283285 3955 283343 3961
rect 298094 3952 298100 3964
rect 298152 3952 298158 4004
rect 313366 3952 313372 4004
rect 313424 3992 313430 4004
rect 358814 3992 358820 4004
rect 313424 3964 358820 3992
rect 313424 3952 313430 3964
rect 358814 3952 358820 3964
rect 358872 3952 358878 4004
rect 359734 3952 359740 4004
rect 359792 3992 359798 4004
rect 376772 3992 376800 4020
rect 359792 3964 376800 3992
rect 359792 3952 359798 3964
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 247678 3924 247684 3936
rect 45796 3896 247684 3924
rect 45796 3884 45802 3896
rect 247678 3884 247684 3896
rect 247736 3884 247742 3936
rect 264606 3884 264612 3936
rect 264664 3924 264670 3936
rect 269117 3927 269175 3933
rect 269117 3924 269129 3927
rect 264664 3896 269129 3924
rect 264664 3884 264670 3896
rect 269117 3893 269129 3896
rect 269163 3893 269175 3927
rect 269117 3887 269175 3893
rect 275278 3884 275284 3936
rect 275336 3924 275342 3936
rect 275922 3924 275928 3936
rect 275336 3896 275928 3924
rect 275336 3884 275342 3896
rect 275922 3884 275928 3896
rect 275980 3884 275986 3936
rect 282454 3884 282460 3936
rect 282512 3924 282518 3936
rect 320821 3927 320879 3933
rect 320821 3924 320833 3927
rect 282512 3896 320833 3924
rect 282512 3884 282518 3896
rect 320821 3893 320833 3896
rect 320867 3893 320879 3927
rect 320821 3887 320879 3893
rect 320913 3927 320971 3933
rect 320913 3893 320925 3927
rect 320959 3924 320971 3927
rect 325602 3924 325608 3936
rect 320959 3896 325608 3924
rect 320959 3893 320971 3896
rect 320913 3887 320971 3893
rect 325602 3884 325608 3896
rect 325660 3884 325666 3936
rect 326341 3927 326399 3933
rect 326341 3893 326353 3927
rect 326387 3924 326399 3927
rect 332229 3927 332287 3933
rect 332229 3924 332241 3927
rect 326387 3896 332241 3924
rect 326387 3893 326399 3896
rect 326341 3887 326399 3893
rect 332229 3893 332241 3896
rect 332275 3893 332287 3927
rect 332229 3887 332287 3893
rect 332321 3927 332379 3933
rect 332321 3893 332333 3927
rect 332367 3924 332379 3927
rect 335909 3927 335967 3933
rect 332367 3896 335860 3924
rect 332367 3893 332379 3896
rect 332321 3887 332379 3893
rect 39758 3816 39764 3868
rect 39816 3856 39822 3868
rect 245930 3856 245936 3868
rect 39816 3828 245936 3856
rect 39816 3816 39822 3828
rect 245930 3816 245936 3828
rect 245988 3816 245994 3868
rect 289538 3816 289544 3868
rect 289596 3856 289602 3868
rect 335832 3856 335860 3896
rect 335909 3893 335921 3927
rect 335955 3924 335967 3927
rect 365806 3924 365812 3936
rect 335955 3896 365812 3924
rect 335955 3893 335967 3896
rect 335909 3887 335967 3893
rect 365806 3884 365812 3896
rect 365864 3884 365870 3936
rect 371602 3884 371608 3936
rect 371660 3924 371666 3936
rect 376757 3927 376815 3933
rect 376757 3924 376769 3927
rect 371660 3896 376769 3924
rect 371660 3884 371666 3896
rect 376757 3893 376769 3896
rect 376803 3893 376815 3927
rect 379900 3924 379928 4100
rect 379974 4088 379980 4140
rect 380032 4128 380038 4140
rect 380802 4128 380808 4140
rect 380032 4100 380808 4128
rect 380032 4088 380038 4100
rect 380802 4088 380808 4100
rect 380860 4088 380866 4140
rect 381170 4088 381176 4140
rect 381228 4128 381234 4140
rect 382182 4128 382188 4140
rect 381228 4100 382188 4128
rect 381228 4088 381234 4100
rect 382182 4088 382188 4100
rect 382240 4088 382246 4140
rect 383562 4088 383568 4140
rect 383620 4128 383626 4140
rect 384298 4128 384304 4140
rect 383620 4100 384304 4128
rect 383620 4088 383626 4100
rect 384298 4088 384304 4100
rect 384356 4088 384362 4140
rect 388254 4088 388260 4140
rect 388312 4128 388318 4140
rect 389082 4128 389088 4140
rect 388312 4100 389088 4128
rect 388312 4088 388318 4100
rect 389082 4088 389088 4100
rect 389140 4088 389146 4140
rect 385862 4020 385868 4072
rect 385920 4060 385926 4072
rect 387058 4060 387064 4072
rect 385920 4032 387064 4060
rect 385920 4020 385926 4032
rect 387058 4020 387064 4032
rect 387116 4020 387122 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 417344 4060 417372 4168
rect 418172 4137 418200 4168
rect 424962 4156 424968 4208
rect 425020 4196 425026 4208
rect 438213 4199 438271 4205
rect 438213 4196 438225 4199
rect 425020 4168 438225 4196
rect 425020 4156 425026 4168
rect 438213 4165 438225 4168
rect 438259 4165 438271 4199
rect 438213 4159 438271 4165
rect 418157 4131 418215 4137
rect 418157 4097 418169 4131
rect 418203 4097 418215 4131
rect 418157 4091 418215 4097
rect 427725 4131 427783 4137
rect 427725 4097 427737 4131
rect 427771 4128 427783 4131
rect 437474 4128 437480 4140
rect 427771 4100 437480 4128
rect 427771 4097 427783 4100
rect 427725 4091 427783 4097
rect 437474 4088 437480 4100
rect 437532 4088 437538 4140
rect 438320 4128 438348 4236
rect 441522 4224 441528 4276
rect 441580 4264 441586 4276
rect 511994 4264 512000 4276
rect 441580 4236 512000 4264
rect 441580 4224 441586 4236
rect 511994 4224 512000 4236
rect 512052 4224 512058 4276
rect 438397 4199 438455 4205
rect 438397 4165 438409 4199
rect 438443 4196 438455 4199
rect 472710 4196 472716 4208
rect 438443 4168 472716 4196
rect 438443 4165 438455 4168
rect 438397 4159 438455 4165
rect 472710 4156 472716 4168
rect 472768 4156 472774 4208
rect 445849 4131 445907 4137
rect 445849 4128 445861 4131
rect 438320 4100 445861 4128
rect 445849 4097 445861 4100
rect 445895 4097 445907 4131
rect 445849 4091 445907 4097
rect 451921 4131 451979 4137
rect 451921 4097 451933 4131
rect 451967 4128 451979 4131
rect 521470 4128 521476 4140
rect 451967 4100 521476 4128
rect 451967 4097 451979 4100
rect 451921 4091 451979 4097
rect 521470 4088 521476 4100
rect 521528 4088 521534 4140
rect 529198 4088 529204 4140
rect 529256 4128 529262 4140
rect 575014 4128 575020 4140
rect 529256 4100 575020 4128
rect 529256 4088 529262 4100
rect 575014 4088 575020 4100
rect 575072 4088 575078 4140
rect 439406 4060 439412 4072
rect 411220 4032 417372 4060
rect 417436 4032 439412 4060
rect 411220 4020 411226 4032
rect 382366 3952 382372 4004
rect 382424 3992 382430 4004
rect 386598 3992 386604 4004
rect 382424 3964 386604 3992
rect 382424 3952 382430 3964
rect 386598 3952 386604 3964
rect 386656 3952 386662 4004
rect 398098 3952 398104 4004
rect 398156 3992 398162 4004
rect 404906 3992 404912 4004
rect 398156 3964 404912 3992
rect 398156 3952 398162 3964
rect 404906 3952 404912 3964
rect 404964 3952 404970 4004
rect 411070 3952 411076 4004
rect 411128 3992 411134 4004
rect 417436 3992 417464 4032
rect 439406 4020 439412 4032
rect 439464 4020 439470 4072
rect 439590 4020 439596 4072
rect 439648 4060 439654 4072
rect 446769 4063 446827 4069
rect 446769 4060 446781 4063
rect 439648 4032 446781 4060
rect 439648 4020 439654 4032
rect 446769 4029 446781 4032
rect 446815 4029 446827 4063
rect 446769 4023 446827 4029
rect 448422 4020 448428 4072
rect 448480 4060 448486 4072
rect 528646 4060 528652 4072
rect 448480 4032 528652 4060
rect 448480 4020 448486 4032
rect 528646 4020 528652 4032
rect 528704 4020 528710 4072
rect 530578 4020 530584 4072
rect 530636 4060 530642 4072
rect 582190 4060 582196 4072
rect 530636 4032 582196 4060
rect 530636 4020 530642 4032
rect 582190 4020 582196 4032
rect 582248 4020 582254 4072
rect 411128 3964 417464 3992
rect 417513 3995 417571 4001
rect 411128 3952 411134 3964
rect 417513 3961 417525 3995
rect 417559 3992 417571 3995
rect 420089 3995 420147 4001
rect 420089 3992 420101 3995
rect 417559 3964 420101 3992
rect 417559 3961 417571 3964
rect 417513 3955 417571 3961
rect 420089 3961 420101 3964
rect 420135 3961 420147 3995
rect 420089 3955 420147 3961
rect 420178 3952 420184 4004
rect 420236 3992 420242 4004
rect 423950 3992 423956 4004
rect 420236 3964 423956 3992
rect 420236 3952 420242 3964
rect 423950 3952 423956 3964
rect 424008 3952 424014 4004
rect 424318 3952 424324 4004
rect 424376 3992 424382 4004
rect 425146 3992 425152 4004
rect 424376 3964 425152 3992
rect 424376 3952 424382 3964
rect 425146 3952 425152 3964
rect 425204 3952 425210 4004
rect 427078 3952 427084 4004
rect 427136 3992 427142 4004
rect 431126 3992 431132 4004
rect 427136 3964 431132 3992
rect 427136 3952 427142 3964
rect 431126 3952 431132 3964
rect 431184 3952 431190 4004
rect 433978 3952 433984 4004
rect 434036 3992 434042 4004
rect 435818 3992 435824 4004
rect 434036 3964 435824 3992
rect 434036 3952 434042 3964
rect 435818 3952 435824 3964
rect 435876 3952 435882 4004
rect 435913 3995 435971 4001
rect 435913 3961 435925 3995
rect 435959 3992 435971 3995
rect 437477 3995 437535 4001
rect 437477 3992 437489 3995
rect 435959 3964 437489 3992
rect 435959 3961 435971 3964
rect 435913 3955 435971 3961
rect 437477 3961 437489 3964
rect 437523 3961 437535 3995
rect 437477 3955 437535 3961
rect 456797 3995 456855 4001
rect 456797 3961 456809 3995
rect 456843 3992 456855 3995
rect 535730 3992 535736 4004
rect 456843 3964 535736 3992
rect 456843 3961 456855 3964
rect 456797 3955 456855 3961
rect 535730 3952 535736 3964
rect 535788 3952 535794 4004
rect 385310 3924 385316 3936
rect 379900 3896 385316 3924
rect 376757 3887 376815 3893
rect 385310 3884 385316 3896
rect 385368 3884 385374 3936
rect 404262 3884 404268 3936
rect 404320 3924 404326 3936
rect 410981 3927 411039 3933
rect 410981 3924 410993 3927
rect 404320 3896 410993 3924
rect 404320 3884 404326 3896
rect 410981 3893 410993 3896
rect 411027 3893 411039 3927
rect 410981 3887 411039 3893
rect 412542 3884 412548 3936
rect 412600 3924 412606 3936
rect 441798 3924 441804 3936
rect 412600 3896 441804 3924
rect 412600 3884 412606 3896
rect 441798 3884 441804 3896
rect 441856 3884 441862 3936
rect 453666 3924 453672 3936
rect 445496 3896 453672 3924
rect 342898 3856 342904 3868
rect 289596 3828 335768 3856
rect 335832 3828 342904 3856
rect 289596 3816 289602 3828
rect 19518 3748 19524 3800
rect 19576 3788 19582 3800
rect 32398 3788 32404 3800
rect 19576 3760 32404 3788
rect 19576 3748 19582 3760
rect 32398 3748 32404 3760
rect 32456 3748 32462 3800
rect 38562 3748 38568 3800
rect 38620 3788 38626 3800
rect 245746 3788 245752 3800
rect 38620 3760 245752 3788
rect 38620 3748 38626 3760
rect 245746 3748 245752 3760
rect 245804 3748 245810 3800
rect 278866 3748 278872 3800
rect 278924 3788 278930 3800
rect 285861 3791 285919 3797
rect 285861 3788 285873 3791
rect 278924 3760 285873 3788
rect 278924 3748 278930 3760
rect 285861 3757 285873 3760
rect 285907 3757 285919 3791
rect 285861 3751 285919 3757
rect 285950 3748 285956 3800
rect 286008 3788 286014 3800
rect 332137 3791 332195 3797
rect 332137 3788 332149 3791
rect 286008 3760 332149 3788
rect 286008 3748 286014 3760
rect 332137 3757 332149 3760
rect 332183 3757 332195 3791
rect 332137 3751 332195 3757
rect 332229 3791 332287 3797
rect 332229 3757 332241 3791
rect 332275 3788 332287 3791
rect 335538 3788 335544 3800
rect 332275 3760 335544 3788
rect 332275 3757 332287 3760
rect 332229 3751 332287 3757
rect 335538 3748 335544 3760
rect 335596 3748 335602 3800
rect 335740 3788 335768 3828
rect 342898 3816 342904 3828
rect 342956 3816 342962 3868
rect 343082 3816 343088 3868
rect 343140 3856 343146 3868
rect 369118 3856 369124 3868
rect 343140 3828 369124 3856
rect 343140 3816 343146 3828
rect 369118 3816 369124 3828
rect 369176 3816 369182 3868
rect 372798 3816 372804 3868
rect 372856 3856 372862 3868
rect 373902 3856 373908 3868
rect 372856 3828 373908 3856
rect 372856 3816 372862 3828
rect 373902 3816 373908 3828
rect 373960 3816 373966 3868
rect 407022 3816 407028 3868
rect 407080 3856 407086 3868
rect 407080 3828 412220 3856
rect 407080 3816 407086 3828
rect 341518 3788 341524 3800
rect 335740 3760 341524 3788
rect 341518 3748 341524 3760
rect 341576 3748 341582 3800
rect 341886 3748 341892 3800
rect 341944 3788 341950 3800
rect 370130 3788 370136 3800
rect 341944 3760 370136 3788
rect 341944 3748 341950 3760
rect 370130 3748 370136 3760
rect 370188 3748 370194 3800
rect 373994 3748 374000 3800
rect 374052 3788 374058 3800
rect 375282 3788 375288 3800
rect 374052 3760 375288 3788
rect 374052 3748 374058 3760
rect 375282 3748 375288 3760
rect 375340 3748 375346 3800
rect 399478 3748 399484 3800
rect 399536 3788 399542 3800
rect 408494 3788 408500 3800
rect 399536 3760 408500 3788
rect 399536 3748 399542 3760
rect 408494 3748 408500 3760
rect 408552 3748 408558 3800
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 243078 3720 243084 3732
rect 32732 3692 243084 3720
rect 32732 3680 32738 3692
rect 243078 3680 243084 3692
rect 243136 3680 243142 3732
rect 292485 3723 292543 3729
rect 292485 3689 292497 3723
rect 292531 3720 292543 3723
rect 326341 3723 326399 3729
rect 326341 3720 326353 3723
rect 292531 3692 326353 3720
rect 292531 3689 292543 3692
rect 292485 3683 292543 3689
rect 326341 3689 326353 3692
rect 326387 3689 326399 3723
rect 326341 3683 326399 3689
rect 326430 3680 326436 3732
rect 326488 3720 326494 3732
rect 328454 3720 328460 3732
rect 326488 3692 328460 3720
rect 326488 3680 326494 3692
rect 328454 3680 328460 3692
rect 328512 3680 328518 3732
rect 331214 3680 331220 3732
rect 331272 3720 331278 3732
rect 335909 3723 335967 3729
rect 335909 3720 335921 3723
rect 331272 3692 335921 3720
rect 331272 3680 331278 3692
rect 335909 3689 335921 3692
rect 335955 3689 335967 3723
rect 335909 3683 335967 3689
rect 338298 3680 338304 3732
rect 338356 3720 338362 3732
rect 361945 3723 362003 3729
rect 361945 3720 361957 3723
rect 338356 3692 361957 3720
rect 338356 3680 338362 3692
rect 361945 3689 361957 3692
rect 361991 3689 362003 3723
rect 361945 3683 362003 3689
rect 362037 3723 362095 3729
rect 362037 3689 362049 3723
rect 362083 3720 362095 3723
rect 370498 3720 370504 3732
rect 362083 3692 370504 3720
rect 362083 3689 362095 3692
rect 362037 3683 362095 3689
rect 370498 3680 370504 3692
rect 370556 3680 370562 3732
rect 375190 3680 375196 3732
rect 375248 3720 375254 3732
rect 383838 3720 383844 3732
rect 375248 3692 383844 3720
rect 375248 3680 375254 3692
rect 383838 3680 383844 3692
rect 383896 3680 383902 3732
rect 393130 3680 393136 3732
rect 393188 3720 393194 3732
rect 396626 3720 396632 3732
rect 393188 3692 396632 3720
rect 393188 3680 393194 3692
rect 396626 3680 396632 3692
rect 396684 3680 396690 3732
rect 400030 3680 400036 3732
rect 400088 3720 400094 3732
rect 412082 3720 412088 3732
rect 400088 3692 412088 3720
rect 400088 3680 400094 3692
rect 412082 3680 412088 3692
rect 412140 3680 412146 3732
rect 412192 3720 412220 3828
rect 413922 3816 413928 3868
rect 413980 3856 413986 3868
rect 445386 3856 445392 3868
rect 413980 3828 445392 3856
rect 413980 3816 413986 3828
rect 445386 3816 445392 3828
rect 445444 3816 445450 3868
rect 412450 3748 412456 3800
rect 412508 3788 412514 3800
rect 442994 3788 443000 3800
rect 412508 3760 443000 3788
rect 412508 3748 412514 3760
rect 442994 3748 443000 3760
rect 443052 3748 443058 3800
rect 417513 3723 417571 3729
rect 417513 3720 417525 3723
rect 412192 3692 417525 3720
rect 417513 3689 417525 3692
rect 417559 3689 417571 3723
rect 422113 3723 422171 3729
rect 422113 3720 422125 3723
rect 417513 3683 417571 3689
rect 417620 3692 422125 3720
rect 25498 3612 25504 3664
rect 25556 3652 25562 3664
rect 240318 3652 240324 3664
rect 25556 3624 240324 3652
rect 25556 3612 25562 3624
rect 240318 3612 240324 3624
rect 240376 3612 240382 3664
rect 262214 3612 262220 3664
rect 262272 3652 262278 3664
rect 322566 3652 322572 3664
rect 262272 3624 322572 3652
rect 262272 3612 262278 3624
rect 322566 3612 322572 3624
rect 322624 3612 322630 3664
rect 325234 3612 325240 3664
rect 325292 3652 325298 3664
rect 352837 3655 352895 3661
rect 352837 3652 352849 3655
rect 325292 3624 352849 3652
rect 325292 3612 325298 3624
rect 352837 3621 352849 3624
rect 352883 3621 352895 3655
rect 352837 3615 352895 3621
rect 352929 3655 352987 3661
rect 352929 3621 352941 3655
rect 352975 3652 352987 3655
rect 355318 3652 355324 3664
rect 352975 3624 355324 3652
rect 352975 3621 352987 3624
rect 352929 3615 352987 3621
rect 355318 3612 355324 3624
rect 355376 3612 355382 3664
rect 355413 3655 355471 3661
rect 355413 3621 355425 3655
rect 355459 3652 355471 3655
rect 358078 3652 358084 3664
rect 355459 3624 358084 3652
rect 355459 3621 355471 3624
rect 355413 3615 355471 3621
rect 358078 3612 358084 3624
rect 358136 3612 358142 3664
rect 360930 3612 360936 3664
rect 360988 3652 360994 3664
rect 377398 3652 377404 3664
rect 360988 3624 377404 3652
rect 360988 3612 360994 3624
rect 377398 3612 377404 3624
rect 377456 3612 377462 3664
rect 400122 3612 400128 3664
rect 400180 3652 400186 3664
rect 413186 3652 413192 3664
rect 400180 3624 413192 3652
rect 400180 3612 400186 3624
rect 413186 3612 413192 3624
rect 413244 3612 413250 3664
rect 416682 3612 416688 3664
rect 416740 3652 416746 3664
rect 417620 3652 417648 3692
rect 422113 3689 422125 3692
rect 422159 3689 422171 3723
rect 423033 3723 423091 3729
rect 423033 3720 423045 3723
rect 422113 3683 422171 3689
rect 422220 3692 423045 3720
rect 416740 3624 417648 3652
rect 416740 3612 416746 3624
rect 418062 3612 418068 3664
rect 418120 3652 418126 3664
rect 420730 3652 420736 3664
rect 418120 3624 420736 3652
rect 418120 3612 418126 3624
rect 420730 3612 420736 3624
rect 420788 3612 420794 3664
rect 420822 3612 420828 3664
rect 420880 3652 420886 3664
rect 422220 3652 422248 3692
rect 423033 3689 423045 3692
rect 423079 3689 423091 3723
rect 423033 3683 423091 3689
rect 423125 3723 423183 3729
rect 423125 3689 423137 3723
rect 423171 3720 423183 3723
rect 426437 3723 426495 3729
rect 426437 3720 426449 3723
rect 423171 3692 426449 3720
rect 423171 3689 423183 3692
rect 423125 3683 423183 3689
rect 426437 3689 426449 3692
rect 426483 3689 426495 3723
rect 426437 3683 426495 3689
rect 428200 3692 428412 3720
rect 420880 3624 422248 3652
rect 422941 3655 422999 3661
rect 420880 3612 420886 3624
rect 422941 3621 422953 3655
rect 422987 3652 422999 3655
rect 428200 3652 428228 3692
rect 422987 3624 428228 3652
rect 428384 3652 428412 3692
rect 428458 3680 428464 3732
rect 428516 3720 428522 3732
rect 430025 3723 430083 3729
rect 430025 3720 430037 3723
rect 428516 3692 430037 3720
rect 428516 3680 428522 3692
rect 430025 3689 430037 3692
rect 430071 3689 430083 3723
rect 430025 3683 430083 3689
rect 430117 3723 430175 3729
rect 430117 3689 430129 3723
rect 430163 3720 430175 3723
rect 441709 3723 441767 3729
rect 441709 3720 441721 3723
rect 430163 3692 441721 3720
rect 430163 3689 430175 3692
rect 430117 3683 430175 3689
rect 441709 3689 441721 3692
rect 441755 3689 441767 3723
rect 445496 3720 445524 3896
rect 453666 3884 453672 3896
rect 453724 3884 453730 3936
rect 453942 3884 453948 3936
rect 454000 3924 454006 3936
rect 542906 3924 542912 3936
rect 454000 3896 542912 3924
rect 454000 3884 454006 3896
rect 542906 3884 542912 3896
rect 542964 3884 542970 3936
rect 445662 3816 445668 3868
rect 445720 3856 445726 3868
rect 451921 3859 451979 3865
rect 451921 3856 451933 3859
rect 445720 3828 451933 3856
rect 445720 3816 445726 3828
rect 451921 3825 451933 3828
rect 451967 3825 451979 3859
rect 451921 3819 451979 3825
rect 456702 3816 456708 3868
rect 456760 3856 456766 3868
rect 550082 3856 550088 3868
rect 456760 3828 550088 3856
rect 456760 3816 456766 3828
rect 550082 3816 550088 3828
rect 550140 3816 550146 3868
rect 445849 3791 445907 3797
rect 445849 3757 445861 3791
rect 445895 3788 445907 3791
rect 459646 3788 459652 3800
rect 445895 3760 459652 3788
rect 445895 3757 445907 3760
rect 445849 3751 445907 3757
rect 459646 3748 459652 3760
rect 459704 3748 459710 3800
rect 460014 3748 460020 3800
rect 460072 3788 460078 3800
rect 463234 3788 463240 3800
rect 460072 3760 463240 3788
rect 460072 3748 460078 3760
rect 463234 3748 463240 3760
rect 463292 3748 463298 3800
rect 466365 3791 466423 3797
rect 466365 3788 466377 3791
rect 463344 3760 466377 3788
rect 441709 3683 441767 3689
rect 442184 3692 445524 3720
rect 442184 3652 442212 3692
rect 451182 3680 451188 3732
rect 451240 3720 451246 3732
rect 456797 3723 456855 3729
rect 456797 3720 456809 3723
rect 451240 3692 456809 3720
rect 451240 3680 451246 3692
rect 456797 3689 456809 3692
rect 456843 3689 456855 3723
rect 456797 3683 456855 3689
rect 456889 3723 456947 3729
rect 456889 3689 456901 3723
rect 456935 3720 456947 3723
rect 456935 3692 457392 3720
rect 456935 3689 456947 3692
rect 456889 3683 456947 3689
rect 428384 3624 442212 3652
rect 422987 3621 422999 3624
rect 422941 3615 422999 3621
rect 442258 3612 442264 3664
rect 442316 3652 442322 3664
rect 449897 3655 449955 3661
rect 449897 3652 449909 3655
rect 442316 3624 449909 3652
rect 442316 3612 442322 3624
rect 449897 3621 449909 3624
rect 449943 3621 449955 3655
rect 449897 3615 449955 3621
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 19978 3584 19984 3596
rect 11296 3556 19984 3584
rect 11296 3544 11302 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 239030 3584 239036 3596
rect 24360 3556 239036 3584
rect 24360 3544 24366 3556
rect 239030 3544 239036 3556
rect 239088 3544 239094 3596
rect 265802 3544 265808 3596
rect 265860 3584 265866 3596
rect 320729 3587 320787 3593
rect 320729 3584 320741 3587
rect 265860 3556 320741 3584
rect 265860 3544 265866 3556
rect 320729 3553 320741 3556
rect 320775 3553 320787 3587
rect 320729 3547 320787 3553
rect 320821 3587 320879 3593
rect 320821 3553 320833 3587
rect 320867 3584 320879 3587
rect 322753 3587 322811 3593
rect 322753 3584 322765 3587
rect 320867 3556 322765 3584
rect 320867 3553 320879 3556
rect 320821 3547 320879 3553
rect 322753 3553 322765 3556
rect 322799 3553 322811 3587
rect 322753 3547 322811 3553
rect 322842 3544 322848 3596
rect 322900 3584 322906 3596
rect 327074 3584 327080 3596
rect 322900 3556 327080 3584
rect 322900 3544 322906 3556
rect 327074 3544 327080 3556
rect 327132 3544 327138 3596
rect 332137 3587 332195 3593
rect 332137 3553 332149 3587
rect 332183 3584 332195 3587
rect 335357 3587 335415 3593
rect 335357 3584 335369 3587
rect 332183 3556 335369 3584
rect 332183 3553 332195 3556
rect 332137 3547 332195 3553
rect 335357 3553 335369 3556
rect 335403 3553 335415 3587
rect 335357 3547 335415 3553
rect 335725 3587 335783 3593
rect 335725 3553 335737 3587
rect 335771 3584 335783 3587
rect 363598 3584 363604 3596
rect 335771 3556 363604 3584
rect 335771 3553 335783 3556
rect 335725 3547 335783 3553
rect 363598 3544 363604 3556
rect 363656 3544 363662 3596
rect 402238 3544 402244 3596
rect 402296 3584 402302 3596
rect 415670 3584 415676 3596
rect 402296 3556 415676 3584
rect 402296 3544 402302 3556
rect 415670 3544 415676 3556
rect 415728 3544 415734 3596
rect 417418 3544 417424 3596
rect 417476 3544 417482 3596
rect 434530 3544 434536 3596
rect 434588 3584 434594 3596
rect 434625 3587 434683 3593
rect 434625 3584 434637 3587
rect 434588 3556 434637 3584
rect 434588 3544 434594 3556
rect 434625 3553 434637 3556
rect 434671 3584 434683 3587
rect 454681 3587 454739 3593
rect 454681 3584 454693 3587
rect 434671 3556 454693 3584
rect 434671 3553 434683 3556
rect 434625 3547 434683 3553
rect 454681 3553 454693 3556
rect 454727 3553 454739 3587
rect 457364 3584 457392 3692
rect 463344 3652 463372 3760
rect 466365 3757 466377 3760
rect 466411 3757 466423 3791
rect 466365 3751 466423 3757
rect 466917 3791 466975 3797
rect 466917 3757 466929 3791
rect 466963 3788 466975 3791
rect 557166 3788 557172 3800
rect 466963 3760 557172 3788
rect 466963 3757 466975 3760
rect 466917 3751 466975 3757
rect 557166 3748 557172 3760
rect 557224 3748 557230 3800
rect 564342 3720 564348 3732
rect 460032 3624 463372 3652
rect 463436 3692 564348 3720
rect 460032 3584 460060 3624
rect 457364 3556 460060 3584
rect 454681 3547 454739 3553
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 236270 3516 236276 3528
rect 16080 3488 236276 3516
rect 16080 3476 16086 3488
rect 236270 3476 236276 3488
rect 236328 3476 236334 3528
rect 258626 3476 258632 3528
rect 258684 3516 258690 3528
rect 320358 3516 320364 3528
rect 258684 3488 320364 3516
rect 258684 3476 258690 3488
rect 320358 3476 320364 3488
rect 320416 3476 320422 3528
rect 320450 3476 320456 3528
rect 320508 3516 320514 3528
rect 321462 3516 321468 3528
rect 320508 3488 321468 3516
rect 320508 3476 320514 3488
rect 321462 3476 321468 3488
rect 321520 3476 321526 3528
rect 324038 3476 324044 3528
rect 324096 3516 324102 3528
rect 363138 3516 363144 3528
rect 324096 3488 363144 3516
rect 324096 3476 324102 3488
rect 363138 3476 363144 3488
rect 363196 3476 363202 3528
rect 368658 3516 368664 3528
rect 363248 3488 368664 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 234890 3448 234896 3460
rect 14884 3420 234896 3448
rect 14884 3408 14890 3420
rect 234890 3408 234896 3420
rect 234948 3408 234954 3460
rect 255038 3408 255044 3460
rect 255096 3448 255102 3460
rect 318702 3448 318708 3460
rect 255096 3420 318708 3448
rect 255096 3408 255102 3420
rect 318702 3408 318708 3420
rect 318760 3408 318766 3460
rect 321646 3408 321652 3460
rect 321704 3448 321710 3460
rect 361850 3448 361856 3460
rect 321704 3420 361856 3448
rect 321704 3408 321710 3420
rect 361850 3408 361856 3420
rect 361908 3408 361914 3460
rect 361945 3451 362003 3457
rect 361945 3417 361957 3451
rect 361991 3448 362003 3451
rect 363248 3448 363276 3488
rect 368658 3476 368664 3488
rect 368716 3476 368722 3528
rect 376757 3519 376815 3525
rect 376757 3516 376769 3519
rect 370240 3488 376769 3516
rect 361991 3420 363276 3448
rect 361991 3417 362003 3420
rect 361945 3411 362003 3417
rect 368014 3408 368020 3460
rect 368072 3448 368078 3460
rect 370240 3448 370268 3488
rect 376757 3485 376769 3488
rect 376803 3485 376815 3519
rect 376757 3479 376815 3485
rect 390830 3476 390836 3528
rect 390888 3516 390894 3528
rect 391842 3516 391848 3528
rect 390888 3488 391848 3516
rect 390888 3476 390894 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 394510 3476 394516 3528
rect 394568 3516 394574 3528
rect 400214 3516 400220 3528
rect 394568 3488 400220 3516
rect 394568 3476 394574 3488
rect 400214 3476 400220 3488
rect 400272 3476 400278 3528
rect 402882 3476 402888 3528
rect 402940 3516 402946 3528
rect 413189 3519 413247 3525
rect 413189 3516 413201 3519
rect 402940 3488 413201 3516
rect 402940 3476 402946 3488
rect 413189 3485 413201 3488
rect 413235 3485 413247 3519
rect 413189 3479 413247 3485
rect 413278 3476 413284 3528
rect 413336 3516 413342 3528
rect 414474 3516 414480 3528
rect 413336 3488 414480 3516
rect 413336 3476 413342 3488
rect 414474 3476 414480 3488
rect 414532 3476 414538 3528
rect 417436 3516 417464 3544
rect 418062 3516 418068 3528
rect 417436 3488 418068 3516
rect 418062 3476 418068 3488
rect 418120 3476 418126 3528
rect 420089 3519 420147 3525
rect 420089 3485 420101 3519
rect 420135 3516 420147 3519
rect 423033 3519 423091 3525
rect 420135 3488 422892 3516
rect 420135 3485 420147 3488
rect 420089 3479 420147 3485
rect 379698 3448 379704 3460
rect 368072 3420 370268 3448
rect 376128 3420 379704 3448
rect 368072 3408 368078 3420
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 35158 3380 35164 3392
rect 29144 3352 35164 3380
rect 29144 3340 29150 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 39298 3380 39304 3392
rect 36228 3352 39304 3380
rect 36228 3340 36234 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 45465 3383 45523 3389
rect 45465 3349 45477 3383
rect 45511 3380 45523 3383
rect 45511 3352 58296 3380
rect 45511 3349 45523 3352
rect 45465 3343 45523 3349
rect 10042 3272 10048 3324
rect 10100 3312 10106 3324
rect 13078 3312 13084 3324
rect 10100 3284 13084 3312
rect 10100 3272 10106 3284
rect 13078 3272 13084 3284
rect 13136 3272 13142 3324
rect 42150 3272 42156 3324
rect 42208 3312 42214 3324
rect 57238 3312 57244 3324
rect 42208 3284 57244 3312
rect 42208 3272 42214 3284
rect 57238 3272 57244 3284
rect 57296 3272 57302 3324
rect 58268 3312 58296 3352
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 251818 3380 251824 3392
rect 71792 3352 251824 3380
rect 61378 3312 61384 3324
rect 58268 3284 61384 3312
rect 61378 3272 61384 3284
rect 61436 3272 61442 3324
rect 52822 3204 52828 3256
rect 52880 3244 52886 3256
rect 53742 3244 53748 3256
rect 52880 3216 53748 3244
rect 52880 3204 52886 3216
rect 53742 3204 53748 3216
rect 53800 3204 53806 3256
rect 54018 3204 54024 3256
rect 54076 3244 54082 3256
rect 54076 3216 59676 3244
rect 54076 3204 54082 3216
rect 43346 3136 43352 3188
rect 43404 3176 43410 3188
rect 45465 3179 45523 3185
rect 45465 3176 45477 3179
rect 43404 3148 45477 3176
rect 43404 3136 43410 3148
rect 45465 3145 45477 3148
rect 45511 3145 45523 3179
rect 45465 3139 45523 3145
rect 59648 3108 59676 3216
rect 64782 3204 64788 3256
rect 64840 3244 64846 3256
rect 71792 3244 71820 3352
rect 251818 3340 251824 3352
rect 251876 3340 251882 3392
rect 282825 3383 282883 3389
rect 282825 3349 282837 3383
rect 282871 3380 282883 3383
rect 289814 3380 289820 3392
rect 282871 3352 289820 3380
rect 282871 3349 282883 3352
rect 282825 3343 282883 3349
rect 289814 3340 289820 3352
rect 289872 3340 289878 3392
rect 299106 3340 299112 3392
rect 299164 3380 299170 3392
rect 302878 3380 302884 3392
rect 299164 3352 302884 3380
rect 299164 3340 299170 3352
rect 302878 3340 302884 3352
rect 302936 3340 302942 3392
rect 310974 3340 310980 3392
rect 311032 3380 311038 3392
rect 344373 3383 344431 3389
rect 344373 3380 344385 3383
rect 311032 3352 344385 3380
rect 311032 3340 311038 3352
rect 344373 3349 344385 3352
rect 344419 3349 344431 3383
rect 344373 3343 344431 3349
rect 345661 3383 345719 3389
rect 345661 3349 345673 3383
rect 345707 3380 345719 3383
rect 352929 3383 352987 3389
rect 352929 3380 352941 3383
rect 345707 3352 352941 3380
rect 345707 3349 345719 3352
rect 345661 3343 345719 3349
rect 352929 3349 352941 3352
rect 352975 3349 352987 3383
rect 352929 3343 352987 3349
rect 353754 3340 353760 3392
rect 353812 3380 353818 3392
rect 375466 3380 375472 3392
rect 353812 3352 375472 3380
rect 353812 3340 353818 3352
rect 375466 3340 375472 3352
rect 375524 3340 375530 3392
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 253198 3312 253204 3324
rect 71924 3284 253204 3312
rect 71924 3272 71930 3284
rect 253198 3272 253204 3284
rect 253256 3272 253262 3324
rect 276400 3284 284708 3312
rect 64840 3216 71820 3244
rect 71884 3216 74580 3244
rect 64840 3204 64846 3216
rect 61194 3136 61200 3188
rect 61252 3176 61258 3188
rect 61252 3148 67956 3176
rect 61252 3136 61258 3148
rect 66898 3108 66904 3120
rect 59648 3080 66904 3108
rect 66898 3068 66904 3080
rect 66956 3068 66962 3120
rect 67928 3108 67956 3148
rect 68278 3136 68284 3188
rect 68336 3176 68342 3188
rect 71884 3176 71912 3216
rect 68336 3148 71912 3176
rect 68336 3136 68342 3148
rect 71038 3108 71044 3120
rect 67928 3080 71044 3108
rect 71038 3068 71044 3080
rect 71096 3068 71102 3120
rect 74552 3040 74580 3216
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 84838 3244 84844 3256
rect 82832 3216 84844 3244
rect 75454 3136 75460 3188
rect 75512 3176 75518 3188
rect 79318 3176 79324 3188
rect 75512 3148 79324 3176
rect 75512 3136 75518 3148
rect 79318 3136 79324 3148
rect 79376 3136 79382 3188
rect 82630 3136 82636 3188
rect 82688 3176 82694 3188
rect 82832 3176 82860 3216
rect 84838 3204 84844 3216
rect 84896 3204 84902 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 88518 3204 88524 3256
rect 88576 3244 88582 3256
rect 89622 3244 89628 3256
rect 88576 3216 89628 3244
rect 88576 3204 88582 3216
rect 89622 3204 89628 3216
rect 89680 3204 89686 3256
rect 254578 3244 254584 3256
rect 89732 3216 254584 3244
rect 82688 3148 82860 3176
rect 82909 3179 82967 3185
rect 82688 3136 82694 3148
rect 82909 3145 82921 3179
rect 82955 3176 82967 3179
rect 89732 3176 89760 3216
rect 254578 3204 254584 3216
rect 254636 3204 254642 3256
rect 269298 3204 269304 3256
rect 269356 3244 269362 3256
rect 276293 3247 276351 3253
rect 276293 3244 276305 3247
rect 269356 3216 276305 3244
rect 269356 3204 269362 3216
rect 276293 3213 276305 3216
rect 276339 3213 276351 3247
rect 276293 3207 276351 3213
rect 255958 3176 255964 3188
rect 82955 3148 89760 3176
rect 94424 3148 255964 3176
rect 82955 3145 82967 3148
rect 82909 3139 82967 3145
rect 89714 3068 89720 3120
rect 89772 3108 89778 3120
rect 94424 3108 94452 3148
rect 255958 3136 255964 3148
rect 256016 3136 256022 3188
rect 272886 3136 272892 3188
rect 272944 3176 272950 3188
rect 276400 3176 276428 3284
rect 276474 3204 276480 3256
rect 276532 3244 276538 3256
rect 284680 3244 284708 3284
rect 284754 3272 284760 3324
rect 284812 3312 284818 3324
rect 285582 3312 285588 3324
rect 284812 3284 285588 3312
rect 284812 3272 284818 3284
rect 285582 3272 285588 3284
rect 285640 3272 285646 3324
rect 285861 3315 285919 3321
rect 285861 3281 285873 3315
rect 285907 3312 285919 3315
rect 292485 3315 292543 3321
rect 292485 3312 292497 3315
rect 285907 3284 292497 3312
rect 285907 3281 285919 3284
rect 285861 3275 285919 3281
rect 292485 3281 292497 3284
rect 292531 3281 292543 3315
rect 292485 3275 292543 3281
rect 303798 3272 303804 3324
rect 303856 3312 303862 3324
rect 344278 3312 344284 3324
rect 303856 3284 344284 3312
rect 303856 3272 303862 3284
rect 344278 3272 344284 3284
rect 344336 3272 344342 3324
rect 345477 3315 345535 3321
rect 345477 3281 345489 3315
rect 345523 3312 345535 3315
rect 349157 3315 349215 3321
rect 349157 3312 349169 3315
rect 345523 3284 349169 3312
rect 345523 3281 345535 3284
rect 345477 3275 345535 3281
rect 349157 3281 349169 3284
rect 349203 3281 349215 3315
rect 349157 3275 349215 3281
rect 350258 3272 350264 3324
rect 350316 3312 350322 3324
rect 374270 3312 374276 3324
rect 350316 3284 374276 3312
rect 350316 3272 350322 3284
rect 374270 3272 374276 3284
rect 374328 3272 374334 3324
rect 288434 3244 288440 3256
rect 276532 3216 284616 3244
rect 284680 3216 288440 3244
rect 276532 3204 276538 3216
rect 272944 3148 276428 3176
rect 272944 3136 272950 3148
rect 277670 3136 277676 3188
rect 277728 3176 277734 3188
rect 284588 3176 284616 3216
rect 288434 3204 288440 3216
rect 288492 3204 288498 3256
rect 291930 3204 291936 3256
rect 291988 3244 291994 3256
rect 316678 3244 316684 3256
rect 291988 3216 316684 3244
rect 291988 3204 291994 3216
rect 316678 3204 316684 3216
rect 316736 3204 316742 3256
rect 318058 3204 318064 3256
rect 318116 3244 318122 3256
rect 343913 3247 343971 3253
rect 343913 3244 343925 3247
rect 318116 3216 343925 3244
rect 318116 3204 318122 3216
rect 343913 3213 343925 3216
rect 343959 3213 343971 3247
rect 343913 3207 343971 3213
rect 344097 3247 344155 3253
rect 344097 3213 344109 3247
rect 344143 3244 344155 3247
rect 348418 3244 348424 3256
rect 344143 3216 348424 3244
rect 344143 3213 344155 3216
rect 344097 3207 344155 3213
rect 348418 3204 348424 3216
rect 348476 3204 348482 3256
rect 349062 3204 349068 3256
rect 349120 3244 349126 3256
rect 355321 3247 355379 3253
rect 355321 3244 355333 3247
rect 349120 3216 355333 3244
rect 349120 3204 349126 3216
rect 355321 3213 355333 3216
rect 355367 3213 355379 3247
rect 355321 3207 355379 3213
rect 355413 3247 355471 3253
rect 355413 3213 355425 3247
rect 355459 3244 355471 3247
rect 356698 3244 356704 3256
rect 355459 3216 356704 3244
rect 355459 3213 355471 3216
rect 355413 3207 355471 3213
rect 356698 3204 356704 3216
rect 356756 3204 356762 3256
rect 357342 3204 357348 3256
rect 357400 3244 357406 3256
rect 376018 3244 376024 3256
rect 357400 3216 376024 3244
rect 357400 3204 357406 3216
rect 376018 3204 376024 3216
rect 376076 3204 376082 3256
rect 288526 3176 288532 3188
rect 277728 3148 284524 3176
rect 284588 3148 288532 3176
rect 277728 3136 277734 3148
rect 89772 3080 94452 3108
rect 89772 3068 89778 3080
rect 94498 3068 94504 3120
rect 94556 3108 94562 3120
rect 95142 3108 95148 3120
rect 94556 3080 95148 3108
rect 94556 3068 94562 3080
rect 95142 3068 95148 3080
rect 95200 3068 95206 3120
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 98086 3068 98092 3120
rect 98144 3108 98150 3120
rect 99190 3108 99196 3120
rect 98144 3080 99196 3108
rect 98144 3068 98150 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 101582 3068 101588 3120
rect 101640 3108 101646 3120
rect 102042 3108 102048 3120
rect 101640 3080 102048 3108
rect 101640 3068 101646 3080
rect 102042 3068 102048 3080
rect 102100 3068 102106 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 105170 3068 105176 3120
rect 105228 3108 105234 3120
rect 106182 3108 106188 3120
rect 105228 3080 106188 3108
rect 105228 3068 105234 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107470 3108 107476 3120
rect 106424 3080 107476 3108
rect 106424 3068 106430 3080
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 257338 3108 257344 3120
rect 108316 3080 257344 3108
rect 77938 3040 77944 3052
rect 74552 3012 77944 3040
rect 77938 3000 77944 3012
rect 77996 3000 78002 3052
rect 93302 3000 93308 3052
rect 93360 3040 93366 3052
rect 102594 3040 102600 3052
rect 93360 3012 102600 3040
rect 93360 3000 93366 3012
rect 102594 3000 102600 3012
rect 102652 3000 102658 3052
rect 79042 2932 79048 2984
rect 79100 2972 79106 2984
rect 82909 2975 82967 2981
rect 82909 2972 82921 2975
rect 79100 2944 82921 2972
rect 79100 2932 79106 2944
rect 82909 2941 82921 2944
rect 82955 2941 82967 2975
rect 82909 2935 82967 2941
rect 86126 2932 86132 2984
rect 86184 2972 86190 2984
rect 93857 2975 93915 2981
rect 93857 2972 93869 2975
rect 86184 2944 93869 2972
rect 86184 2932 86190 2944
rect 93857 2941 93869 2944
rect 93903 2941 93915 2975
rect 93857 2935 93915 2941
rect 96890 2932 96896 2984
rect 96948 2972 96954 2984
rect 108316 2972 108344 3080
rect 257338 3068 257344 3080
rect 257396 3068 257402 3120
rect 284496 3108 284524 3148
rect 288526 3136 288532 3148
rect 288584 3136 288590 3188
rect 309778 3136 309784 3188
rect 309836 3176 309842 3188
rect 335817 3179 335875 3185
rect 335817 3176 335829 3179
rect 309836 3148 335829 3176
rect 309836 3136 309842 3148
rect 335817 3145 335829 3148
rect 335863 3145 335875 3179
rect 335817 3139 335875 3145
rect 335906 3136 335912 3188
rect 335964 3176 335970 3188
rect 340601 3179 340659 3185
rect 340601 3176 340613 3179
rect 335964 3148 340613 3176
rect 335964 3136 335970 3148
rect 340601 3145 340613 3148
rect 340647 3145 340659 3179
rect 340601 3139 340659 3145
rect 340690 3136 340696 3188
rect 340748 3176 340754 3188
rect 345661 3179 345719 3185
rect 345661 3176 345673 3179
rect 340748 3148 345673 3176
rect 340748 3136 340754 3148
rect 345661 3145 345673 3148
rect 345707 3145 345719 3179
rect 345661 3139 345719 3145
rect 346670 3136 346676 3188
rect 346728 3176 346734 3188
rect 362037 3179 362095 3185
rect 362037 3176 362049 3179
rect 346728 3148 362049 3176
rect 346728 3136 346734 3148
rect 362037 3145 362049 3148
rect 362083 3145 362095 3179
rect 362037 3139 362095 3145
rect 362126 3136 362132 3188
rect 362184 3176 362190 3188
rect 362862 3176 362868 3188
rect 362184 3148 362868 3176
rect 362184 3136 362190 3148
rect 362862 3136 362868 3148
rect 362920 3136 362926 3188
rect 363322 3136 363328 3188
rect 363380 3176 363386 3188
rect 364242 3176 364248 3188
rect 363380 3148 364248 3176
rect 363380 3136 363386 3148
rect 364242 3136 364248 3148
rect 364300 3136 364306 3188
rect 364518 3136 364524 3188
rect 364576 3176 364582 3188
rect 365717 3179 365775 3185
rect 365717 3176 365729 3179
rect 364576 3148 365729 3176
rect 364576 3136 364582 3148
rect 365717 3145 365729 3148
rect 365763 3145 365775 3179
rect 365717 3139 365775 3145
rect 290458 3108 290464 3120
rect 284496 3080 290464 3108
rect 290458 3068 290464 3080
rect 290516 3068 290522 3120
rect 295518 3068 295524 3120
rect 295576 3108 295582 3120
rect 319438 3108 319444 3120
rect 295576 3080 319444 3108
rect 295576 3068 295582 3080
rect 319438 3068 319444 3080
rect 319496 3068 319502 3120
rect 322753 3111 322811 3117
rect 322753 3077 322765 3111
rect 322799 3108 322811 3111
rect 327718 3108 327724 3120
rect 322799 3080 327724 3108
rect 322799 3077 322811 3080
rect 322753 3071 322811 3077
rect 327718 3068 327724 3080
rect 327776 3068 327782 3120
rect 328822 3068 328828 3120
rect 328880 3108 328886 3120
rect 362218 3108 362224 3120
rect 328880 3080 362224 3108
rect 328880 3068 328886 3080
rect 362218 3068 362224 3080
rect 362276 3068 362282 3120
rect 375285 3111 375343 3117
rect 375285 3077 375297 3111
rect 375331 3108 375343 3111
rect 376128 3108 376156 3420
rect 379698 3408 379704 3420
rect 379756 3408 379762 3460
rect 406378 3408 406384 3460
rect 406436 3448 406442 3460
rect 410886 3448 410892 3460
rect 406436 3420 410892 3448
rect 406436 3408 406442 3420
rect 410886 3408 410892 3420
rect 410944 3408 410950 3460
rect 410981 3451 411039 3457
rect 410981 3417 410993 3451
rect 411027 3448 411039 3451
rect 422754 3448 422760 3460
rect 411027 3420 422760 3448
rect 411027 3417 411039 3420
rect 410981 3411 411039 3417
rect 422754 3408 422760 3420
rect 422812 3408 422818 3460
rect 422864 3448 422892 3488
rect 423033 3485 423045 3519
rect 423079 3516 423091 3519
rect 460842 3516 460848 3528
rect 423079 3488 460848 3516
rect 423079 3485 423091 3488
rect 423033 3479 423091 3485
rect 460842 3476 460848 3488
rect 460900 3476 460906 3528
rect 462222 3476 462228 3528
rect 462280 3516 462286 3528
rect 463436 3516 463464 3692
rect 564342 3680 564348 3692
rect 564400 3680 564406 3732
rect 463602 3612 463608 3664
rect 463660 3652 463666 3664
rect 566734 3652 566740 3664
rect 463660 3624 566740 3652
rect 463660 3612 463666 3624
rect 566734 3612 566740 3624
rect 566792 3612 566798 3664
rect 466362 3544 466368 3596
rect 466420 3584 466426 3596
rect 571426 3584 571432 3596
rect 466420 3556 571432 3584
rect 466420 3544 466426 3556
rect 571426 3544 571432 3556
rect 571484 3544 571490 3596
rect 462280 3488 463464 3516
rect 462280 3476 462286 3488
rect 466270 3476 466276 3528
rect 466328 3516 466334 3528
rect 573818 3516 573824 3528
rect 466328 3488 573824 3516
rect 466328 3476 466334 3488
rect 573818 3476 573824 3488
rect 573876 3476 573882 3528
rect 429930 3448 429936 3460
rect 422864 3420 429936 3448
rect 429930 3408 429936 3420
rect 429988 3408 429994 3460
rect 430025 3451 430083 3457
rect 430025 3417 430037 3451
rect 430071 3448 430083 3451
rect 432509 3451 432567 3457
rect 432509 3448 432521 3451
rect 430071 3420 432521 3448
rect 430071 3417 430083 3420
rect 430025 3411 430083 3417
rect 432509 3417 432521 3420
rect 432555 3417 432567 3451
rect 432509 3411 432567 3417
rect 432601 3451 432659 3457
rect 432601 3417 432613 3451
rect 432647 3448 432659 3451
rect 467926 3448 467932 3460
rect 432647 3420 467932 3448
rect 432647 3417 432659 3420
rect 432601 3411 432659 3417
rect 467926 3408 467932 3420
rect 467984 3408 467990 3460
rect 469030 3408 469036 3460
rect 469088 3448 469094 3460
rect 578602 3448 578608 3460
rect 469088 3420 578608 3448
rect 469088 3408 469094 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 403618 3340 403624 3392
rect 403676 3380 403682 3392
rect 407298 3380 407304 3392
rect 403676 3352 407304 3380
rect 403676 3340 403682 3352
rect 407298 3340 407304 3352
rect 407356 3340 407362 3392
rect 409782 3340 409788 3392
rect 409840 3380 409846 3392
rect 437014 3380 437020 3392
rect 409840 3352 437020 3380
rect 409840 3340 409846 3352
rect 437014 3340 437020 3352
rect 437072 3340 437078 3392
rect 437474 3340 437480 3392
rect 437532 3380 437538 3392
rect 438210 3380 438216 3392
rect 437532 3352 438216 3380
rect 437532 3340 437538 3352
rect 438210 3340 438216 3352
rect 438268 3340 438274 3392
rect 443638 3340 443644 3392
rect 443696 3380 443702 3392
rect 443696 3352 510108 3380
rect 443696 3340 443702 3352
rect 395982 3272 395988 3324
rect 396040 3312 396046 3324
rect 402514 3312 402520 3324
rect 396040 3284 402520 3312
rect 396040 3272 396046 3284
rect 402514 3272 402520 3284
rect 402572 3272 402578 3324
rect 402790 3272 402796 3324
rect 402848 3312 402854 3324
rect 419166 3312 419172 3324
rect 402848 3284 419172 3312
rect 402848 3272 402854 3284
rect 419166 3272 419172 3284
rect 419224 3272 419230 3324
rect 420270 3272 420276 3324
rect 420328 3312 420334 3324
rect 446582 3312 446588 3324
rect 420328 3284 446588 3312
rect 420328 3272 420334 3284
rect 446582 3272 446588 3284
rect 446640 3272 446646 3324
rect 503622 3312 503628 3324
rect 446692 3284 503628 3312
rect 409138 3204 409144 3256
rect 409196 3244 409202 3256
rect 423125 3247 423183 3253
rect 423125 3244 423137 3247
rect 409196 3216 423137 3244
rect 409196 3204 409202 3216
rect 423125 3213 423137 3216
rect 423171 3213 423183 3247
rect 423125 3207 423183 3213
rect 431218 3204 431224 3256
rect 431276 3244 431282 3256
rect 435913 3247 435971 3253
rect 435913 3244 435925 3247
rect 431276 3216 435925 3244
rect 431276 3204 431282 3216
rect 435913 3213 435925 3216
rect 435959 3213 435971 3247
rect 435913 3207 435971 3213
rect 442350 3204 442356 3256
rect 442408 3244 442414 3256
rect 446692 3244 446720 3284
rect 503622 3272 503628 3284
rect 503680 3272 503686 3324
rect 510080 3312 510108 3352
rect 514018 3340 514024 3392
rect 514076 3380 514082 3392
rect 517882 3380 517888 3392
rect 514076 3352 517888 3380
rect 514076 3340 514082 3352
rect 517882 3340 517888 3352
rect 517940 3340 517946 3392
rect 525058 3380 525064 3392
rect 517992 3352 525064 3380
rect 514386 3312 514392 3324
rect 510080 3284 514392 3312
rect 514386 3272 514392 3284
rect 514444 3272 514450 3324
rect 516870 3272 516876 3324
rect 516928 3312 516934 3324
rect 517992 3312 518020 3352
rect 525058 3340 525064 3352
rect 525116 3340 525122 3392
rect 527818 3340 527824 3392
rect 527876 3380 527882 3392
rect 567838 3380 567844 3392
rect 527876 3352 567844 3380
rect 527876 3340 527882 3352
rect 567838 3340 567844 3352
rect 567896 3340 567902 3392
rect 577406 3312 577412 3324
rect 516928 3284 518020 3312
rect 518084 3284 577412 3312
rect 516928 3272 516934 3284
rect 442408 3216 446720 3244
rect 446769 3247 446827 3253
rect 442408 3204 442414 3216
rect 446769 3213 446781 3247
rect 446815 3244 446827 3247
rect 496538 3244 496544 3256
rect 446815 3216 496544 3244
rect 446815 3213 446827 3216
rect 446769 3207 446827 3213
rect 496538 3204 496544 3216
rect 496596 3204 496602 3256
rect 512638 3204 512644 3256
rect 512696 3244 512702 3256
rect 518084 3244 518112 3284
rect 577406 3272 577412 3284
rect 577464 3272 577470 3324
rect 512696 3216 518112 3244
rect 518161 3247 518219 3253
rect 512696 3204 512702 3216
rect 518161 3213 518173 3247
rect 518207 3244 518219 3247
rect 570230 3244 570236 3256
rect 518207 3216 570236 3244
rect 518207 3213 518219 3216
rect 518161 3207 518219 3213
rect 570230 3204 570236 3216
rect 570288 3204 570294 3256
rect 405642 3136 405648 3188
rect 405700 3176 405706 3188
rect 426342 3176 426348 3188
rect 405700 3148 426348 3176
rect 405700 3136 405706 3148
rect 426342 3136 426348 3148
rect 426400 3136 426406 3188
rect 426437 3179 426495 3185
rect 426437 3145 426449 3179
rect 426483 3176 426495 3179
rect 432322 3176 432328 3188
rect 426483 3148 432328 3176
rect 426483 3145 426495 3148
rect 426437 3139 426495 3145
rect 432322 3136 432328 3148
rect 432380 3136 432386 3188
rect 432432 3148 477632 3176
rect 375331 3080 376156 3108
rect 375331 3077 375343 3080
rect 375285 3071 375343 3077
rect 393222 3068 393228 3120
rect 393280 3108 393286 3120
rect 395430 3108 395436 3120
rect 393280 3080 395436 3108
rect 393280 3068 393286 3080
rect 395430 3068 395436 3080
rect 395488 3068 395494 3120
rect 404998 3068 405004 3120
rect 405056 3108 405062 3120
rect 416866 3108 416872 3120
rect 405056 3080 416872 3108
rect 405056 3068 405062 3080
rect 416866 3068 416872 3080
rect 416924 3068 416930 3120
rect 422941 3111 422999 3117
rect 422941 3108 422953 3111
rect 416976 3080 422953 3108
rect 258718 3040 258724 3052
rect 96948 2944 108344 2972
rect 108408 3012 258724 3040
rect 96948 2932 96954 2944
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 108408 2904 108436 3012
rect 258718 3000 258724 3012
rect 258776 3000 258782 3052
rect 276293 3043 276351 3049
rect 276293 3009 276305 3043
rect 276339 3040 276351 3043
rect 282825 3043 282883 3049
rect 282825 3040 282837 3043
rect 276339 3012 282837 3040
rect 276339 3009 276351 3012
rect 276293 3003 276351 3009
rect 282825 3009 282837 3012
rect 282871 3009 282883 3043
rect 282825 3003 282883 3009
rect 293126 3000 293132 3052
rect 293184 3040 293190 3052
rect 312538 3040 312544 3052
rect 293184 3012 312544 3040
rect 293184 3000 293190 3012
rect 312538 3000 312544 3012
rect 312596 3000 312602 3052
rect 315758 3000 315764 3052
rect 315816 3040 315822 3052
rect 324222 3040 324228 3052
rect 315816 3012 324228 3040
rect 315816 3000 315822 3012
rect 324222 3000 324228 3012
rect 324280 3000 324286 3052
rect 327626 3000 327632 3052
rect 327684 3040 327690 3052
rect 335725 3043 335783 3049
rect 335725 3040 335737 3043
rect 327684 3012 335737 3040
rect 327684 3000 327690 3012
rect 335725 3009 335737 3012
rect 335771 3009 335783 3043
rect 335725 3003 335783 3009
rect 335906 3000 335912 3052
rect 335964 3040 335970 3052
rect 367278 3040 367284 3052
rect 335964 3012 367284 3040
rect 335964 3000 335970 3012
rect 367278 3000 367284 3012
rect 367336 3000 367342 3052
rect 376386 3000 376392 3052
rect 376444 3040 376450 3052
rect 381630 3040 381636 3052
rect 376444 3012 381636 3040
rect 376444 3000 376450 3012
rect 381630 3000 381636 3012
rect 381688 3000 381694 3052
rect 394602 3000 394608 3052
rect 394660 3040 394666 3052
rect 399018 3040 399024 3052
rect 394660 3012 399024 3040
rect 394660 3000 394666 3012
rect 399018 3000 399024 3012
rect 399076 3000 399082 3052
rect 112346 2932 112352 2984
rect 112404 2972 112410 2984
rect 113082 2972 113088 2984
rect 112404 2944 113088 2972
rect 112404 2932 112410 2944
rect 113082 2932 113088 2944
rect 113140 2932 113146 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 115934 2932 115940 2984
rect 115992 2972 115998 2984
rect 116946 2972 116952 2984
rect 115992 2944 116952 2972
rect 115992 2932 115998 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 119430 2932 119436 2984
rect 119488 2972 119494 2984
rect 119982 2972 119988 2984
rect 119488 2944 119988 2972
rect 119488 2932 119494 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 258810 2972 258816 2984
rect 121472 2944 258816 2972
rect 104032 2876 108436 2904
rect 104032 2864 104038 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 121472 2904 121500 2944
rect 258810 2932 258816 2944
rect 258868 2932 258874 2984
rect 316954 2932 316960 2984
rect 317012 2972 317018 2984
rect 335633 2975 335691 2981
rect 335633 2972 335645 2975
rect 317012 2944 335645 2972
rect 317012 2932 317018 2944
rect 335633 2941 335645 2944
rect 335679 2941 335691 2975
rect 335633 2935 335691 2941
rect 335817 2975 335875 2981
rect 335817 2941 335829 2975
rect 335863 2972 335875 2975
rect 344186 2972 344192 2984
rect 335863 2944 344192 2972
rect 335863 2941 335875 2944
rect 335817 2935 335875 2941
rect 344186 2932 344192 2944
rect 344244 2932 344250 2984
rect 344373 2975 344431 2981
rect 344373 2941 344385 2975
rect 344419 2972 344431 2975
rect 347777 2975 347835 2981
rect 347777 2972 347789 2975
rect 344419 2944 347789 2972
rect 344419 2941 344431 2944
rect 344373 2935 344431 2941
rect 347777 2941 347789 2944
rect 347823 2941 347835 2975
rect 347777 2935 347835 2941
rect 350077 2975 350135 2981
rect 350077 2941 350089 2975
rect 350123 2972 350135 2975
rect 351914 2972 351920 2984
rect 350123 2944 351920 2972
rect 350123 2941 350135 2944
rect 350077 2935 350135 2941
rect 351914 2932 351920 2944
rect 351972 2932 351978 2984
rect 352558 2932 352564 2984
rect 352616 2972 352622 2984
rect 374086 2972 374092 2984
rect 352616 2944 374092 2972
rect 352616 2932 352622 2944
rect 374086 2932 374092 2944
rect 374144 2932 374150 2984
rect 395890 2932 395896 2984
rect 395948 2972 395954 2984
rect 401318 2972 401324 2984
rect 395948 2944 401324 2972
rect 395948 2932 395954 2944
rect 401318 2932 401324 2944
rect 401376 2932 401382 2984
rect 416590 2932 416596 2984
rect 416648 2972 416654 2984
rect 416976 2972 417004 3080
rect 422941 3077 422953 3080
rect 422987 3077 422999 3111
rect 422941 3071 422999 3077
rect 423033 3111 423091 3117
rect 423033 3077 423045 3111
rect 423079 3108 423091 3111
rect 427725 3111 427783 3117
rect 427725 3108 427737 3111
rect 423079 3080 427737 3108
rect 423079 3077 423091 3080
rect 423033 3071 423091 3077
rect 427725 3077 427737 3080
rect 427771 3077 427783 3111
rect 427725 3071 427783 3077
rect 431310 3068 431316 3120
rect 431368 3108 431374 3120
rect 432432 3108 432460 3148
rect 431368 3080 432460 3108
rect 432509 3111 432567 3117
rect 431368 3068 431374 3080
rect 432509 3077 432521 3111
rect 432555 3108 432567 3111
rect 475102 3108 475108 3120
rect 432555 3080 475108 3108
rect 432555 3077 432567 3080
rect 432509 3071 432567 3077
rect 475102 3068 475108 3080
rect 475160 3068 475166 3120
rect 475378 3068 475384 3120
rect 475436 3108 475442 3120
rect 477494 3108 477500 3120
rect 475436 3080 477500 3108
rect 475436 3068 475442 3080
rect 477494 3068 477500 3080
rect 477552 3068 477558 3120
rect 477604 3108 477632 3148
rect 505738 3136 505744 3188
rect 505796 3176 505802 3188
rect 563146 3176 563152 3188
rect 505796 3148 563152 3176
rect 505796 3136 505802 3148
rect 563146 3136 563152 3148
rect 563204 3136 563210 3188
rect 482278 3108 482284 3120
rect 477604 3080 482284 3108
rect 482278 3068 482284 3080
rect 482336 3068 482342 3120
rect 524966 3068 524972 3120
rect 525024 3108 525030 3120
rect 560754 3108 560760 3120
rect 525024 3080 560760 3108
rect 525024 3068 525030 3080
rect 560754 3068 560760 3080
rect 560812 3068 560818 3120
rect 421558 3000 421564 3052
rect 421616 3040 421622 3052
rect 450170 3040 450176 3052
rect 421616 3012 450176 3040
rect 421616 3000 421622 3012
rect 450170 3000 450176 3012
rect 450228 3000 450234 3052
rect 450265 3043 450323 3049
rect 450265 3009 450277 3043
rect 450311 3040 450323 3043
rect 489362 3040 489368 3052
rect 450311 3012 489368 3040
rect 450311 3009 450323 3012
rect 450265 3003 450323 3009
rect 489362 3000 489368 3012
rect 489420 3000 489426 3052
rect 509878 3000 509884 3052
rect 509936 3040 509942 3052
rect 518161 3043 518219 3049
rect 518161 3040 518173 3043
rect 509936 3012 518173 3040
rect 509936 3000 509942 3012
rect 518161 3009 518173 3012
rect 518207 3009 518219 3043
rect 518161 3003 518219 3009
rect 523678 3000 523684 3052
rect 523736 3040 523742 3052
rect 553578 3040 553584 3052
rect 523736 3012 553584 3040
rect 523736 3000 523742 3012
rect 553578 3000 553584 3012
rect 553636 3000 553642 3052
rect 416648 2944 417004 2972
rect 416648 2932 416654 2944
rect 418062 2932 418068 2984
rect 418120 2972 418126 2984
rect 428734 2972 428740 2984
rect 418120 2944 428740 2972
rect 418120 2932 418126 2944
rect 428734 2932 428740 2944
rect 428792 2932 428798 2984
rect 429838 2932 429844 2984
rect 429896 2972 429902 2984
rect 448974 2972 448980 2984
rect 429896 2944 448980 2972
rect 429896 2932 429902 2944
rect 448974 2932 448980 2944
rect 449032 2932 449038 2984
rect 449897 2975 449955 2981
rect 449897 2941 449909 2975
rect 449943 2972 449955 2975
rect 481082 2972 481088 2984
rect 449943 2944 481088 2972
rect 449943 2941 449955 2944
rect 449897 2935 449955 2941
rect 481082 2932 481088 2944
rect 481140 2932 481146 2984
rect 520918 2932 520924 2984
rect 520976 2972 520982 2984
rect 546494 2972 546500 2984
rect 520976 2944 546500 2972
rect 520976 2932 520982 2944
rect 546494 2932 546500 2944
rect 546552 2932 546558 2984
rect 260098 2904 260104 2916
rect 111208 2876 121500 2904
rect 121564 2876 260104 2904
rect 111208 2864 111214 2876
rect 93857 2839 93915 2845
rect 93857 2805 93869 2839
rect 93903 2836 93915 2839
rect 95878 2836 95884 2848
rect 93903 2808 95884 2836
rect 93903 2805 93915 2808
rect 93857 2799 93915 2805
rect 95878 2796 95884 2808
rect 95936 2796 95942 2848
rect 114738 2796 114744 2848
rect 114796 2836 114802 2848
rect 121564 2836 121592 2876
rect 260098 2864 260104 2876
rect 260156 2864 260162 2916
rect 319254 2864 319260 2916
rect 319312 2904 319318 2916
rect 326522 2904 326528 2916
rect 319312 2876 326528 2904
rect 319312 2864 319318 2876
rect 326522 2864 326528 2876
rect 326580 2864 326586 2916
rect 340693 2907 340751 2913
rect 340693 2873 340705 2907
rect 340739 2904 340751 2907
rect 344097 2907 344155 2913
rect 344097 2904 344109 2907
rect 340739 2876 344109 2904
rect 340739 2873 340751 2876
rect 340693 2867 340751 2873
rect 344097 2873 344109 2876
rect 344143 2873 344155 2907
rect 344097 2867 344155 2873
rect 344278 2864 344284 2916
rect 344336 2904 344342 2916
rect 352653 2907 352711 2913
rect 352653 2904 352665 2907
rect 344336 2876 352665 2904
rect 344336 2864 344342 2876
rect 352653 2873 352665 2876
rect 352699 2873 352711 2907
rect 354861 2907 354919 2913
rect 354861 2904 354873 2907
rect 352653 2867 352711 2873
rect 352760 2876 354873 2904
rect 114796 2808 121592 2836
rect 114796 2796 114802 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 261478 2836 261484 2848
rect 121880 2808 261484 2836
rect 121880 2796 121886 2808
rect 261478 2796 261484 2808
rect 261536 2796 261542 2848
rect 330018 2796 330024 2848
rect 330076 2836 330082 2848
rect 335538 2836 335544 2848
rect 330076 2808 335544 2836
rect 330076 2796 330082 2808
rect 335538 2796 335544 2808
rect 335596 2796 335602 2848
rect 335633 2839 335691 2845
rect 335633 2805 335645 2839
rect 335679 2836 335691 2839
rect 340785 2839 340843 2845
rect 340785 2836 340797 2839
rect 335679 2808 340797 2836
rect 335679 2805 335691 2808
rect 335633 2799 335691 2805
rect 340785 2805 340797 2808
rect 340831 2805 340843 2839
rect 340785 2799 340843 2805
rect 343913 2839 343971 2845
rect 343913 2805 343925 2839
rect 343959 2836 343971 2839
rect 352760 2836 352788 2876
rect 354861 2873 354873 2876
rect 354907 2873 354919 2907
rect 354861 2867 354919 2873
rect 354950 2864 354956 2916
rect 355008 2904 355014 2916
rect 355962 2904 355968 2916
rect 355008 2876 355968 2904
rect 355008 2864 355014 2876
rect 355962 2864 355968 2876
rect 356020 2864 356026 2916
rect 359458 2904 359464 2916
rect 356072 2876 359464 2904
rect 343959 2808 352788 2836
rect 352837 2839 352895 2845
rect 343959 2805 343971 2808
rect 343913 2799 343971 2805
rect 352837 2805 352849 2839
rect 352883 2836 352895 2839
rect 356072 2836 356100 2876
rect 359458 2864 359464 2876
rect 359516 2864 359522 2916
rect 365717 2907 365775 2913
rect 365717 2873 365729 2907
rect 365763 2904 365775 2907
rect 375285 2907 375343 2913
rect 375285 2904 375297 2907
rect 365763 2876 375297 2904
rect 365763 2873 365775 2876
rect 365717 2867 365775 2873
rect 375285 2873 375297 2876
rect 375331 2873 375343 2907
rect 375285 2867 375343 2873
rect 398190 2864 398196 2916
rect 398248 2904 398254 2916
rect 403710 2904 403716 2916
rect 398248 2876 403716 2904
rect 398248 2864 398254 2876
rect 403710 2864 403716 2876
rect 403768 2864 403774 2916
rect 413189 2907 413247 2913
rect 413189 2873 413201 2907
rect 413235 2904 413247 2907
rect 420362 2904 420368 2916
rect 413235 2876 420368 2904
rect 413235 2873 413247 2876
rect 413189 2867 413247 2873
rect 420362 2864 420368 2876
rect 420420 2864 420426 2916
rect 423033 2907 423091 2913
rect 423033 2904 423045 2907
rect 420472 2876 423045 2904
rect 352883 2808 356100 2836
rect 352883 2805 352895 2808
rect 352837 2799 352895 2805
rect 356146 2796 356152 2848
rect 356204 2836 356210 2848
rect 375558 2836 375564 2848
rect 356204 2808 375564 2836
rect 356204 2796 356210 2808
rect 375558 2796 375564 2808
rect 375616 2796 375622 2848
rect 388438 2836 388444 2848
rect 387076 2808 388444 2836
rect 387076 2780 387104 2808
rect 388438 2796 388444 2808
rect 388496 2796 388502 2848
rect 418157 2839 418215 2845
rect 418157 2805 418169 2839
rect 418203 2836 418215 2839
rect 420472 2836 420500 2876
rect 423033 2873 423045 2876
rect 423079 2873 423091 2907
rect 423033 2867 423091 2873
rect 424410 2864 424416 2916
rect 424468 2904 424474 2916
rect 432601 2907 432659 2913
rect 432601 2904 432613 2907
rect 424468 2876 432613 2904
rect 424468 2864 424474 2876
rect 432601 2873 432613 2876
rect 432647 2873 432659 2907
rect 432601 2867 432659 2873
rect 438118 2864 438124 2916
rect 438176 2904 438182 2916
rect 438176 2876 446444 2904
rect 438176 2864 438182 2876
rect 418203 2808 420500 2836
rect 422113 2839 422171 2845
rect 418203 2805 418215 2808
rect 418157 2799 418215 2805
rect 422113 2805 422125 2839
rect 422159 2836 422171 2839
rect 422159 2808 429792 2836
rect 422159 2805 422171 2808
rect 422113 2799 422171 2805
rect 347777 2771 347835 2777
rect 347777 2737 347789 2771
rect 347823 2768 347835 2771
rect 350077 2771 350135 2777
rect 350077 2768 350089 2771
rect 347823 2740 350089 2768
rect 347823 2737 347835 2740
rect 347777 2731 347835 2737
rect 350077 2737 350089 2740
rect 350123 2737 350135 2771
rect 350077 2731 350135 2737
rect 387058 2728 387064 2780
rect 387116 2728 387122 2780
rect 429764 2768 429792 2808
rect 439498 2796 439504 2848
rect 439556 2836 439562 2848
rect 441709 2839 441767 2845
rect 439556 2808 441476 2836
rect 439556 2796 439562 2808
rect 430117 2771 430175 2777
rect 430117 2768 430129 2771
rect 429764 2740 430129 2768
rect 430117 2737 430129 2740
rect 430163 2737 430175 2771
rect 441448 2768 441476 2808
rect 441709 2805 441721 2839
rect 441755 2836 441767 2839
rect 444837 2839 444895 2845
rect 444837 2836 444849 2839
rect 441755 2808 444849 2836
rect 441755 2805 441767 2808
rect 441709 2799 441767 2805
rect 444837 2805 444849 2808
rect 444883 2805 444895 2839
rect 446416 2836 446444 2876
rect 449158 2864 449164 2916
rect 449216 2904 449222 2916
rect 450265 2907 450323 2913
rect 450265 2904 450277 2907
rect 449216 2876 450277 2904
rect 449216 2864 449222 2876
rect 450265 2873 450277 2876
rect 450311 2873 450323 2907
rect 456797 2907 456855 2913
rect 456797 2904 456809 2907
rect 450265 2867 450323 2873
rect 451292 2876 456809 2904
rect 451185 2839 451243 2845
rect 451185 2836 451197 2839
rect 446416 2808 451197 2836
rect 444837 2799 444895 2805
rect 451185 2805 451197 2808
rect 451231 2805 451243 2839
rect 451185 2799 451243 2805
rect 441448 2740 441660 2768
rect 430117 2731 430175 2737
rect 441632 2700 441660 2740
rect 451292 2700 451320 2876
rect 456797 2873 456809 2876
rect 456843 2873 456855 2907
rect 456797 2867 456855 2873
rect 460290 2864 460296 2916
rect 460348 2904 460354 2916
rect 466181 2907 466239 2913
rect 466181 2904 466193 2907
rect 460348 2876 466193 2904
rect 460348 2864 460354 2876
rect 466181 2873 466193 2876
rect 466227 2873 466239 2907
rect 466181 2867 466239 2873
rect 466365 2907 466423 2913
rect 466365 2873 466377 2907
rect 466411 2904 466423 2907
rect 473906 2904 473912 2916
rect 466411 2876 473912 2904
rect 466411 2873 466423 2876
rect 466365 2867 466423 2873
rect 473906 2864 473912 2876
rect 473964 2864 473970 2916
rect 521010 2864 521016 2916
rect 521068 2904 521074 2916
rect 539318 2904 539324 2916
rect 521068 2876 539324 2904
rect 521068 2864 521074 2876
rect 539318 2864 539324 2876
rect 539376 2864 539382 2916
rect 451461 2839 451519 2845
rect 451461 2805 451473 2839
rect 451507 2836 451519 2839
rect 466822 2836 466828 2848
rect 451507 2808 466828 2836
rect 451507 2805 451519 2808
rect 451461 2799 451519 2805
rect 466822 2796 466828 2808
rect 466880 2796 466886 2848
rect 466917 2839 466975 2845
rect 466917 2805 466929 2839
rect 466963 2836 466975 2839
rect 466963 2808 466997 2836
rect 466963 2805 466975 2808
rect 466917 2799 466975 2805
rect 466181 2771 466239 2777
rect 466181 2737 466193 2771
rect 466227 2768 466239 2771
rect 466932 2768 466960 2799
rect 518158 2796 518164 2848
rect 518216 2836 518222 2848
rect 532234 2836 532240 2848
rect 518216 2808 532240 2836
rect 518216 2796 518222 2808
rect 532234 2796 532240 2808
rect 532292 2796 532298 2848
rect 466227 2740 466960 2768
rect 466227 2737 466239 2740
rect 466181 2731 466239 2737
rect 441632 2672 451320 2700
rect 454681 2159 454739 2165
rect 454681 2125 454693 2159
rect 454727 2156 454739 2159
rect 457254 2156 457260 2168
rect 454727 2128 457260 2156
rect 454727 2125 454739 2128
rect 454681 2119 454739 2125
rect 457254 2116 457260 2128
rect 457312 2116 457318 2168
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 164694 552 164700 604
rect 164752 592 164758 604
rect 165522 592 165528 604
rect 164752 564 165528 592
rect 164752 552 164758 564
rect 165522 552 165528 564
rect 165580 552 165586 604
rect 165890 552 165896 604
rect 165948 592 165954 604
rect 166902 592 166908 604
rect 165948 564 166908 592
rect 165948 552 165954 564
rect 166902 552 166908 564
rect 166960 552 166966 604
rect 169386 552 169392 604
rect 169444 592 169450 604
rect 169662 592 169668 604
rect 169444 564 169668 592
rect 169444 552 169450 564
rect 169662 552 169668 564
rect 169720 552 169726 604
rect 182542 552 182548 604
rect 182600 592 182606 604
rect 183462 592 183468 604
rect 182600 564 183468 592
rect 182600 552 182606 564
rect 183462 552 183468 564
rect 183520 552 183526 604
rect 183738 552 183744 604
rect 183796 592 183802 604
rect 184750 592 184756 604
rect 183796 564 184756 592
rect 183796 552 183802 564
rect 184750 552 184756 564
rect 184808 552 184814 604
rect 187234 552 187240 604
rect 187292 592 187298 604
rect 187602 592 187608 604
rect 187292 564 187608 592
rect 187292 552 187298 564
rect 187602 552 187608 564
rect 187660 552 187666 604
rect 189626 552 189632 604
rect 189684 592 189690 604
rect 190362 592 190368 604
rect 189684 564 190368 592
rect 189684 552 189690 564
rect 190362 552 190368 564
rect 190420 552 190426 604
rect 281258 552 281264 604
rect 281316 592 281322 604
rect 281442 592 281448 604
rect 281316 564 281448 592
rect 281316 552 281322 564
rect 281442 552 281448 564
rect 281500 552 281506 604
rect 345474 592 345480 604
rect 345435 564 345480 592
rect 345474 552 345480 564
rect 345532 552 345538 604
rect 384666 552 384672 604
rect 384724 592 384730 604
rect 384942 592 384948 604
rect 384724 564 384948 592
rect 384724 552 384730 564
rect 384942 552 384948 564
rect 385000 552 385006 604
rect 392118 552 392124 604
rect 392176 592 392182 604
rect 393038 592 393044 604
rect 392176 564 393044 592
rect 392176 552 392182 564
rect 393038 552 393044 564
rect 393096 552 393102 604
rect 405918 552 405924 604
rect 405976 592 405982 604
rect 406102 592 406108 604
rect 405976 564 406108 592
rect 405976 552 405982 564
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 444837 595 444895 601
rect 444837 561 444849 595
rect 444883 592 444895 595
rect 452470 592 452476 604
rect 444883 564 452476 592
rect 444883 561 444895 564
rect 444837 555 444895 561
rect 452470 552 452476 564
rect 452528 552 452534 604
rect 463694 552 463700 604
rect 463752 592 463758 604
rect 464430 592 464436 604
rect 463752 564 464436 592
rect 463752 552 463758 564
rect 464430 552 464436 564
rect 464488 552 464494 604
rect 471514 592 471520 604
rect 471475 564 471520 592
rect 471514 552 471520 564
rect 471572 552 471578 604
<< via1 >>
rect 202788 700952 202840 701004
rect 358820 700952 358872 701004
rect 170312 700884 170364 700936
rect 362960 700884 363012 700936
rect 328368 700816 328420 700868
rect 527180 700816 527232 700868
rect 329748 700748 329800 700800
rect 543464 700748 543516 700800
rect 154120 700680 154172 700732
rect 367100 700680 367152 700732
rect 137836 700612 137888 700664
rect 364340 700612 364392 700664
rect 105452 700544 105504 700596
rect 368480 700544 368532 700596
rect 89168 700476 89220 700528
rect 374000 700476 374052 700528
rect 72976 700408 73028 700460
rect 371240 700408 371292 700460
rect 40500 700340 40552 700392
rect 375380 700340 375432 700392
rect 24308 700272 24360 700324
rect 379520 700272 379572 700324
rect 218980 700204 219032 700256
rect 360200 700204 360252 700256
rect 336648 700136 336700 700188
rect 478512 700136 478564 700188
rect 335268 700068 335320 700120
rect 462320 700068 462372 700120
rect 235172 700000 235224 700052
rect 356060 700000 356112 700052
rect 267648 699932 267700 699984
rect 351920 699932 351972 699984
rect 283840 699864 283892 699916
rect 354680 699864 354732 699916
rect 343548 699796 343600 699848
rect 413652 699796 413704 699848
rect 340788 699728 340840 699780
rect 397460 699728 397512 699780
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 332508 699660 332560 699712
rect 346400 699660 346452 699712
rect 347780 699660 347832 699712
rect 348792 699660 348844 699712
rect 321468 696940 321520 696992
rect 580172 696940 580224 696992
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 364616 687760 364668 687812
rect 365168 687760 365220 687812
rect 324228 685856 324280 685908
rect 580172 685856 580224 685908
rect 364616 685788 364668 685840
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 382280 681708 382332 681760
rect 364524 676243 364576 676252
rect 364524 676209 364533 676243
rect 364533 676209 364567 676243
rect 364567 676209 364576 676243
rect 364524 676200 364576 676209
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 320088 673480 320140 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 386420 667904 386472 667956
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 383660 652740 383712 652792
rect 315948 650020 316000 650072
rect 580172 650020 580224 650072
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 317328 638936 317380 638988
rect 580172 638936 580224 638988
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 313188 626560 313240 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 387800 623772 387852 623824
rect 364616 618196 364668 618248
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3424 609968 3476 610020
rect 391940 609968 391992 610020
rect 364524 608651 364576 608660
rect 364524 608617 364533 608651
rect 364533 608617 364567 608651
rect 364567 608617 364576 608651
rect 364524 608608 364576 608617
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 309048 603100 309100 603152
rect 580172 603100 580224 603152
rect 429568 601672 429620 601724
rect 559288 601672 559340 601724
rect 364616 598927 364668 598936
rect 364616 598893 364625 598927
rect 364625 598893 364659 598927
rect 364659 598893 364668 598927
rect 364616 598884 364668 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 390560 594804 390612 594856
rect 311808 592016 311860 592068
rect 580172 592016 580224 592068
rect 364708 589296 364760 589348
rect 429660 589296 429712 589348
rect 559380 589296 559432 589348
rect 344468 584672 344520 584724
rect 364708 584672 364760 584724
rect 300768 584604 300820 584656
rect 350816 584604 350868 584656
rect 338212 584536 338264 584588
rect 429660 584536 429712 584588
rect 331864 584468 331916 584520
rect 494244 584468 494296 584520
rect 325516 584400 325568 584452
rect 559380 584400 559432 584452
rect 304540 583652 304592 583704
rect 471428 583652 471480 583704
rect 298192 583584 298244 583636
rect 471336 583584 471388 583636
rect 256056 583516 256108 583568
rect 580632 583516 580684 583568
rect 245568 583448 245620 583500
rect 580448 583448 580500 583500
rect 243452 583380 243504 583432
rect 580264 583380 580316 583432
rect 4712 583312 4764 583364
rect 399208 583312 399260 583364
rect 5448 583244 5500 583296
rect 405556 583244 405608 583296
rect 10324 583176 10376 583228
rect 411904 583176 411956 583228
rect 6276 583108 6328 583160
rect 409788 583108 409840 583160
rect 3148 583040 3200 583092
rect 407672 583040 407724 583092
rect 13084 582972 13136 583024
rect 418160 582972 418212 583024
rect 14464 582904 14516 582956
rect 424508 582904 424560 582956
rect 3240 582836 3292 582888
rect 414020 582836 414072 582888
rect 5356 582768 5408 582820
rect 422392 582768 422444 582820
rect 15844 582700 15896 582752
rect 437112 582700 437164 582752
rect 4068 582632 4120 582684
rect 430856 582632 430908 582684
rect 5264 582564 5316 582616
rect 432972 582564 433024 582616
rect 3884 582496 3936 582548
rect 434996 582496 435048 582548
rect 5172 582428 5224 582480
rect 445576 582428 445628 582480
rect 3700 582360 3752 582412
rect 443460 582360 443512 582412
rect 302424 581612 302476 581664
rect 469588 581612 469640 581664
rect 296076 581544 296128 581596
rect 469680 581544 469732 581596
rect 289728 581476 289780 581528
rect 469772 581476 469824 581528
rect 287612 581408 287664 581460
rect 470508 581408 470560 581460
rect 283472 581340 283524 581392
rect 470416 581340 470468 581392
rect 281356 581272 281408 581324
rect 470324 581272 470376 581324
rect 275008 581204 275060 581256
rect 470232 581204 470284 581256
rect 268660 581136 268712 581188
rect 470048 581136 470100 581188
rect 251824 581068 251876 581120
rect 469864 581068 469916 581120
rect 264520 581000 264572 581052
rect 580080 581000 580132 581052
rect 262404 580252 262456 580304
rect 469956 580252 470008 580304
rect 306564 580184 306616 580236
rect 580172 580184 580224 580236
rect 6644 580116 6696 580168
rect 395068 580116 395120 580168
rect 6552 580048 6604 580100
rect 397092 580048 397144 580100
rect 6460 579980 6512 580032
rect 400956 579980 401008 580032
rect 6368 579912 6420 579964
rect 403164 579912 403216 579964
rect 3792 579844 3844 579896
rect 438860 579844 438912 579896
rect 4988 579776 5040 579828
rect 451556 579776 451608 579828
rect 4896 579708 4948 579760
rect 458272 579708 458324 579760
rect 6184 579640 6236 579692
rect 464252 579640 464304 579692
rect 271144 579368 271196 579420
rect 247960 579343 248012 579352
rect 247960 579309 247969 579343
rect 247969 579309 248003 579343
rect 248003 579309 248012 579343
rect 247960 579300 248012 579309
rect 254216 579343 254268 579352
rect 254216 579309 254225 579343
rect 254225 579309 254259 579343
rect 254259 579309 254268 579343
rect 254216 579300 254268 579309
rect 258448 579300 258500 579352
rect 260656 579300 260708 579352
rect 266912 579300 266964 579352
rect 273168 579300 273220 579352
rect 277308 579300 277360 579352
rect 279608 579300 279660 579352
rect 285772 579300 285824 579352
rect 292120 579343 292172 579352
rect 292120 579309 292129 579343
rect 292129 579309 292163 579343
rect 292163 579309 292172 579343
rect 292120 579300 292172 579309
rect 415676 579343 415728 579352
rect 415676 579309 415685 579343
rect 415685 579309 415719 579343
rect 415719 579309 415728 579343
rect 415676 579300 415728 579309
rect 428372 579343 428424 579352
rect 428372 579309 428381 579343
rect 428381 579309 428415 579343
rect 428415 579309 428424 579343
rect 428372 579300 428424 579309
rect 441068 579343 441120 579352
rect 441068 579309 441077 579343
rect 441077 579309 441111 579343
rect 441111 579309 441120 579343
rect 441068 579300 441120 579309
rect 453580 579343 453632 579352
rect 453580 579309 453589 579343
rect 453589 579309 453623 579343
rect 453623 579309 453632 579343
rect 453580 579300 453632 579309
rect 455788 579343 455840 579352
rect 455788 579309 455797 579343
rect 455797 579309 455831 579343
rect 455831 579309 455840 579343
rect 455788 579300 455840 579309
rect 471244 579232 471296 579284
rect 470140 579164 470192 579216
rect 579804 579096 579856 579148
rect 579988 579028 580040 579080
rect 579896 578960 579948 579012
rect 580080 578892 580132 578944
rect 580908 578824 580960 578876
rect 580724 578756 580776 578808
rect 580816 578688 580868 578740
rect 580540 578620 580592 578672
rect 580356 578552 580408 578604
rect 3332 578484 3384 578536
rect 3976 578416 4028 578468
rect 3608 578348 3660 578400
rect 3424 578280 3476 578332
rect 3516 578212 3568 578264
rect 3056 567332 3108 567384
rect 6644 567332 6696 567384
rect 469588 557472 469640 557524
rect 579712 557472 579764 557524
rect 2780 553052 2832 553104
rect 4712 553052 4764 553104
rect 471428 546388 471480 546440
rect 579712 546388 579764 546440
rect 3056 538636 3108 538688
rect 6552 538636 6604 538688
rect 469680 510552 469732 510604
rect 579712 510552 579764 510604
rect 3056 510212 3108 510264
rect 6460 510212 6512 510264
rect 471336 499468 471388 499520
rect 579712 499468 579764 499520
rect 2780 496680 2832 496732
rect 5448 496680 5500 496732
rect 2964 481108 3016 481160
rect 6368 481108 6420 481160
rect 469772 463632 469824 463684
rect 579712 463632 579764 463684
rect 470508 440172 470560 440224
rect 579804 440172 579856 440224
rect 3148 438812 3200 438864
rect 10324 438812 10376 438864
rect 3148 424056 3200 424108
rect 6276 424056 6328 424108
rect 470416 416712 470468 416764
rect 579804 416712 579856 416764
rect 471244 405628 471296 405680
rect 579804 405628 579856 405680
rect 470324 393252 470376 393304
rect 579804 393252 579856 393304
rect 3240 380808 3292 380860
rect 13084 380808 13136 380860
rect 470232 346332 470284 346384
rect 579988 346332 580040 346384
rect 348516 338648 348568 338700
rect 316132 338104 316184 338156
rect 316316 338104 316368 338156
rect 318800 338104 318852 338156
rect 319812 338104 319864 338156
rect 340328 338104 340380 338156
rect 340696 338104 340748 338156
rect 71044 338036 71096 338088
rect 254952 338036 255004 338088
rect 314660 338036 314712 338088
rect 315396 338036 315448 338088
rect 354404 338036 354456 338088
rect 358084 338036 358136 338088
rect 371516 338036 371568 338088
rect 378876 338036 378928 338088
rect 403348 338036 403400 338088
rect 414664 338036 414716 338088
rect 429844 338036 429896 338088
rect 483020 338036 483072 338088
rect 66904 337968 66956 338020
rect 252008 337968 252060 338020
rect 306196 337968 306248 338020
rect 355876 337968 355928 338020
rect 364248 337968 364300 338020
rect 379336 337968 379388 338020
rect 397460 337968 397512 338020
rect 403624 337968 403676 338020
rect 406292 337968 406344 338020
rect 417424 337968 417476 338020
rect 424968 337968 425020 338020
rect 430120 337968 430172 338020
rect 454776 337968 454828 338020
rect 459744 337968 459796 338020
rect 460848 337968 460900 338020
rect 483388 338036 483440 338088
rect 499580 338036 499632 338088
rect 61384 337900 61436 337952
rect 247592 337900 247644 337952
rect 258724 337900 258776 337952
rect 272616 337900 272668 337952
rect 303160 337900 303212 337952
rect 352932 337900 352984 337952
rect 355324 337900 355376 337952
rect 370044 337900 370096 337952
rect 380348 337900 380400 337952
rect 400404 337900 400456 337952
rect 413284 337900 413336 337952
rect 413652 337900 413704 337952
rect 420276 337900 420328 337952
rect 431316 337900 431368 337952
rect 435732 337900 435784 337952
rect 57244 337832 57296 337884
rect 247132 337832 247184 337884
rect 290464 337832 290516 337884
rect 347044 337832 347096 337884
rect 348424 337832 348476 337884
rect 365628 337832 365680 337884
rect 411720 337832 411772 337884
rect 412548 337832 412600 337884
rect 50344 337764 50396 337816
rect 244188 337764 244240 337816
rect 259644 337764 259696 337816
rect 260104 337764 260156 337816
rect 288256 337764 288308 337816
rect 351920 337764 351972 337816
rect 362868 337764 362920 337816
rect 39304 337696 39356 337748
rect 57980 337696 58032 337748
rect 67548 337696 67600 337748
rect 249064 337696 249116 337748
rect 250536 337696 250588 337748
rect 251456 337696 251508 337748
rect 252468 337696 252520 337748
rect 254584 337696 254636 337748
rect 262312 337696 262364 337748
rect 307760 337696 307812 337748
rect 317328 337696 317380 337748
rect 356704 337696 356756 337748
rect 360752 337696 360804 337748
rect 377404 337764 377456 337816
rect 388444 337764 388496 337816
rect 389180 337764 389232 337816
rect 396080 337764 396132 337816
rect 398196 337764 398248 337816
rect 404360 337764 404412 337816
rect 416136 337764 416188 337816
rect 416688 337764 416740 337816
rect 417608 337832 417660 337884
rect 451832 337900 451884 337952
rect 460664 337832 460716 337884
rect 525064 337968 525116 338020
rect 463608 337900 463660 337952
rect 467104 337900 467156 337952
rect 467748 337900 467800 337952
rect 468024 337900 468076 337952
rect 469128 337900 469180 337952
rect 527824 337900 527876 337952
rect 483020 337832 483072 337884
rect 483388 337832 483440 337884
rect 523684 337832 523736 337884
rect 420184 337764 420236 337816
rect 422024 337764 422076 337816
rect 438676 337764 438728 337816
rect 32404 337628 32456 337680
rect 230664 337628 230716 337680
rect 231124 337628 231176 337680
rect 255964 337628 256016 337680
rect 260104 337628 260156 337680
rect 277032 337628 277084 337680
rect 285588 337628 285640 337680
rect 336096 337628 336148 337680
rect 344560 337628 344612 337680
rect 349988 337628 350040 337680
rect 35164 337560 35216 337612
rect 241704 337560 241756 337612
rect 261392 337560 261444 337612
rect 279976 337560 280028 337612
rect 281448 337560 281500 337612
rect 345572 337560 345624 337612
rect 345756 337560 345808 337612
rect 350172 337560 350224 337612
rect 28264 337492 28316 337544
rect 237840 337492 237892 337544
rect 244648 337492 244700 337544
rect 253204 337492 253256 337544
rect 259368 337492 259420 337544
rect 19984 337424 20036 337476
rect 234344 337424 234396 337476
rect 238300 337424 238352 337476
rect 258816 337424 258868 337476
rect 275560 337492 275612 337544
rect 275928 337492 275980 337544
rect 13084 337356 13136 337408
rect 233516 337356 233568 337408
rect 233884 337356 233936 337408
rect 241244 337356 241296 337408
rect 250444 337356 250496 337408
rect 253480 337356 253532 337408
rect 257344 337356 257396 337408
rect 269672 337424 269724 337476
rect 271788 337424 271840 337476
rect 341616 337492 341668 337544
rect 342720 337492 342772 337544
rect 344376 337492 344428 337544
rect 354864 337628 354916 337680
rect 358728 337628 358780 337680
rect 375932 337696 375984 337748
rect 392584 337696 392636 337748
rect 393228 337696 393280 337748
rect 394056 337696 394108 337748
rect 394608 337696 394660 337748
rect 396540 337696 396592 337748
rect 398104 337696 398156 337748
rect 410248 337696 410300 337748
rect 411168 337696 411220 337748
rect 411260 337696 411312 337748
rect 412364 337696 412416 337748
rect 414204 337696 414256 337748
rect 415308 337696 415360 337748
rect 415584 337696 415636 337748
rect 416504 337696 416556 337748
rect 417056 337696 417108 337748
rect 417976 337696 418028 337748
rect 425428 337696 425480 337748
rect 428464 337696 428516 337748
rect 373908 337628 373960 337680
rect 383292 337628 383344 337680
rect 393596 337628 393648 337680
rect 397460 337628 397512 337680
rect 398012 337628 398064 337680
rect 399484 337628 399536 337680
rect 404820 337628 404872 337680
rect 424324 337628 424376 337680
rect 426440 337628 426492 337680
rect 437480 337696 437532 337748
rect 442356 337696 442408 337748
rect 446036 337764 446088 337816
rect 455696 337764 455748 337816
rect 520924 337764 520976 337816
rect 483020 337696 483072 337748
rect 483388 337696 483440 337748
rect 506480 337696 506532 337748
rect 351184 337560 351236 337612
rect 371148 337560 371200 337612
rect 382280 337560 382332 337612
rect 398932 337560 398984 337612
rect 406384 337560 406436 337612
rect 407304 337560 407356 337612
rect 427084 337560 427136 337612
rect 427912 337560 427964 337612
rect 351828 337492 351880 337544
rect 374460 337492 374512 337544
rect 375288 337492 375340 337544
rect 383752 337492 383804 337544
rect 395068 337492 395120 337544
rect 395896 337492 395948 337544
rect 405832 337492 405884 337544
rect 426440 337492 426492 337544
rect 266728 337356 266780 337408
rect 269028 337356 269080 337408
rect 344100 337424 344152 337476
rect 347504 337424 347556 337476
rect 349068 337424 349120 337476
rect 79324 337288 79376 337340
rect 260840 337288 260892 337340
rect 272800 337288 272852 337340
rect 84844 337220 84896 337272
rect 263784 337220 263836 337272
rect 271328 337220 271380 337272
rect 77944 337152 77996 337204
rect 257896 337152 257948 337204
rect 297916 337152 297968 337204
rect 100668 337084 100720 337136
rect 271144 337084 271196 337136
rect 309784 337288 309836 337340
rect 316040 337288 316092 337340
rect 316868 337288 316920 337340
rect 317420 337288 317472 337340
rect 318340 337288 318392 337340
rect 318892 337288 318944 337340
rect 319260 337288 319312 337340
rect 320180 337288 320232 337340
rect 320732 337288 320784 337340
rect 361764 337288 361816 337340
rect 312544 337220 312596 337272
rect 341800 337220 341852 337272
rect 348976 337220 349028 337272
rect 359464 337220 359516 337272
rect 363696 337220 363748 337272
rect 372068 337424 372120 337476
rect 381820 337424 381872 337476
rect 397000 337424 397052 337476
rect 405924 337424 405976 337476
rect 420552 337424 420604 337476
rect 436652 337560 436704 337612
rect 437388 337560 437440 337612
rect 432788 337424 432840 337476
rect 437204 337424 437256 337476
rect 437480 337424 437532 337476
rect 439596 337492 439648 337544
rect 442264 337424 442316 337476
rect 455604 337628 455656 337680
rect 457720 337628 457772 337680
rect 521016 337628 521068 337680
rect 443092 337560 443144 337612
rect 448980 337560 449032 337612
rect 483020 337560 483072 337612
rect 483480 337560 483532 337612
rect 518164 337560 518216 337612
rect 463608 337492 463660 337544
rect 483112 337492 483164 337544
rect 483296 337492 483348 337544
rect 514024 337492 514076 337544
rect 449164 337424 449216 337476
rect 516784 337424 516836 337476
rect 369768 337356 369820 337408
rect 400956 337356 401008 337408
rect 402244 337356 402296 337408
rect 367008 337288 367060 337340
rect 380808 337288 380860 337340
rect 398472 337288 398524 337340
rect 408776 337356 408828 337408
rect 409144 337356 409196 337408
rect 372988 337220 373040 337272
rect 412732 337356 412784 337408
rect 413836 337356 413888 337408
rect 421196 337356 421248 337408
rect 438124 337356 438176 337408
rect 440148 337356 440200 337408
rect 510620 337356 510672 337408
rect 421012 337288 421064 337340
rect 423496 337220 423548 337272
rect 459192 337220 459244 337272
rect 460296 337220 460348 337272
rect 464620 337288 464672 337340
rect 466552 337288 466604 337340
rect 529204 337288 529256 337340
rect 469496 337220 469548 337272
rect 530584 337220 530636 337272
rect 314200 337152 314252 337204
rect 321468 337152 321520 337204
rect 312728 337084 312780 337136
rect 316684 337084 316736 337136
rect 342904 337152 342956 337204
rect 355968 337152 356020 337204
rect 335268 337084 335320 337136
rect 95884 337016 95936 337068
rect 265256 337016 265308 337068
rect 366640 337084 366692 337136
rect 369124 337084 369176 337136
rect 371056 337084 371108 337136
rect 367652 337016 367704 337068
rect 107568 336948 107620 337000
rect 274088 336948 274140 337000
rect 319444 336948 319496 337000
rect 102784 336880 102836 336932
rect 268200 336880 268252 336932
rect 333244 336880 333296 336932
rect 338764 336880 338816 336932
rect 118608 336812 118660 336864
rect 278504 336812 278556 336864
rect 327724 336812 327776 336864
rect 340788 336880 340840 336932
rect 125508 336744 125560 336796
rect 281172 336744 281224 336796
rect 340236 336744 340288 336796
rect 251824 336676 251876 336728
rect 256424 336676 256476 336728
rect 262864 336676 262916 336728
rect 263048 336676 263100 336728
rect 284392 336719 284444 336728
rect 284392 336685 284401 336719
rect 284401 336685 284435 336719
rect 284435 336685 284444 336719
rect 284392 336676 284444 336685
rect 288992 336676 289044 336728
rect 327632 336676 327684 336728
rect 340328 336676 340380 336728
rect 343088 336744 343140 336796
rect 344284 336812 344336 336864
rect 345572 336744 345624 336796
rect 353392 336948 353444 337000
rect 345940 336880 345992 336932
rect 360292 336880 360344 336932
rect 366916 336948 366968 337000
rect 378048 336948 378100 337000
rect 385224 337152 385276 337204
rect 401876 337152 401928 337204
rect 416964 337152 417016 337204
rect 380808 337084 380860 337136
rect 386236 337084 386288 337136
rect 415124 337084 415176 337136
rect 421564 337084 421616 337136
rect 407764 337016 407816 337068
rect 409144 337016 409196 337068
rect 419080 337016 419132 337068
rect 431224 337152 431276 337204
rect 433524 337152 433576 337204
rect 434260 337152 434312 337204
rect 492680 337152 492732 337204
rect 433984 337084 434036 337136
rect 485780 337084 485832 337136
rect 422484 337016 422536 337068
rect 424416 337016 424468 337068
rect 382188 336948 382240 337000
rect 386696 336948 386748 337000
rect 401416 336948 401468 337000
rect 405004 336948 405056 337000
rect 409236 336948 409288 337000
rect 369584 336880 369636 336932
rect 384304 336880 384356 336932
rect 387708 336880 387760 336932
rect 357348 336812 357400 336864
rect 362224 336812 362276 336864
rect 365168 336812 365220 336864
rect 381636 336812 381688 336864
rect 384764 336812 384816 336864
rect 384948 336812 385000 336864
rect 388168 336812 388220 336864
rect 420000 336812 420052 336864
rect 420736 336812 420788 336864
rect 351460 336744 351512 336796
rect 352564 336744 352616 336796
rect 357808 336744 357860 336796
rect 363604 336744 363656 336796
rect 364708 336744 364760 336796
rect 370504 336744 370556 336796
rect 372528 336744 372580 336796
rect 376024 336744 376076 336796
rect 376944 336744 376996 336796
rect 377680 336744 377732 336796
rect 378416 336744 378468 336796
rect 380164 336744 380216 336796
rect 381360 336744 381412 336796
rect 381544 336744 381596 336796
rect 382832 336744 382884 336796
rect 387064 336744 387116 336796
rect 388720 336744 388772 336796
rect 392400 336744 392452 336796
rect 393596 336744 393648 336796
rect 418528 336744 418580 336796
rect 419448 336744 419500 336796
rect 419540 336744 419592 336796
rect 420828 336744 420880 336796
rect 421472 336744 421524 336796
rect 422208 336744 422260 336796
rect 428372 336948 428424 337000
rect 431316 336948 431368 337000
rect 423956 336880 424008 336932
rect 426900 336812 426952 336864
rect 477592 337016 477644 337068
rect 475384 336948 475436 337000
rect 469220 336880 469272 336932
rect 434720 336812 434772 336864
rect 436008 336812 436060 336864
rect 429384 336744 429436 336796
rect 430488 336744 430540 336796
rect 430856 336744 430908 336796
rect 431868 336744 431920 336796
rect 432328 336744 432380 336796
rect 433156 336744 433208 336796
rect 433708 336744 433760 336796
rect 434628 336744 434680 336796
rect 435180 336744 435232 336796
rect 435916 336744 435968 336796
rect 436192 336744 436244 336796
rect 437296 336744 437348 336796
rect 439504 336812 439556 336864
rect 441620 336812 441672 336864
rect 443644 336812 443696 336864
rect 444564 336812 444616 336864
rect 445668 336812 445720 336864
rect 450452 336812 450504 336864
rect 451188 336812 451240 336864
rect 453304 336812 453356 336864
rect 453948 336812 454000 336864
rect 456800 336812 456852 336864
rect 458088 336812 458140 336864
rect 439136 336744 439188 336796
rect 440148 336744 440200 336796
rect 440608 336744 440660 336796
rect 441528 336744 441580 336796
rect 442080 336744 442132 336796
rect 442908 336744 442960 336796
rect 443552 336744 443604 336796
rect 444288 336744 444340 336796
rect 445024 336744 445076 336796
rect 445576 336744 445628 336796
rect 446496 336744 446548 336796
rect 447048 336744 447100 336796
rect 447508 336744 447560 336796
rect 421196 336719 421248 336728
rect 421196 336685 421205 336719
rect 421205 336685 421239 336719
rect 421239 336685 421248 336719
rect 421196 336676 421248 336685
rect 448244 336744 448296 336796
rect 448428 336744 448480 336796
rect 449900 336744 449952 336796
rect 451004 336744 451056 336796
rect 451372 336744 451424 336796
rect 452476 336744 452528 336796
rect 452844 336744 452896 336796
rect 453764 336744 453816 336796
rect 454316 336744 454368 336796
rect 455236 336744 455288 336796
rect 455788 336744 455840 336796
rect 456616 336744 456668 336796
rect 457260 336744 457312 336796
rect 457996 336744 458048 336796
rect 459652 336812 459704 336864
rect 458272 336744 458324 336796
rect 459468 336744 459520 336796
rect 463792 336812 463844 336864
rect 461216 336744 461268 336796
rect 462136 336744 462188 336796
rect 462688 336744 462740 336796
rect 463516 336744 463568 336796
rect 464160 336744 464212 336796
rect 464988 336744 465040 336796
rect 461952 336676 462004 336728
rect 448428 336608 448480 336660
rect 470600 336812 470652 336864
rect 509884 336812 509936 336864
rect 505744 336744 505796 336796
rect 247684 336472 247736 336524
rect 248604 336472 248656 336524
rect 248512 336064 248564 336116
rect 249524 336064 249576 336116
rect 236184 335656 236236 335708
rect 237012 335656 237064 335708
rect 302240 335656 302292 335708
rect 302700 335656 302752 335708
rect 332692 335656 332744 335708
rect 333428 335656 333480 335708
rect 334072 335656 334124 335708
rect 334900 335656 334952 335708
rect 236092 335588 236144 335640
rect 236552 335588 236604 335640
rect 241612 335588 241664 335640
rect 242348 335588 242400 335640
rect 260932 335588 260984 335640
rect 261484 335588 261536 335640
rect 263692 335588 263744 335640
rect 264428 335588 264480 335640
rect 265072 335588 265124 335640
rect 265900 335588 265952 335640
rect 266452 335588 266504 335640
rect 267372 335588 267424 335640
rect 280252 335588 280304 335640
rect 280620 335588 280672 335640
rect 281540 335588 281592 335640
rect 282092 335588 282144 335640
rect 283012 335588 283064 335640
rect 283564 335588 283616 335640
rect 285680 335588 285732 335640
rect 285956 335588 286008 335640
rect 286048 335588 286100 335640
rect 286600 335588 286652 335640
rect 287060 335588 287112 335640
rect 287980 335588 288032 335640
rect 288440 335588 288492 335640
rect 289452 335588 289504 335640
rect 292764 335588 292816 335640
rect 293316 335588 293368 335640
rect 298284 335588 298336 335640
rect 298652 335588 298704 335640
rect 300860 335588 300912 335640
rect 301228 335588 301280 335640
rect 303620 335588 303672 335640
rect 304172 335588 304224 335640
rect 305000 335588 305052 335640
rect 305644 335588 305696 335640
rect 307760 335588 307812 335640
rect 308588 335588 308640 335640
rect 309140 335588 309192 335640
rect 310060 335588 310112 335640
rect 321652 335588 321704 335640
rect 322204 335588 322256 335640
rect 329840 335588 329892 335640
rect 330116 335588 330168 335640
rect 332600 335588 332652 335640
rect 333060 335588 333112 335640
rect 333980 335588 334032 335640
rect 334532 335588 334584 335640
rect 335360 335588 335412 335640
rect 336004 335588 336056 335640
rect 338120 335588 338172 335640
rect 338948 335588 339000 335640
rect 363052 335588 363104 335640
rect 363788 335588 363840 335640
rect 367284 335588 367336 335640
rect 367928 335588 367980 335640
rect 374092 335588 374144 335640
rect 374644 335588 374696 335640
rect 465448 335588 465500 335640
rect 466368 335588 466420 335640
rect 245844 335452 245896 335504
rect 246672 335452 246724 335504
rect 438032 335452 438084 335504
rect 438676 335452 438728 335504
rect 284484 335180 284536 335232
rect 258172 334704 258224 334756
rect 258540 334704 258592 334756
rect 303068 334704 303120 334756
rect 234988 334500 235040 334552
rect 235632 334500 235684 334552
rect 250628 334432 250680 334484
rect 270776 334296 270828 334348
rect 271236 334296 271288 334348
rect 272248 334296 272300 334348
rect 272708 334296 272760 334348
rect 247132 334160 247184 334212
rect 248144 334160 248196 334212
rect 278780 333276 278832 333328
rect 278964 333276 279016 333328
rect 325976 333276 326028 333328
rect 326528 333276 326580 333328
rect 336740 333276 336792 333328
rect 336924 333276 336976 333328
rect 361672 333276 361724 333328
rect 362316 333276 362368 333328
rect 356152 332800 356204 332852
rect 356612 332800 356664 332852
rect 284668 332528 284720 332580
rect 285128 332528 285180 332580
rect 331220 332120 331272 332172
rect 331496 332120 331548 332172
rect 242992 332052 243044 332104
rect 243452 332052 243504 332104
rect 310520 332052 310572 332104
rect 311532 332052 311584 332104
rect 301044 331848 301096 331900
rect 301688 331848 301740 331900
rect 331312 331712 331364 331764
rect 331956 331712 332008 331764
rect 328552 331304 328604 331356
rect 329012 331304 329064 331356
rect 299572 331236 299624 331288
rect 336832 331236 336884 331288
rect 259644 331168 259696 331220
rect 259828 331168 259880 331220
rect 341156 331168 341208 331220
rect 341340 331168 341392 331220
rect 360292 331168 360344 331220
rect 360476 331168 360528 331220
rect 459652 331168 459704 331220
rect 460112 331168 460164 331220
rect 299572 331100 299624 331152
rect 299756 331100 299808 331152
rect 300216 331100 300268 331152
rect 336832 331100 336884 331152
rect 299480 331032 299532 331084
rect 299664 331032 299716 331084
rect 306472 331032 306524 331084
rect 306656 331032 306708 331084
rect 284300 329536 284352 329588
rect 284576 329536 284628 329588
rect 250168 328491 250220 328500
rect 250168 328457 250177 328491
rect 250177 328457 250211 328491
rect 250211 328457 250220 328491
rect 250168 328448 250220 328457
rect 278872 328448 278924 328500
rect 279056 328448 279108 328500
rect 302516 328491 302568 328500
rect 302516 328457 302525 328491
rect 302525 328457 302559 328491
rect 302559 328457 302568 328491
rect 302516 328448 302568 328457
rect 303896 328448 303948 328500
rect 304632 328448 304684 328500
rect 323308 328448 323360 328500
rect 323676 328448 323728 328500
rect 324688 328448 324740 328500
rect 325148 328448 325200 328500
rect 337292 328448 337344 328500
rect 337384 328448 337436 328500
rect 372712 328448 372764 328500
rect 373264 328448 373316 328500
rect 375656 328448 375708 328500
rect 376116 328448 376168 328500
rect 259828 328423 259880 328432
rect 259828 328389 259837 328423
rect 259837 328389 259871 328423
rect 259871 328389 259880 328423
rect 259828 328380 259880 328389
rect 295524 328380 295576 328432
rect 295708 328380 295760 328432
rect 296812 328380 296864 328432
rect 296996 328380 297048 328432
rect 341340 328423 341392 328432
rect 341340 328389 341349 328423
rect 341349 328389 341383 328423
rect 341383 328389 341392 328423
rect 341340 328380 341392 328389
rect 358728 328423 358780 328432
rect 358728 328389 358737 328423
rect 358737 328389 358771 328423
rect 358771 328389 358780 328423
rect 358728 328380 358780 328389
rect 470600 328423 470652 328432
rect 470600 328389 470609 328423
rect 470609 328389 470643 328423
rect 470643 328389 470652 328423
rect 470600 328380 470652 328389
rect 330484 327156 330536 327208
rect 327264 327131 327316 327140
rect 327264 327097 327273 327131
rect 327273 327097 327307 327131
rect 327307 327097 327316 327131
rect 327264 327088 327316 327097
rect 330116 327088 330168 327140
rect 421196 327131 421248 327140
rect 421196 327097 421205 327131
rect 421205 327097 421239 327131
rect 421239 327097 421248 327131
rect 421196 327088 421248 327097
rect 299848 327063 299900 327072
rect 299848 327029 299857 327063
rect 299857 327029 299891 327063
rect 299891 327029 299900 327063
rect 299848 327020 299900 327029
rect 301136 327020 301188 327072
rect 301320 327020 301372 327072
rect 359188 327063 359240 327072
rect 359188 327029 359197 327063
rect 359197 327029 359231 327063
rect 359231 327029 359240 327063
rect 359188 327020 359240 327029
rect 272156 324300 272208 324352
rect 272248 324300 272300 324352
rect 3332 324232 3384 324284
rect 14464 324232 14516 324284
rect 470140 322872 470192 322924
rect 579988 322872 580040 322924
rect 262772 322260 262824 322312
rect 251456 321580 251508 321632
rect 266728 321580 266780 321632
rect 267832 321580 267884 321632
rect 310796 321580 310848 321632
rect 337292 321580 337344 321632
rect 377128 321580 377180 321632
rect 232228 321512 232280 321564
rect 232412 321512 232464 321564
rect 310888 321444 310940 321496
rect 337384 321444 337436 321496
rect 251548 321376 251600 321428
rect 377220 321376 377272 321428
rect 288808 319107 288860 319116
rect 288808 319073 288817 319107
rect 288817 319073 288851 319107
rect 288851 319073 288860 319107
rect 288808 319064 288860 319073
rect 265256 318903 265308 318912
rect 265256 318869 265265 318903
rect 265265 318869 265299 318903
rect 265299 318869 265308 318903
rect 265256 318860 265308 318869
rect 259920 318792 259972 318844
rect 266636 318835 266688 318844
rect 266636 318801 266645 318835
rect 266645 318801 266679 318835
rect 266679 318801 266688 318835
rect 266636 318792 266688 318801
rect 267740 318835 267792 318844
rect 267740 318801 267749 318835
rect 267749 318801 267783 318835
rect 267783 318801 267792 318835
rect 267740 318792 267792 318801
rect 284668 318792 284720 318844
rect 284760 318792 284812 318844
rect 302516 318792 302568 318844
rect 302608 318792 302660 318844
rect 306748 318792 306800 318844
rect 306840 318792 306892 318844
rect 330116 318792 330168 318844
rect 339776 318835 339828 318844
rect 339776 318801 339785 318835
rect 339785 318801 339819 318835
rect 339819 318801 339828 318835
rect 339776 318792 339828 318801
rect 341432 318792 341484 318844
rect 358728 318835 358780 318844
rect 358728 318801 358737 318835
rect 358737 318801 358771 318835
rect 358771 318801 358780 318835
rect 358728 318792 358780 318801
rect 470600 318835 470652 318844
rect 470600 318801 470609 318835
rect 470609 318801 470643 318835
rect 470643 318801 470652 318835
rect 470600 318792 470652 318801
rect 372712 318767 372764 318776
rect 372712 318733 372721 318767
rect 372721 318733 372755 318767
rect 372755 318733 372764 318767
rect 372712 318724 372764 318733
rect 330208 318656 330260 318708
rect 359188 317747 359240 317756
rect 359188 317713 359197 317747
rect 359197 317713 359231 317747
rect 359231 317713 359240 317747
rect 359188 317704 359240 317713
rect 262680 317475 262732 317484
rect 262680 317441 262689 317475
rect 262689 317441 262723 317475
rect 262723 317441 262732 317475
rect 262680 317432 262732 317441
rect 265256 317475 265308 317484
rect 265256 317441 265265 317475
rect 265265 317441 265299 317475
rect 265299 317441 265308 317475
rect 265256 317432 265308 317441
rect 299848 317475 299900 317484
rect 299848 317441 299857 317475
rect 299857 317441 299891 317475
rect 299891 317441 299900 317475
rect 299848 317432 299900 317441
rect 358728 317407 358780 317416
rect 358728 317373 358737 317407
rect 358737 317373 358771 317407
rect 358771 317373 358780 317407
rect 358728 317364 358780 317373
rect 421196 317407 421248 317416
rect 421196 317373 421205 317407
rect 421205 317373 421239 317407
rect 421239 317373 421248 317407
rect 421196 317364 421248 317373
rect 460204 317407 460256 317416
rect 460204 317373 460213 317407
rect 460213 317373 460247 317407
rect 460247 317373 460256 317407
rect 460204 317364 460256 317373
rect 386788 316072 386840 316124
rect 386972 316072 387024 316124
rect 270500 316004 270552 316056
rect 270684 316004 270736 316056
rect 273536 316004 273588 316056
rect 273628 316004 273680 316056
rect 294144 316004 294196 316056
rect 294236 316004 294288 316056
rect 262680 315979 262732 315988
rect 262680 315945 262689 315979
rect 262689 315945 262723 315979
rect 262723 315945 262732 315979
rect 262680 315936 262732 315945
rect 386788 315979 386840 315988
rect 386788 315945 386797 315979
rect 386797 315945 386831 315979
rect 386831 315945 386840 315979
rect 386788 315936 386840 315945
rect 272156 314619 272208 314628
rect 272156 314585 272165 314619
rect 272165 314585 272199 314619
rect 272199 314585 272208 314619
rect 272156 314576 272208 314585
rect 250168 313964 250220 314016
rect 250168 313828 250220 313880
rect 232412 311924 232464 311976
rect 288808 311924 288860 311976
rect 310888 311967 310940 311976
rect 310888 311933 310897 311967
rect 310897 311933 310931 311967
rect 310931 311933 310940 311967
rect 310888 311924 310940 311933
rect 323308 311924 323360 311976
rect 259736 311856 259788 311908
rect 259920 311856 259972 311908
rect 284668 311856 284720 311908
rect 285956 311899 286008 311908
rect 285956 311865 285965 311899
rect 285965 311865 285999 311899
rect 285999 311865 286008 311899
rect 285956 311856 286008 311865
rect 323216 311856 323268 311908
rect 337200 311856 337252 311908
rect 337384 311856 337436 311908
rect 341248 311856 341300 311908
rect 341432 311856 341484 311908
rect 232320 311788 232372 311840
rect 244464 311831 244516 311840
rect 244464 311797 244473 311831
rect 244473 311797 244507 311831
rect 244507 311797 244516 311831
rect 244464 311788 244516 311797
rect 339684 311788 339736 311840
rect 339868 311788 339920 311840
rect 273444 309315 273496 309324
rect 273444 309281 273453 309315
rect 273453 309281 273487 309315
rect 273487 309281 273496 309315
rect 273444 309272 273496 309281
rect 266636 309204 266688 309256
rect 244464 309179 244516 309188
rect 244464 309145 244473 309179
rect 244473 309145 244507 309179
rect 244507 309145 244516 309179
rect 244464 309136 244516 309145
rect 290004 309136 290056 309188
rect 290096 309136 290148 309188
rect 372712 309179 372764 309188
rect 372712 309145 372721 309179
rect 372721 309145 372755 309179
rect 372755 309145 372764 309179
rect 372712 309136 372764 309145
rect 236276 309111 236328 309120
rect 236276 309077 236285 309111
rect 236285 309077 236319 309111
rect 236319 309077 236328 309111
rect 236276 309068 236328 309077
rect 259736 309068 259788 309120
rect 265256 309111 265308 309120
rect 265256 309077 265265 309111
rect 265265 309077 265299 309111
rect 265299 309077 265308 309111
rect 265256 309068 265308 309077
rect 266636 309068 266688 309120
rect 339868 309111 339920 309120
rect 339868 309077 339877 309111
rect 339877 309077 339911 309111
rect 339911 309077 339920 309111
rect 339868 309068 339920 309077
rect 341248 309068 341300 309120
rect 470600 309111 470652 309120
rect 470600 309077 470609 309111
rect 470609 309077 470643 309111
rect 470643 309077 470652 309111
rect 470600 309068 470652 309077
rect 327264 309000 327316 309052
rect 327356 309000 327408 309052
rect 2780 308796 2832 308848
rect 5356 308796 5408 308848
rect 310704 307844 310756 307896
rect 301044 307776 301096 307828
rect 301228 307776 301280 307828
rect 358728 307819 358780 307828
rect 358728 307785 358737 307819
rect 358737 307785 358771 307819
rect 358771 307785 358780 307819
rect 358728 307776 358780 307785
rect 421196 307819 421248 307828
rect 421196 307785 421205 307819
rect 421205 307785 421239 307819
rect 421239 307785 421248 307819
rect 421196 307776 421248 307785
rect 460204 307819 460256 307828
rect 460204 307785 460213 307819
rect 460213 307785 460247 307819
rect 460247 307785 460256 307819
rect 460204 307776 460256 307785
rect 310704 307751 310756 307760
rect 310704 307717 310713 307751
rect 310713 307717 310747 307751
rect 310747 307717 310756 307751
rect 310704 307708 310756 307717
rect 325608 307708 325660 307760
rect 325976 307708 326028 307760
rect 337200 307708 337252 307760
rect 285772 306416 285824 306468
rect 262680 306391 262732 306400
rect 262680 306357 262689 306391
rect 262689 306357 262723 306391
rect 262723 306357 262732 306391
rect 284576 306391 284628 306400
rect 262680 306348 262732 306357
rect 284576 306357 284585 306391
rect 284585 306357 284619 306391
rect 284619 306357 284628 306391
rect 284576 306348 284628 306357
rect 317512 306348 317564 306400
rect 317696 306348 317748 306400
rect 463700 306348 463752 306400
rect 463884 306348 463936 306400
rect 357808 302268 357860 302320
rect 295616 302132 295668 302184
rect 327356 302132 327408 302184
rect 295708 302064 295760 302116
rect 357900 302064 357952 302116
rect 386788 302107 386840 302116
rect 386788 302073 386797 302107
rect 386797 302073 386831 302107
rect 386831 302073 386840 302107
rect 386788 302064 386840 302073
rect 273536 301520 273588 301572
rect 339868 299931 339920 299940
rect 339868 299897 339877 299931
rect 339877 299897 339911 299931
rect 339911 299897 339920 299931
rect 339868 299888 339920 299897
rect 259644 299591 259696 299600
rect 259644 299557 259653 299591
rect 259653 299557 259687 299591
rect 259687 299557 259696 299591
rect 259644 299548 259696 299557
rect 236460 299480 236512 299532
rect 239128 299480 239180 299532
rect 239312 299480 239364 299532
rect 262588 299480 262640 299532
rect 265256 299523 265308 299532
rect 265256 299489 265265 299523
rect 265265 299489 265299 299523
rect 265299 299489 265308 299523
rect 265256 299480 265308 299489
rect 267832 299548 267884 299600
rect 341156 299523 341208 299532
rect 341156 299489 341165 299523
rect 341165 299489 341199 299523
rect 341199 299489 341208 299523
rect 341156 299480 341208 299489
rect 359280 299548 359332 299600
rect 470600 299523 470652 299532
rect 470600 299489 470609 299523
rect 470609 299489 470643 299523
rect 470643 299489 470652 299523
rect 470600 299480 470652 299489
rect 259644 299412 259696 299464
rect 259828 299412 259880 299464
rect 262680 299412 262732 299464
rect 267740 299412 267792 299464
rect 323308 299455 323360 299464
rect 323308 299421 323317 299455
rect 323317 299421 323351 299455
rect 323351 299421 323360 299455
rect 323308 299412 323360 299421
rect 324688 299455 324740 299464
rect 324688 299421 324697 299455
rect 324697 299421 324731 299455
rect 324731 299421 324740 299455
rect 324688 299412 324740 299421
rect 359096 299412 359148 299464
rect 372712 299455 372764 299464
rect 372712 299421 372721 299455
rect 372721 299421 372755 299455
rect 372755 299421 372764 299455
rect 372712 299412 372764 299421
rect 375748 299412 375800 299464
rect 470048 299412 470100 299464
rect 579804 299412 579856 299464
rect 337016 298231 337068 298240
rect 337016 298197 337025 298231
rect 337025 298197 337059 298231
rect 337059 298197 337068 298231
rect 337016 298188 337068 298197
rect 266636 298163 266688 298172
rect 266636 298129 266645 298163
rect 266645 298129 266679 298163
rect 266679 298129 266688 298163
rect 266636 298120 266688 298129
rect 310888 298120 310940 298172
rect 327264 298163 327316 298172
rect 327264 298129 327273 298163
rect 327273 298129 327307 298163
rect 327307 298129 327316 298163
rect 327264 298120 327316 298129
rect 337016 298052 337068 298104
rect 358728 298095 358780 298104
rect 358728 298061 358737 298095
rect 358737 298061 358771 298095
rect 358771 298061 358780 298095
rect 358728 298052 358780 298061
rect 359096 298095 359148 298104
rect 359096 298061 359105 298095
rect 359105 298061 359139 298095
rect 359139 298061 359148 298095
rect 359096 298052 359148 298061
rect 421196 298095 421248 298104
rect 421196 298061 421205 298095
rect 421205 298061 421239 298095
rect 421239 298061 421248 298095
rect 421196 298052 421248 298061
rect 460020 298095 460072 298104
rect 460020 298061 460029 298095
rect 460029 298061 460063 298095
rect 460063 298061 460072 298095
rect 460020 298052 460072 298061
rect 329932 297712 329984 297764
rect 330392 297712 330444 297764
rect 266636 296735 266688 296744
rect 266636 296701 266645 296735
rect 266645 296701 266679 296735
rect 266679 296701 266688 296735
rect 266636 296692 266688 296701
rect 270776 296692 270828 296744
rect 270960 296692 271012 296744
rect 272248 296692 272300 296744
rect 285772 296692 285824 296744
rect 286048 296692 286100 296744
rect 294144 296692 294196 296744
rect 294328 296692 294380 296744
rect 270776 295264 270828 295316
rect 270960 295264 271012 295316
rect 272248 295264 272300 295316
rect 251548 294652 251600 294704
rect 290004 294584 290056 294636
rect 290188 294584 290240 294636
rect 306748 294584 306800 294636
rect 306932 294584 306984 294636
rect 310888 293063 310940 293072
rect 310888 293029 310897 293063
rect 310897 293029 310931 293063
rect 310931 293029 310940 293063
rect 310888 293020 310940 293029
rect 386788 293063 386840 293072
rect 386788 293029 386797 293063
rect 386797 293029 386831 293063
rect 386831 293029 386840 293063
rect 386788 293020 386840 293029
rect 236276 292544 236328 292596
rect 236460 292544 236512 292596
rect 296812 292544 296864 292596
rect 301044 292544 301096 292596
rect 357440 292544 357492 292596
rect 357900 292544 357952 292596
rect 239036 292476 239088 292528
rect 239220 292476 239272 292528
rect 296904 292476 296956 292528
rect 301136 292476 301188 292528
rect 337200 292451 337252 292460
rect 337200 292417 337209 292451
rect 337209 292417 337243 292451
rect 337243 292417 337252 292451
rect 337200 292408 337252 292417
rect 285772 291864 285824 291916
rect 286048 291864 286100 291916
rect 288716 290003 288768 290012
rect 288716 289969 288725 290003
rect 288725 289969 288759 290003
rect 288759 289969 288768 290003
rect 288716 289960 288768 289969
rect 251456 289867 251508 289876
rect 251456 289833 251465 289867
rect 251465 289833 251499 289867
rect 251499 289833 251508 289867
rect 251456 289824 251508 289833
rect 299756 289824 299808 289876
rect 299848 289824 299900 289876
rect 324688 289867 324740 289876
rect 324688 289833 324697 289867
rect 324697 289833 324731 289867
rect 324731 289833 324740 289867
rect 324688 289824 324740 289833
rect 372712 289867 372764 289876
rect 372712 289833 372721 289867
rect 372721 289833 372755 289867
rect 372755 289833 372764 289867
rect 372712 289824 372764 289833
rect 375656 289867 375708 289876
rect 375656 289833 375665 289867
rect 375665 289833 375699 289867
rect 375699 289833 375708 289867
rect 375656 289824 375708 289833
rect 377128 289824 377180 289876
rect 377220 289824 377272 289876
rect 250076 289756 250128 289808
rect 250352 289756 250404 289808
rect 259736 289756 259788 289808
rect 259920 289756 259972 289808
rect 284576 289756 284628 289808
rect 288716 289756 288768 289808
rect 288808 289756 288860 289808
rect 290004 289756 290056 289808
rect 290188 289756 290240 289808
rect 302516 289756 302568 289808
rect 302700 289756 302752 289808
rect 306748 289756 306800 289808
rect 306932 289756 306984 289808
rect 327264 289756 327316 289808
rect 341248 289756 341300 289808
rect 470600 289799 470652 289808
rect 470600 289765 470609 289799
rect 470609 289765 470643 289799
rect 470643 289765 470652 289799
rect 470600 289756 470652 289765
rect 284760 289688 284812 289740
rect 327356 289688 327408 289740
rect 295708 288464 295760 288516
rect 323492 288464 323544 288516
rect 267740 288396 267792 288448
rect 267832 288396 267884 288448
rect 359188 288396 359240 288448
rect 421196 288439 421248 288448
rect 421196 288405 421205 288439
rect 421205 288405 421239 288439
rect 421239 288405 421248 288439
rect 421196 288396 421248 288405
rect 460112 288396 460164 288448
rect 325884 288328 325936 288380
rect 326068 288328 326120 288380
rect 329932 288328 329984 288380
rect 330300 288328 330352 288380
rect 266636 287036 266688 287088
rect 266728 287036 266780 287088
rect 291568 287036 291620 287088
rect 291752 287036 291804 287088
rect 294236 287036 294288 287088
rect 294328 287036 294380 287088
rect 295524 287079 295576 287088
rect 295524 287045 295533 287079
rect 295533 287045 295567 287079
rect 295567 287045 295576 287079
rect 295524 287036 295576 287045
rect 296904 286968 296956 287020
rect 272156 285719 272208 285728
rect 272156 285685 272165 285719
rect 272165 285685 272199 285719
rect 272199 285685 272208 285719
rect 272156 285676 272208 285685
rect 266728 285651 266780 285660
rect 266728 285617 266737 285651
rect 266737 285617 266771 285651
rect 266771 285617 266780 285651
rect 266728 285608 266780 285617
rect 236276 282888 236328 282940
rect 301136 282956 301188 283008
rect 460112 282956 460164 283008
rect 337108 282931 337160 282940
rect 337108 282897 337117 282931
rect 337117 282897 337151 282931
rect 337151 282897 337160 282931
rect 337108 282888 337160 282897
rect 339684 282888 339736 282940
rect 339868 282888 339920 282940
rect 357440 282888 357492 282940
rect 301044 282820 301096 282872
rect 360292 282888 360344 282940
rect 360476 282888 360528 282940
rect 236460 282752 236512 282804
rect 310888 282795 310940 282804
rect 310888 282761 310897 282795
rect 310897 282761 310931 282795
rect 310931 282761 310940 282795
rect 310888 282752 310940 282761
rect 357716 282752 357768 282804
rect 386788 282795 386840 282804
rect 386788 282761 386797 282795
rect 386797 282761 386831 282795
rect 386831 282761 386840 282795
rect 386788 282752 386840 282761
rect 460112 282752 460164 282804
rect 270776 282208 270828 282260
rect 270960 282208 271012 282260
rect 295524 280780 295576 280832
rect 295800 280780 295852 280832
rect 358728 280279 358780 280288
rect 358728 280245 358737 280279
rect 358737 280245 358771 280279
rect 358771 280245 358780 280279
rect 358728 280236 358780 280245
rect 325884 280211 325936 280220
rect 325884 280177 325893 280211
rect 325893 280177 325927 280211
rect 325927 280177 325936 280211
rect 325884 280168 325936 280177
rect 341156 280211 341208 280220
rect 341156 280177 341165 280211
rect 341165 280177 341199 280211
rect 341199 280177 341208 280211
rect 341156 280168 341208 280177
rect 470600 280211 470652 280220
rect 470600 280177 470609 280211
rect 470609 280177 470643 280211
rect 470643 280177 470652 280211
rect 470600 280168 470652 280177
rect 236460 280100 236512 280152
rect 239128 280143 239180 280152
rect 239128 280109 239137 280143
rect 239137 280109 239171 280143
rect 239171 280109 239180 280143
rect 239128 280100 239180 280109
rect 251456 280143 251508 280152
rect 251456 280109 251465 280143
rect 251465 280109 251499 280143
rect 251499 280109 251508 280143
rect 251456 280100 251508 280109
rect 259552 280143 259604 280152
rect 259552 280109 259561 280143
rect 259561 280109 259595 280143
rect 259595 280109 259604 280143
rect 259552 280100 259604 280109
rect 273536 280100 273588 280152
rect 273628 280100 273680 280152
rect 284576 280100 284628 280152
rect 284760 280100 284812 280152
rect 336924 280143 336976 280152
rect 336924 280109 336933 280143
rect 336933 280109 336967 280143
rect 336967 280109 336976 280143
rect 336924 280100 336976 280109
rect 359096 280100 359148 280152
rect 359188 280100 359240 280152
rect 372712 280143 372764 280152
rect 372712 280109 372721 280143
rect 372721 280109 372755 280143
rect 372755 280109 372764 280143
rect 372712 280100 372764 280109
rect 377128 280143 377180 280152
rect 377128 280109 377137 280143
rect 377137 280109 377171 280143
rect 377171 280109 377180 280143
rect 377128 280100 377180 280109
rect 460112 280143 460164 280152
rect 460112 280109 460121 280143
rect 460121 280109 460155 280143
rect 460155 280109 460164 280143
rect 460112 280100 460164 280109
rect 250076 278740 250128 278792
rect 250168 278740 250220 278792
rect 265256 278876 265308 278928
rect 285772 278740 285824 278792
rect 286048 278740 286100 278792
rect 288716 278740 288768 278792
rect 288808 278740 288860 278792
rect 294236 278740 294288 278792
rect 294328 278740 294380 278792
rect 323216 278740 323268 278792
rect 323308 278740 323360 278792
rect 325884 278783 325936 278792
rect 325884 278749 325893 278783
rect 325893 278749 325927 278783
rect 325927 278749 325936 278783
rect 325884 278740 325936 278749
rect 337108 278783 337160 278792
rect 337108 278749 337117 278783
rect 337117 278749 337151 278783
rect 337151 278749 337160 278783
rect 337108 278740 337160 278749
rect 265348 278672 265400 278724
rect 310888 278715 310940 278724
rect 310888 278681 310897 278715
rect 310897 278681 310931 278715
rect 310931 278681 310940 278715
rect 310888 278672 310940 278681
rect 386788 278715 386840 278724
rect 386788 278681 386797 278715
rect 386797 278681 386831 278715
rect 386831 278681 386840 278715
rect 386788 278672 386840 278681
rect 291568 277448 291620 277500
rect 291568 277312 291620 277364
rect 266728 276063 266780 276072
rect 266728 276029 266737 276063
rect 266737 276029 266771 276063
rect 266771 276029 266780 276063
rect 266728 276020 266780 276029
rect 297088 276020 297140 276072
rect 463792 275315 463844 275324
rect 463792 275281 463801 275315
rect 463801 275281 463835 275315
rect 463835 275281 463844 275315
rect 463792 275272 463844 275281
rect 266636 274635 266688 274644
rect 266636 274601 266645 274635
rect 266645 274601 266679 274635
rect 266679 274601 266688 274635
rect 266636 274592 266688 274601
rect 330116 273955 330168 273964
rect 330116 273921 330125 273955
rect 330125 273921 330159 273955
rect 330159 273921 330168 273955
rect 330116 273912 330168 273921
rect 250168 273300 250220 273352
rect 250076 273164 250128 273216
rect 460112 273139 460164 273148
rect 460112 273105 460121 273139
rect 460121 273105 460155 273139
rect 460155 273105 460164 273139
rect 460112 273096 460164 273105
rect 259552 273071 259604 273080
rect 259552 273037 259561 273071
rect 259561 273037 259595 273071
rect 259595 273037 259604 273071
rect 259552 273028 259604 273037
rect 367008 270648 367060 270700
rect 236276 270555 236328 270564
rect 236276 270521 236285 270555
rect 236285 270521 236319 270555
rect 236319 270521 236328 270555
rect 236276 270512 236328 270521
rect 239220 270512 239272 270564
rect 251456 270555 251508 270564
rect 251456 270521 251465 270555
rect 251465 270521 251499 270555
rect 251499 270521 251508 270555
rect 251456 270512 251508 270521
rect 324688 270512 324740 270564
rect 324780 270512 324832 270564
rect 325884 270512 325936 270564
rect 325976 270512 326028 270564
rect 336924 270555 336976 270564
rect 336924 270521 336933 270555
rect 336933 270521 336967 270555
rect 336967 270521 336976 270555
rect 336924 270512 336976 270521
rect 367008 270512 367060 270564
rect 372712 270555 372764 270564
rect 372712 270521 372721 270555
rect 372721 270521 372755 270555
rect 372755 270521 372764 270555
rect 372712 270512 372764 270521
rect 377128 270555 377180 270564
rect 377128 270521 377137 270555
rect 377137 270521 377171 270555
rect 377171 270521 377180 270555
rect 377128 270512 377180 270521
rect 463884 270512 463936 270564
rect 341248 270444 341300 270496
rect 460112 270444 460164 270496
rect 470600 270487 470652 270496
rect 470600 270453 470609 270487
rect 470609 270453 470643 270487
rect 470643 270453 470652 270487
rect 470600 270444 470652 270453
rect 302700 269152 302752 269204
rect 306932 269152 306984 269204
rect 262496 269084 262548 269136
rect 262588 269084 262640 269136
rect 284576 269084 284628 269136
rect 284760 269084 284812 269136
rect 290096 269084 290148 269136
rect 290188 269084 290240 269136
rect 301044 269084 301096 269136
rect 301228 269084 301280 269136
rect 302608 269084 302660 269136
rect 306840 269084 306892 269136
rect 358544 269084 358596 269136
rect 358636 269084 358688 269136
rect 421196 269084 421248 269136
rect 421380 269084 421432 269136
rect 250076 269059 250128 269068
rect 250076 269025 250085 269059
rect 250085 269025 250119 269059
rect 250119 269025 250128 269059
rect 250076 269016 250128 269025
rect 288716 267724 288768 267776
rect 288808 267724 288860 267776
rect 291568 267724 291620 267776
rect 291660 267724 291712 267776
rect 295616 267724 295668 267776
rect 295800 267724 295852 267776
rect 294236 264936 294288 264988
rect 294328 264936 294380 264988
rect 270684 263576 270736 263628
rect 339684 263576 339736 263628
rect 339868 263576 339920 263628
rect 360292 263576 360344 263628
rect 360476 263576 360528 263628
rect 270684 263440 270736 263492
rect 310888 263483 310940 263492
rect 310888 263449 310897 263483
rect 310897 263449 310931 263483
rect 310931 263449 310940 263483
rect 310888 263440 310940 263449
rect 386788 263483 386840 263492
rect 386788 263449 386797 263483
rect 386797 263449 386831 263483
rect 386831 263449 386840 263483
rect 386788 263440 386840 263449
rect 325976 260924 326028 260976
rect 460020 260967 460072 260976
rect 460020 260933 460029 260967
rect 460029 260933 460063 260967
rect 460063 260933 460072 260967
rect 460020 260924 460072 260933
rect 284576 260856 284628 260908
rect 284760 260856 284812 260908
rect 236460 260788 236512 260840
rect 239128 260831 239180 260840
rect 239128 260797 239137 260831
rect 239137 260797 239171 260831
rect 239171 260797 239180 260831
rect 239128 260788 239180 260797
rect 251456 260831 251508 260840
rect 251456 260797 251465 260831
rect 251465 260797 251499 260831
rect 251499 260797 251508 260831
rect 251456 260788 251508 260797
rect 259552 260831 259604 260840
rect 259552 260797 259561 260831
rect 259561 260797 259595 260831
rect 259595 260797 259604 260831
rect 259552 260788 259604 260797
rect 262588 260788 262640 260840
rect 266636 260831 266688 260840
rect 266636 260797 266645 260831
rect 266645 260797 266679 260831
rect 266679 260797 266688 260831
rect 266636 260788 266688 260797
rect 267740 260788 267792 260840
rect 270684 260831 270736 260840
rect 270684 260797 270693 260831
rect 270693 260797 270727 260831
rect 270727 260797 270736 260831
rect 270684 260788 270736 260797
rect 273536 260788 273588 260840
rect 273628 260788 273680 260840
rect 262680 260720 262732 260772
rect 330116 260899 330168 260908
rect 330116 260865 330125 260899
rect 330125 260865 330159 260899
rect 330159 260865 330168 260899
rect 330116 260856 330168 260865
rect 341156 260899 341208 260908
rect 341156 260865 341165 260899
rect 341165 260865 341199 260899
rect 341199 260865 341208 260899
rect 341156 260856 341208 260865
rect 470600 260899 470652 260908
rect 470600 260865 470609 260899
rect 470609 260865 470643 260899
rect 470643 260865 470652 260899
rect 470600 260856 470652 260865
rect 336924 260831 336976 260840
rect 336924 260797 336933 260831
rect 336933 260797 336967 260831
rect 336967 260797 336976 260831
rect 336924 260788 336976 260797
rect 372712 260831 372764 260840
rect 372712 260797 372721 260831
rect 372721 260797 372755 260831
rect 372755 260797 372764 260831
rect 372712 260788 372764 260797
rect 377128 260831 377180 260840
rect 377128 260797 377137 260831
rect 377137 260797 377171 260831
rect 377171 260797 377180 260831
rect 377128 260788 377180 260797
rect 460020 260788 460072 260840
rect 460204 260788 460256 260840
rect 463792 260788 463844 260840
rect 267832 260720 267884 260772
rect 325976 260720 326028 260772
rect 327264 259564 327316 259616
rect 250168 259428 250220 259480
rect 272064 259428 272116 259480
rect 272156 259428 272208 259480
rect 336924 259428 336976 259480
rect 337108 259428 337160 259480
rect 299848 259360 299900 259412
rect 300032 259360 300084 259412
rect 302608 259360 302660 259412
rect 302792 259360 302844 259412
rect 327264 259360 327316 259412
rect 358728 259403 358780 259412
rect 358728 259369 358737 259403
rect 358737 259369 358771 259403
rect 358771 259369 358780 259403
rect 358728 259360 358780 259369
rect 250168 259335 250220 259344
rect 250168 259301 250177 259335
rect 250177 259301 250211 259335
rect 250211 259301 250220 259335
rect 250168 259292 250220 259301
rect 267832 258000 267884 258052
rect 272432 258000 272484 258052
rect 268016 257932 268068 257984
rect 295708 256640 295760 256692
rect 295892 256640 295944 256692
rect 310888 256071 310940 256080
rect 310888 256037 310897 256071
rect 310897 256037 310931 256071
rect 310931 256037 310940 256071
rect 310888 256028 310940 256037
rect 265348 255935 265400 255944
rect 265348 255901 265357 255935
rect 265357 255901 265391 255935
rect 265391 255901 265400 255935
rect 265348 255892 265400 255901
rect 337292 254600 337344 254652
rect 323400 253988 323452 254040
rect 327264 253920 327316 253972
rect 386788 253988 386840 254040
rect 323308 253852 323360 253904
rect 357532 253852 357584 253904
rect 357716 253852 357768 253904
rect 359004 253852 359056 253904
rect 359188 253852 359240 253904
rect 386696 253852 386748 253904
rect 259552 253759 259604 253768
rect 259552 253725 259561 253759
rect 259561 253725 259595 253759
rect 259595 253725 259604 253759
rect 259552 253716 259604 253725
rect 2780 252492 2832 252544
rect 5264 252492 5316 252544
rect 469956 252492 470008 252544
rect 580172 252492 580224 252544
rect 236276 251243 236328 251252
rect 236276 251209 236285 251243
rect 236285 251209 236319 251243
rect 236319 251209 236328 251243
rect 236276 251200 236328 251209
rect 239220 251200 239272 251252
rect 251456 251243 251508 251252
rect 251456 251209 251465 251243
rect 251465 251209 251499 251243
rect 251499 251209 251508 251243
rect 251456 251200 251508 251209
rect 290004 251200 290056 251252
rect 290096 251200 290148 251252
rect 259552 251175 259604 251184
rect 259552 251141 259561 251175
rect 259561 251141 259595 251175
rect 259595 251141 259604 251175
rect 259552 251132 259604 251141
rect 266728 251132 266780 251184
rect 266820 251132 266872 251184
rect 296996 251268 297048 251320
rect 310704 251268 310756 251320
rect 372712 251243 372764 251252
rect 372712 251209 372721 251243
rect 372721 251209 372755 251243
rect 372755 251209 372764 251243
rect 372712 251200 372764 251209
rect 377128 251243 377180 251252
rect 377128 251209 377137 251243
rect 377137 251209 377171 251243
rect 377171 251209 377180 251243
rect 377128 251200 377180 251209
rect 463700 251243 463752 251252
rect 463700 251209 463709 251243
rect 463709 251209 463743 251243
rect 463743 251209 463752 251243
rect 463700 251200 463752 251209
rect 310704 251175 310756 251184
rect 310704 251141 310713 251175
rect 310713 251141 310747 251175
rect 310747 251141 310756 251175
rect 310704 251132 310756 251141
rect 367008 251175 367060 251184
rect 367008 251141 367017 251175
rect 367017 251141 367051 251175
rect 367051 251141 367060 251175
rect 367008 251132 367060 251141
rect 470600 251175 470652 251184
rect 470600 251141 470609 251175
rect 470609 251141 470643 251175
rect 470643 251141 470652 251175
rect 470600 251132 470652 251141
rect 250352 251064 250404 251116
rect 296812 251064 296864 251116
rect 284668 249840 284720 249892
rect 284760 249840 284812 249892
rect 285956 249772 286008 249824
rect 286048 249772 286100 249824
rect 336924 249815 336976 249824
rect 336924 249781 336933 249815
rect 336933 249781 336967 249815
rect 336967 249781 336976 249815
rect 336924 249772 336976 249781
rect 421196 249772 421248 249824
rect 421380 249772 421432 249824
rect 272432 249704 272484 249756
rect 284668 249747 284720 249756
rect 284668 249713 284677 249747
rect 284677 249713 284711 249747
rect 284711 249713 284720 249747
rect 284668 249704 284720 249713
rect 265348 248251 265400 248260
rect 265348 248217 265357 248251
rect 265357 248217 265391 248251
rect 265391 248217 265400 248251
rect 265348 248208 265400 248217
rect 290004 246984 290056 247036
rect 290372 246984 290424 247036
rect 294236 246984 294288 247036
rect 294420 246848 294472 246900
rect 288900 245599 288952 245608
rect 288900 245565 288909 245599
rect 288909 245565 288943 245599
rect 288943 245565 288952 245599
rect 288900 245556 288952 245565
rect 285956 244987 286008 244996
rect 285956 244953 285965 244987
rect 285965 244953 285999 244987
rect 285999 244953 286008 244987
rect 285956 244944 286008 244953
rect 339684 244264 339736 244316
rect 339868 244264 339920 244316
rect 341248 244332 341300 244384
rect 360292 244264 360344 244316
rect 360476 244264 360528 244316
rect 460112 244332 460164 244384
rect 341156 244196 341208 244248
rect 460020 244196 460072 244248
rect 259644 244128 259696 244180
rect 271880 243040 271932 243092
rect 272432 243040 272484 243092
rect 306840 241544 306892 241596
rect 236552 241476 236604 241528
rect 236644 241476 236696 241528
rect 266728 241476 266780 241528
rect 266820 241476 266872 241528
rect 324688 241544 324740 241596
rect 325976 241544 326028 241596
rect 337108 241587 337160 241596
rect 337108 241553 337117 241587
rect 337117 241553 337151 241587
rect 337151 241553 337160 241587
rect 337108 241544 337160 241553
rect 310888 241476 310940 241528
rect 323308 241476 323360 241528
rect 323400 241476 323452 241528
rect 324596 241476 324648 241528
rect 325884 241476 325936 241528
rect 357624 241476 357676 241528
rect 357716 241476 357768 241528
rect 359096 241476 359148 241528
rect 359188 241476 359240 241528
rect 367008 241519 367060 241528
rect 367008 241485 367017 241519
rect 367017 241485 367051 241519
rect 367051 241485 367060 241519
rect 367008 241476 367060 241485
rect 470600 241519 470652 241528
rect 470600 241485 470609 241519
rect 470609 241485 470643 241519
rect 470643 241485 470652 241519
rect 470600 241476 470652 241485
rect 299480 241451 299532 241460
rect 299480 241417 299489 241451
rect 299489 241417 299523 241451
rect 299523 241417 299532 241451
rect 299480 241408 299532 241417
rect 306840 241408 306892 241460
rect 259644 241340 259696 241392
rect 259828 241340 259880 241392
rect 270684 240227 270736 240236
rect 270684 240193 270693 240227
rect 270693 240193 270727 240227
rect 270727 240193 270736 240227
rect 270684 240184 270736 240193
rect 327172 240227 327224 240236
rect 327172 240193 327181 240227
rect 327181 240193 327215 240227
rect 327215 240193 327224 240227
rect 327172 240184 327224 240193
rect 284852 240116 284904 240168
rect 299940 240116 299992 240168
rect 300032 240116 300084 240168
rect 302700 240116 302752 240168
rect 302792 240116 302844 240168
rect 358728 240159 358780 240168
rect 358728 240125 358737 240159
rect 358737 240125 358771 240159
rect 358771 240125 358780 240159
rect 358728 240116 358780 240125
rect 267740 240048 267792 240100
rect 267924 240048 267976 240100
rect 291568 240048 291620 240100
rect 291844 240048 291896 240100
rect 324596 240091 324648 240100
rect 324596 240057 324605 240091
rect 324605 240057 324639 240091
rect 324639 240057 324648 240091
rect 324596 240048 324648 240057
rect 327172 240091 327224 240100
rect 327172 240057 327181 240091
rect 327181 240057 327215 240091
rect 327215 240057 327224 240091
rect 327172 240048 327224 240057
rect 270684 238731 270736 238740
rect 270684 238697 270693 238731
rect 270693 238697 270727 238731
rect 270727 238697 270736 238731
rect 270684 238688 270736 238697
rect 3056 237328 3108 237380
rect 15844 237328 15896 237380
rect 288992 235968 289044 236020
rect 262772 235900 262824 235952
rect 265164 234676 265216 234728
rect 265348 234676 265400 234728
rect 310888 234676 310940 234728
rect 323400 234719 323452 234728
rect 323400 234685 323409 234719
rect 323409 234685 323443 234719
rect 323443 234685 323452 234719
rect 323400 234676 323452 234685
rect 337200 234608 337252 234660
rect 273444 234540 273496 234592
rect 273628 234540 273680 234592
rect 310796 234540 310848 234592
rect 357532 234540 357584 234592
rect 357716 234540 357768 234592
rect 359004 234540 359056 234592
rect 359188 234540 359240 234592
rect 285956 234515 286008 234524
rect 285956 234481 285965 234515
rect 285965 234481 285999 234515
rect 285999 234481 286008 234515
rect 285956 234472 286008 234481
rect 270684 233835 270736 233844
rect 270684 233801 270693 233835
rect 270693 233801 270727 233835
rect 270727 233801 270736 233835
rect 270684 233792 270736 233801
rect 244280 231820 244332 231872
rect 244464 231820 244516 231872
rect 250076 231820 250128 231872
rect 250352 231820 250404 231872
rect 251456 231820 251508 231872
rect 251640 231820 251692 231872
rect 299480 231863 299532 231872
rect 299480 231829 299489 231863
rect 299489 231829 299523 231863
rect 299523 231829 299532 231863
rect 299480 231820 299532 231829
rect 299940 231820 299992 231872
rect 301136 231888 301188 231940
rect 372528 231820 372580 231872
rect 372712 231820 372764 231872
rect 376944 231820 376996 231872
rect 377128 231820 377180 231872
rect 299756 231752 299808 231804
rect 301044 231752 301096 231804
rect 310796 231795 310848 231804
rect 310796 231761 310805 231795
rect 310805 231761 310839 231795
rect 310839 231761 310848 231795
rect 310796 231752 310848 231761
rect 323400 231795 323452 231804
rect 323400 231761 323409 231795
rect 323409 231761 323443 231795
rect 323443 231761 323452 231795
rect 323400 231752 323452 231761
rect 324780 231752 324832 231804
rect 327172 230571 327224 230580
rect 327172 230537 327181 230571
rect 327181 230537 327215 230571
rect 327215 230537 327224 230571
rect 327172 230528 327224 230537
rect 325976 230460 326028 230512
rect 326160 230460 326212 230512
rect 336740 230460 336792 230512
rect 336924 230460 336976 230512
rect 337108 230503 337160 230512
rect 337108 230469 337117 230503
rect 337117 230469 337151 230503
rect 337151 230469 337160 230503
rect 337108 230460 337160 230469
rect 341248 230460 341300 230512
rect 341432 230460 341484 230512
rect 358452 230460 358504 230512
rect 358636 230460 358688 230512
rect 421196 230460 421248 230512
rect 421380 230460 421432 230512
rect 459836 230460 459888 230512
rect 460112 230460 460164 230512
rect 358544 230392 358596 230444
rect 265164 229032 265216 229084
rect 265532 229032 265584 229084
rect 272064 229075 272116 229084
rect 272064 229041 272073 229075
rect 272073 229041 272107 229075
rect 272107 229041 272116 229075
rect 272064 229032 272116 229041
rect 262588 226355 262640 226364
rect 262588 226321 262597 226355
rect 262597 226321 262631 226355
rect 262631 226321 262640 226355
rect 262588 226312 262640 226321
rect 336740 225428 336792 225480
rect 336924 225428 336976 225480
rect 284852 225020 284904 225072
rect 236276 224952 236328 225004
rect 339684 224952 339736 225004
rect 339868 224952 339920 225004
rect 341248 225020 341300 225072
rect 360292 224952 360344 225004
rect 360476 224952 360528 225004
rect 460112 225020 460164 225072
rect 284852 224884 284904 224936
rect 341156 224884 341208 224936
rect 460020 224884 460072 224936
rect 236460 224816 236512 224868
rect 306840 222300 306892 222352
rect 306932 222300 306984 222352
rect 259644 222164 259696 222216
rect 259828 222164 259880 222216
rect 294328 222164 294380 222216
rect 294420 222164 294472 222216
rect 295524 222164 295576 222216
rect 295616 222164 295668 222216
rect 296812 222164 296864 222216
rect 296904 222164 296956 222216
rect 299756 222164 299808 222216
rect 299940 222164 299992 222216
rect 310888 222164 310940 222216
rect 325884 222164 325936 222216
rect 326068 222164 326120 222216
rect 359096 222164 359148 222216
rect 359188 222164 359240 222216
rect 386604 222164 386656 222216
rect 386788 222164 386840 222216
rect 463792 222164 463844 222216
rect 464068 222164 464120 222216
rect 470416 222164 470468 222216
rect 470600 222164 470652 222216
rect 299480 222139 299532 222148
rect 299480 222105 299489 222139
rect 299489 222105 299523 222139
rect 299523 222105 299532 222139
rect 299480 222096 299532 222105
rect 259644 222028 259696 222080
rect 259828 222028 259880 222080
rect 273536 220804 273588 220856
rect 273628 220804 273680 220856
rect 327356 220804 327408 220856
rect 327540 220804 327592 220856
rect 330208 220804 330260 220856
rect 330392 220804 330444 220856
rect 358728 220847 358780 220856
rect 358728 220813 358737 220847
rect 358737 220813 358771 220847
rect 358771 220813 358780 220847
rect 358728 220804 358780 220813
rect 272156 220736 272208 220788
rect 341156 220779 341208 220788
rect 341156 220745 341165 220779
rect 341165 220745 341199 220779
rect 341199 220745 341208 220779
rect 341156 220736 341208 220745
rect 262588 219444 262640 219496
rect 270776 219376 270828 219428
rect 270960 219376 271012 219428
rect 317512 219376 317564 219428
rect 317696 219376 317748 219428
rect 262680 219308 262732 219360
rect 290096 217991 290148 218000
rect 290096 217957 290105 217991
rect 290105 217957 290139 217991
rect 290139 217957 290148 217991
rect 290096 217948 290148 217957
rect 310888 215364 310940 215416
rect 386420 215296 386472 215348
rect 386604 215296 386656 215348
rect 464068 215364 464120 215416
rect 273444 215228 273496 215280
rect 273628 215228 273680 215280
rect 310796 215228 310848 215280
rect 341156 215271 341208 215280
rect 341156 215237 341165 215271
rect 341165 215237 341199 215271
rect 341199 215237 341208 215271
rect 341156 215228 341208 215237
rect 459836 215228 459888 215280
rect 460020 215228 460072 215280
rect 463976 215228 464028 215280
rect 291660 214591 291712 214600
rect 291660 214557 291669 214591
rect 291669 214557 291703 214591
rect 291703 214557 291712 214591
rect 291660 214548 291712 214557
rect 244280 212508 244332 212560
rect 244464 212508 244516 212560
rect 250076 212508 250128 212560
rect 250352 212508 250404 212560
rect 251456 212508 251508 212560
rect 251640 212508 251692 212560
rect 299480 212551 299532 212560
rect 299480 212517 299489 212551
rect 299489 212517 299523 212551
rect 299523 212517 299532 212551
rect 299480 212508 299532 212517
rect 299940 212576 299992 212628
rect 301136 212576 301188 212628
rect 324688 212508 324740 212560
rect 324780 212508 324832 212560
rect 325884 212508 325936 212560
rect 325976 212508 326028 212560
rect 336740 212508 336792 212560
rect 336924 212508 336976 212560
rect 357624 212508 357676 212560
rect 357716 212508 357768 212560
rect 359096 212508 359148 212560
rect 359188 212508 359240 212560
rect 372528 212508 372580 212560
rect 372712 212508 372764 212560
rect 376944 212508 376996 212560
rect 377128 212508 377180 212560
rect 284668 212440 284720 212492
rect 284852 212440 284904 212492
rect 299756 212440 299808 212492
rect 301044 212440 301096 212492
rect 310796 212483 310848 212492
rect 310796 212449 310805 212483
rect 310805 212449 310839 212483
rect 310839 212449 310848 212483
rect 310796 212440 310848 212449
rect 330208 212440 330260 212492
rect 330300 212440 330352 212492
rect 250076 211080 250128 211132
rect 250260 211080 250312 211132
rect 284668 211080 284720 211132
rect 284944 211080 284996 211132
rect 317512 209788 317564 209840
rect 317696 209788 317748 209840
rect 290096 208403 290148 208412
rect 290096 208369 290105 208403
rect 290105 208369 290139 208403
rect 290139 208369 290148 208403
rect 290096 208360 290148 208369
rect 323308 205640 323360 205692
rect 339684 205640 339736 205692
rect 339868 205640 339920 205692
rect 360292 205640 360344 205692
rect 360476 205640 360528 205692
rect 460112 205708 460164 205760
rect 460020 205572 460072 205624
rect 323400 205504 323452 205556
rect 291660 204051 291712 204060
rect 291660 204017 291669 204051
rect 291669 204017 291703 204051
rect 291703 204017 291712 204051
rect 291660 204008 291712 204017
rect 262588 202852 262640 202904
rect 262680 202852 262732 202904
rect 266636 202852 266688 202904
rect 266728 202852 266780 202904
rect 285956 202852 286008 202904
rect 286140 202852 286192 202904
rect 294236 202852 294288 202904
rect 294328 202852 294380 202904
rect 295524 202852 295576 202904
rect 295616 202852 295668 202904
rect 296812 202852 296864 202904
rect 296904 202852 296956 202904
rect 299756 202852 299808 202904
rect 299940 202852 299992 202904
rect 310888 202852 310940 202904
rect 324596 202852 324648 202904
rect 324688 202852 324740 202904
rect 325884 202852 325936 202904
rect 325976 202852 326028 202904
rect 341156 202852 341208 202904
rect 341248 202852 341300 202904
rect 463792 202852 463844 202904
rect 464068 202852 464120 202904
rect 470416 202852 470468 202904
rect 470600 202852 470652 202904
rect 239128 202784 239180 202836
rect 239220 202784 239272 202836
rect 273536 202784 273588 202836
rect 273628 202784 273680 202836
rect 299480 202827 299532 202836
rect 299480 202793 299489 202827
rect 299489 202793 299523 202827
rect 299523 202793 299532 202827
rect 336924 202827 336976 202836
rect 299480 202784 299532 202793
rect 336924 202793 336933 202827
rect 336933 202793 336967 202827
rect 336967 202793 336976 202827
rect 336924 202784 336976 202793
rect 270500 202104 270552 202156
rect 270960 202104 271012 202156
rect 290096 201492 290148 201544
rect 250076 201424 250128 201476
rect 250352 201424 250404 201476
rect 262588 201424 262640 201476
rect 262772 201424 262824 201476
rect 272340 201467 272392 201476
rect 272340 201433 272349 201467
rect 272349 201433 272383 201467
rect 272383 201433 272392 201467
rect 272340 201424 272392 201433
rect 267740 201356 267792 201408
rect 267924 201356 267976 201408
rect 358452 201424 358504 201476
rect 358728 201424 358780 201476
rect 421196 201424 421248 201476
rect 421380 201424 421432 201476
rect 290188 201356 290240 201408
rect 250076 200107 250128 200116
rect 250076 200073 250085 200107
rect 250085 200073 250119 200107
rect 250119 200073 250128 200107
rect 250076 200064 250128 200073
rect 265164 200107 265216 200116
rect 265164 200073 265173 200107
rect 265173 200073 265207 200107
rect 265207 200073 265216 200107
rect 265164 200064 265216 200073
rect 317512 200064 317564 200116
rect 317696 200064 317748 200116
rect 285772 198024 285824 198076
rect 285956 198024 286008 198076
rect 294236 198024 294288 198076
rect 294420 198024 294472 198076
rect 232228 195984 232280 196036
rect 310888 196052 310940 196104
rect 337108 195984 337160 196036
rect 460020 195984 460072 196036
rect 232320 195916 232372 195968
rect 310796 195916 310848 195968
rect 337200 195916 337252 195968
rect 357532 195916 357584 195968
rect 357716 195916 357768 195968
rect 359004 195916 359056 195968
rect 359188 195916 359240 195968
rect 464068 196052 464120 196104
rect 463976 195916 464028 195968
rect 460112 195848 460164 195900
rect 270500 195780 270552 195832
rect 270684 195780 270736 195832
rect 265164 195279 265216 195288
rect 265164 195245 265173 195279
rect 265173 195245 265207 195279
rect 265207 195245 265216 195279
rect 265164 195236 265216 195245
rect 244280 193196 244332 193248
rect 244464 193196 244516 193248
rect 251456 193196 251508 193248
rect 251640 193196 251692 193248
rect 259736 193196 259788 193248
rect 259920 193196 259972 193248
rect 290188 193264 290240 193316
rect 299480 193239 299532 193248
rect 299480 193205 299489 193239
rect 299489 193205 299523 193239
rect 299523 193205 299532 193239
rect 299480 193196 299532 193205
rect 302700 193264 302752 193316
rect 323308 193196 323360 193248
rect 323492 193196 323544 193248
rect 324596 193196 324648 193248
rect 324688 193196 324740 193248
rect 325884 193196 325936 193248
rect 325976 193196 326028 193248
rect 336924 193239 336976 193248
rect 336924 193205 336933 193239
rect 336933 193205 336967 193239
rect 336967 193205 336976 193239
rect 336924 193196 336976 193205
rect 341248 193196 341300 193248
rect 341432 193196 341484 193248
rect 372528 193196 372580 193248
rect 372712 193196 372764 193248
rect 376944 193196 376996 193248
rect 377128 193196 377180 193248
rect 386696 193196 386748 193248
rect 386880 193196 386932 193248
rect 272340 193171 272392 193180
rect 272340 193137 272349 193171
rect 272349 193137 272383 193171
rect 272383 193137 272392 193171
rect 272340 193128 272392 193137
rect 290096 193128 290148 193180
rect 302516 193128 302568 193180
rect 367008 193171 367060 193180
rect 367008 193137 367017 193171
rect 367017 193137 367051 193171
rect 367051 193137 367060 193171
rect 367008 193128 367060 193137
rect 266636 191811 266688 191820
rect 266636 191777 266645 191811
rect 266645 191777 266679 191811
rect 266679 191777 266688 191811
rect 266636 191768 266688 191777
rect 270684 191768 270736 191820
rect 270868 191768 270920 191820
rect 288808 191811 288860 191820
rect 288808 191777 288817 191811
rect 288817 191777 288851 191811
rect 288851 191777 288860 191811
rect 288808 191768 288860 191777
rect 291568 191768 291620 191820
rect 291660 191768 291712 191820
rect 317512 190476 317564 190528
rect 317696 190476 317748 190528
rect 270868 190408 270920 190460
rect 271052 190408 271104 190460
rect 290096 188640 290148 188692
rect 299848 188479 299900 188488
rect 299848 188445 299857 188479
rect 299857 188445 299891 188479
rect 299891 188445 299900 188479
rect 299848 188436 299900 188445
rect 306840 188479 306892 188488
rect 306840 188445 306849 188479
rect 306849 188445 306883 188479
rect 306883 188445 306892 188479
rect 306840 188436 306892 188445
rect 264980 186940 265032 186992
rect 265164 186940 265216 186992
rect 295616 186396 295668 186448
rect 296904 186396 296956 186448
rect 327264 186396 327316 186448
rect 330208 186396 330260 186448
rect 250076 186303 250128 186312
rect 250076 186269 250085 186303
rect 250085 186269 250119 186303
rect 250119 186269 250128 186303
rect 250076 186260 250128 186269
rect 266636 186303 266688 186312
rect 266636 186269 266645 186303
rect 266645 186269 266679 186303
rect 266679 186269 266688 186303
rect 266636 186260 266688 186269
rect 272156 186260 272208 186312
rect 272432 186260 272484 186312
rect 295524 186260 295576 186312
rect 296812 186260 296864 186312
rect 327172 186260 327224 186312
rect 460020 186328 460072 186380
rect 460112 186260 460164 186312
rect 330208 186192 330260 186244
rect 294420 184220 294472 184272
rect 285956 183676 286008 183728
rect 284668 183608 284720 183660
rect 236460 183540 236512 183592
rect 236552 183540 236604 183592
rect 302516 183608 302568 183660
rect 285956 183540 286008 183592
rect 299848 183583 299900 183592
rect 299848 183549 299857 183583
rect 299857 183549 299891 183583
rect 299891 183549 299900 183583
rect 299848 183540 299900 183549
rect 301044 183540 301096 183592
rect 301228 183540 301280 183592
rect 302608 183540 302660 183592
rect 306840 183583 306892 183592
rect 306840 183549 306849 183583
rect 306849 183549 306883 183583
rect 306883 183549 306892 183583
rect 306840 183540 306892 183549
rect 310888 183540 310940 183592
rect 311072 183540 311124 183592
rect 358636 183540 358688 183592
rect 358728 183540 358780 183592
rect 359096 183540 359148 183592
rect 359188 183540 359240 183592
rect 360476 183540 360528 183592
rect 360660 183540 360712 183592
rect 367008 183583 367060 183592
rect 367008 183549 367017 183583
rect 367017 183549 367051 183583
rect 367051 183549 367060 183583
rect 367008 183540 367060 183549
rect 463792 183540 463844 183592
rect 464068 183540 464120 183592
rect 470416 183540 470468 183592
rect 470600 183540 470652 183592
rect 239128 183472 239180 183524
rect 239220 183472 239272 183524
rect 273536 183472 273588 183524
rect 273628 183472 273680 183524
rect 284668 183472 284720 183524
rect 337108 183515 337160 183524
rect 337108 183481 337117 183515
rect 337117 183481 337151 183515
rect 337151 183481 337160 183515
rect 337108 183472 337160 183481
rect 460112 183515 460164 183524
rect 460112 183481 460121 183515
rect 460121 183481 460155 183515
rect 460155 183481 460164 183515
rect 460112 183472 460164 183481
rect 341156 182112 341208 182164
rect 341248 182112 341300 182164
rect 358544 182112 358596 182164
rect 358728 182112 358780 182164
rect 360476 182112 360528 182164
rect 360660 182112 360712 182164
rect 421196 182112 421248 182164
rect 421380 182112 421432 182164
rect 469864 182112 469916 182164
rect 580172 182112 580224 182164
rect 357624 180820 357676 180872
rect 357716 180820 357768 180872
rect 284668 180795 284720 180804
rect 284668 180761 284677 180795
rect 284677 180761 284711 180795
rect 284711 180761 284720 180795
rect 284668 180752 284720 180761
rect 299848 180795 299900 180804
rect 299848 180761 299857 180795
rect 299857 180761 299891 180795
rect 299891 180761 299900 180795
rect 299848 180752 299900 180761
rect 301044 180795 301096 180804
rect 301044 180761 301053 180795
rect 301053 180761 301087 180795
rect 301087 180761 301096 180795
rect 301044 180752 301096 180761
rect 302608 180795 302660 180804
rect 302608 180761 302617 180795
rect 302617 180761 302651 180795
rect 302651 180761 302660 180795
rect 302608 180752 302660 180761
rect 317512 180752 317564 180804
rect 317696 180752 317748 180804
rect 259644 179571 259696 179580
rect 259644 179537 259653 179571
rect 259653 179537 259687 179571
rect 259687 179537 259696 179571
rect 259644 179528 259696 179537
rect 288808 179435 288860 179444
rect 288808 179401 288817 179435
rect 288817 179401 288851 179435
rect 288851 179401 288860 179435
rect 288808 179392 288860 179401
rect 290004 179435 290056 179444
rect 290004 179401 290013 179435
rect 290013 179401 290047 179435
rect 290047 179401 290056 179435
rect 290004 179392 290056 179401
rect 294328 179435 294380 179444
rect 294328 179401 294337 179435
rect 294337 179401 294371 179435
rect 294371 179401 294380 179435
rect 294328 179392 294380 179401
rect 295524 178712 295576 178764
rect 295708 178712 295760 178764
rect 296812 178712 296864 178764
rect 296996 178712 297048 178764
rect 294328 177964 294380 178016
rect 250076 177284 250128 177336
rect 250352 177284 250404 177336
rect 232228 176672 232280 176724
rect 310888 176740 310940 176792
rect 357624 176740 357676 176792
rect 463884 176672 463936 176724
rect 464068 176672 464120 176724
rect 232320 176604 232372 176656
rect 288808 176647 288860 176656
rect 288808 176613 288817 176647
rect 288817 176613 288851 176647
rect 288851 176613 288860 176647
rect 288808 176604 288860 176613
rect 310796 176604 310848 176656
rect 357624 176604 357676 176656
rect 372712 176604 372764 176656
rect 372804 176536 372856 176588
rect 460112 176511 460164 176520
rect 460112 176477 460121 176511
rect 460121 176477 460155 176511
rect 460155 176477 460164 176511
rect 460112 176468 460164 176477
rect 259736 173952 259788 174004
rect 236276 173884 236328 173936
rect 236644 173884 236696 173936
rect 251456 173884 251508 173936
rect 251640 173884 251692 173936
rect 262588 173884 262640 173936
rect 262680 173884 262732 173936
rect 266636 173884 266688 173936
rect 266820 173884 266872 173936
rect 267740 173884 267792 173936
rect 267832 173884 267884 173936
rect 323308 173884 323360 173936
rect 323492 173884 323544 173936
rect 324688 173884 324740 173936
rect 324780 173884 324832 173936
rect 325884 173884 325936 173936
rect 325976 173884 326028 173936
rect 327172 173884 327224 173936
rect 327264 173884 327316 173936
rect 336740 173884 336792 173936
rect 336924 173884 336976 173936
rect 376944 173884 376996 173936
rect 377036 173884 377088 173936
rect 386788 173884 386840 173936
rect 386972 173884 387024 173936
rect 339684 173816 339736 173868
rect 339960 173816 340012 173868
rect 270776 172524 270828 172576
rect 272248 172524 272300 172576
rect 272340 172524 272392 172576
rect 337108 172567 337160 172576
rect 337108 172533 337117 172567
rect 337117 172533 337151 172567
rect 337151 172533 337160 172567
rect 337108 172524 337160 172533
rect 330116 172499 330168 172508
rect 330116 172465 330125 172499
rect 330125 172465 330159 172499
rect 330159 172465 330168 172499
rect 330116 172456 330168 172465
rect 270868 172388 270920 172440
rect 284760 171096 284812 171148
rect 299848 171139 299900 171148
rect 299848 171105 299857 171139
rect 299857 171105 299891 171139
rect 299891 171105 299900 171139
rect 299848 171096 299900 171105
rect 301044 171139 301096 171148
rect 301044 171105 301053 171139
rect 301053 171105 301087 171139
rect 301087 171105 301096 171139
rect 301044 171096 301096 171105
rect 302608 171139 302660 171148
rect 302608 171105 302617 171139
rect 302617 171105 302651 171139
rect 302651 171105 302660 171139
rect 302608 171096 302660 171105
rect 306656 171096 306708 171148
rect 306932 171096 306984 171148
rect 286048 171028 286100 171080
rect 337108 169260 337160 169312
rect 337384 169260 337436 169312
rect 259736 169056 259788 169108
rect 259920 169056 259972 169108
rect 294328 168376 294380 168428
rect 272064 167628 272116 167680
rect 272248 167628 272300 167680
rect 357440 167628 357492 167680
rect 357624 167628 357676 167680
rect 270868 167084 270920 167136
rect 288808 167059 288860 167068
rect 288808 167025 288817 167059
rect 288817 167025 288851 167059
rect 288851 167025 288860 167059
rect 288808 167016 288860 167025
rect 310796 167016 310848 167068
rect 270684 166948 270736 167000
rect 460112 166991 460164 167000
rect 460112 166957 460121 166991
rect 460121 166957 460155 166991
rect 460155 166957 460164 166991
rect 460112 166948 460164 166957
rect 310888 166880 310940 166932
rect 2780 165452 2832 165504
rect 5172 165452 5224 165504
rect 262680 164296 262732 164348
rect 265256 164296 265308 164348
rect 267832 164296 267884 164348
rect 262588 164228 262640 164280
rect 265164 164228 265216 164280
rect 267740 164228 267792 164280
rect 239128 164160 239180 164212
rect 239220 164160 239272 164212
rect 244280 164160 244332 164212
rect 244464 164160 244516 164212
rect 251456 164160 251508 164212
rect 251640 164160 251692 164212
rect 259644 164160 259696 164212
rect 259828 164160 259880 164212
rect 372804 164203 372856 164212
rect 372804 164169 372813 164203
rect 372813 164169 372847 164203
rect 372847 164169 372856 164203
rect 372804 164160 372856 164169
rect 386512 164160 386564 164212
rect 386696 164160 386748 164212
rect 330116 162979 330168 162988
rect 330116 162945 330125 162979
rect 330125 162945 330159 162979
rect 330159 162945 330168 162979
rect 330116 162936 330168 162945
rect 232136 162800 232188 162852
rect 232228 162800 232280 162852
rect 358544 162800 358596 162852
rect 358728 162800 358780 162852
rect 421196 162843 421248 162852
rect 421196 162809 421205 162843
rect 421205 162809 421239 162843
rect 421239 162809 421248 162843
rect 421196 162800 421248 162809
rect 357532 162732 357584 162784
rect 357624 162732 357676 162784
rect 285956 161483 286008 161492
rect 285956 161449 285965 161483
rect 285965 161449 285999 161483
rect 285999 161449 286008 161483
rect 285956 161440 286008 161449
rect 460112 161483 460164 161492
rect 460112 161449 460121 161483
rect 460121 161449 460155 161483
rect 460155 161449 460164 161483
rect 460112 161440 460164 161449
rect 302516 161372 302568 161424
rect 302608 161372 302660 161424
rect 330116 161415 330168 161424
rect 330116 161381 330125 161415
rect 330125 161381 330159 161415
rect 330159 161381 330168 161415
rect 330116 161372 330168 161381
rect 295616 160080 295668 160132
rect 295708 160080 295760 160132
rect 296904 160080 296956 160132
rect 296996 160080 297048 160132
rect 306380 160012 306432 160064
rect 306840 160012 306892 160064
rect 285956 158652 286008 158704
rect 294328 158695 294380 158704
rect 294328 158661 294337 158695
rect 294337 158661 294371 158695
rect 294371 158661 294380 158695
rect 294328 158652 294380 158661
rect 272156 158015 272208 158024
rect 272156 157981 272165 158015
rect 272165 157981 272199 158015
rect 272199 157981 272208 158015
rect 272156 157972 272208 157981
rect 337016 157972 337068 158024
rect 337200 157972 337252 158024
rect 364340 157564 364392 157616
rect 373816 157564 373868 157616
rect 396080 157496 396132 157548
rect 400772 157496 400824 157548
rect 417884 157496 417936 157548
rect 418160 157496 418212 157548
rect 437204 157496 437256 157548
rect 437480 157496 437532 157548
rect 456524 157496 456576 157548
rect 458272 157496 458324 157548
rect 267740 157428 267792 157480
rect 265164 157360 265216 157412
rect 325884 157360 325936 157412
rect 327172 157360 327224 157412
rect 267740 157292 267792 157344
rect 265256 157224 265308 157276
rect 359096 157292 359148 157344
rect 372804 157335 372856 157344
rect 372804 157301 372813 157335
rect 372813 157301 372847 157335
rect 372847 157301 372856 157335
rect 372804 157292 372856 157301
rect 377128 157292 377180 157344
rect 327264 157224 327316 157276
rect 359188 157224 359240 157276
rect 377220 157224 377272 157276
rect 325976 157156 326028 157208
rect 247224 154572 247276 154624
rect 247316 154572 247368 154624
rect 299756 154504 299808 154556
rect 299848 154504 299900 154556
rect 470416 154504 470468 154556
rect 470600 154504 470652 154556
rect 301044 154436 301096 154488
rect 301228 154436 301280 154488
rect 259828 154164 259880 154216
rect 421196 153255 421248 153264
rect 421196 153221 421205 153255
rect 421205 153221 421239 153255
rect 421239 153221 421248 153255
rect 421196 153212 421248 153221
rect 290004 153144 290056 153196
rect 290096 153144 290148 153196
rect 291476 153144 291528 153196
rect 291568 153144 291620 153196
rect 295524 153144 295576 153196
rect 295616 153144 295668 153196
rect 310796 153187 310848 153196
rect 310796 153153 310805 153187
rect 310805 153153 310839 153187
rect 310839 153153 310848 153187
rect 310796 153144 310848 153153
rect 341156 153187 341208 153196
rect 341156 153153 341165 153187
rect 341165 153153 341199 153187
rect 341199 153153 341208 153187
rect 341156 153144 341208 153153
rect 330116 151827 330168 151836
rect 330116 151793 330125 151827
rect 330125 151793 330159 151827
rect 330159 151793 330168 151827
rect 330116 151784 330168 151793
rect 3332 151716 3384 151768
rect 17224 151716 17276 151768
rect 460112 151759 460164 151768
rect 460112 151725 460121 151759
rect 460121 151725 460155 151759
rect 460155 151725 460164 151759
rect 460112 151716 460164 151725
rect 339500 149676 339552 149728
rect 339776 149676 339828 149728
rect 294328 149107 294380 149116
rect 294328 149073 294337 149107
rect 294337 149073 294371 149107
rect 294371 149073 294380 149107
rect 294328 149064 294380 149073
rect 272156 148971 272208 148980
rect 272156 148937 272165 148971
rect 272165 148937 272199 148971
rect 272199 148937 272208 148971
rect 272156 148928 272208 148937
rect 360384 147704 360436 147756
rect 463792 147704 463844 147756
rect 330116 147636 330168 147688
rect 310796 147611 310848 147620
rect 310796 147577 310805 147611
rect 310805 147577 310839 147611
rect 310839 147577 310848 147611
rect 310796 147568 310848 147577
rect 330208 147568 330260 147620
rect 266728 144916 266780 144968
rect 463700 144959 463752 144968
rect 463700 144925 463709 144959
rect 463709 144925 463743 144959
rect 463743 144925 463752 144959
rect 463700 144916 463752 144925
rect 244280 144848 244332 144900
rect 244464 144848 244516 144900
rect 247132 144848 247184 144900
rect 247224 144848 247276 144900
rect 262588 144848 262640 144900
rect 262772 144848 262824 144900
rect 267740 144848 267792 144900
rect 267924 144848 267976 144900
rect 270684 144891 270736 144900
rect 270684 144857 270693 144891
rect 270693 144857 270727 144891
rect 270727 144857 270736 144891
rect 270684 144848 270736 144857
rect 272156 144848 272208 144900
rect 272432 144848 272484 144900
rect 323308 144848 323360 144900
rect 323400 144848 323452 144900
rect 325884 144848 325936 144900
rect 326068 144848 326120 144900
rect 327172 144848 327224 144900
rect 327356 144848 327408 144900
rect 341340 144848 341392 144900
rect 360200 144891 360252 144900
rect 360200 144857 360209 144891
rect 360209 144857 360243 144891
rect 360243 144857 360252 144891
rect 360200 144848 360252 144857
rect 367008 144891 367060 144900
rect 367008 144857 367017 144891
rect 367017 144857 367051 144891
rect 367051 144857 367060 144891
rect 367008 144848 367060 144857
rect 386512 144848 386564 144900
rect 386696 144848 386748 144900
rect 266728 144780 266780 144832
rect 339684 144780 339736 144832
rect 339868 144780 339920 144832
rect 232320 143531 232372 143540
rect 232320 143497 232329 143531
rect 232329 143497 232363 143531
rect 232363 143497 232372 143531
rect 232320 143488 232372 143497
rect 272432 143531 272484 143540
rect 272432 143497 272441 143531
rect 272441 143497 272475 143531
rect 272475 143497 272484 143531
rect 272432 143488 272484 143497
rect 301044 143488 301096 143540
rect 301228 143488 301280 143540
rect 323308 143531 323360 143540
rect 323308 143497 323317 143531
rect 323317 143497 323351 143531
rect 323351 143497 323360 143531
rect 323308 143488 323360 143497
rect 324596 143531 324648 143540
rect 324596 143497 324605 143531
rect 324605 143497 324639 143531
rect 324639 143497 324648 143531
rect 324596 143488 324648 143497
rect 330208 143488 330260 143540
rect 421196 143531 421248 143540
rect 421196 143497 421205 143531
rect 421205 143497 421239 143531
rect 421239 143497 421248 143531
rect 421196 143488 421248 143497
rect 460112 142239 460164 142248
rect 460112 142205 460121 142239
rect 460121 142205 460155 142239
rect 460155 142205 460164 142239
rect 460112 142196 460164 142205
rect 259644 142171 259696 142180
rect 259644 142137 259653 142171
rect 259653 142137 259687 142171
rect 259687 142137 259696 142171
rect 259644 142128 259696 142137
rect 306380 142128 306432 142180
rect 307024 142128 307076 142180
rect 317512 142128 317564 142180
rect 317696 142128 317748 142180
rect 460112 142103 460164 142112
rect 460112 142069 460121 142103
rect 460121 142069 460155 142103
rect 460155 142069 460164 142103
rect 460112 142060 460164 142069
rect 259736 141992 259788 142044
rect 286048 140811 286100 140820
rect 286048 140777 286057 140811
rect 286057 140777 286091 140811
rect 286091 140777 286100 140811
rect 286048 140768 286100 140777
rect 288808 140700 288860 140752
rect 294236 140700 294288 140752
rect 294420 140700 294472 140752
rect 295524 140743 295576 140752
rect 295524 140709 295533 140743
rect 295533 140709 295567 140743
rect 295567 140709 295576 140743
rect 295524 140700 295576 140709
rect 377220 140020 377272 140072
rect 270684 139995 270736 140004
rect 270684 139961 270693 139995
rect 270693 139961 270727 139995
rect 270727 139961 270736 139995
rect 270684 139952 270736 139961
rect 294420 139383 294472 139392
rect 294420 139349 294429 139383
rect 294429 139349 294463 139383
rect 294463 139349 294472 139383
rect 294420 139340 294472 139349
rect 372804 138116 372856 138168
rect 290096 138048 290148 138100
rect 375748 138048 375800 138100
rect 239128 137980 239180 138032
rect 296812 137980 296864 138032
rect 297272 137980 297324 138032
rect 337108 137980 337160 138032
rect 375656 137980 375708 138032
rect 463700 137980 463752 138032
rect 239036 137912 239088 137964
rect 317512 137912 317564 137964
rect 317788 137912 317840 137964
rect 330116 137955 330168 137964
rect 330116 137921 330125 137955
rect 330125 137921 330159 137955
rect 330159 137921 330168 137955
rect 330116 137912 330168 137921
rect 337200 137912 337252 137964
rect 463884 137912 463936 137964
rect 2780 136484 2832 136536
rect 5080 136484 5132 136536
rect 367008 135303 367060 135312
rect 367008 135269 367017 135303
rect 367017 135269 367051 135303
rect 367051 135269 367060 135303
rect 367008 135260 367060 135269
rect 372712 135303 372764 135312
rect 372712 135269 372721 135303
rect 372721 135269 372755 135303
rect 372755 135269 372764 135303
rect 372712 135260 372764 135269
rect 377128 135303 377180 135312
rect 377128 135269 377137 135303
rect 377137 135269 377171 135303
rect 377171 135269 377180 135303
rect 377128 135260 377180 135269
rect 266636 135192 266688 135244
rect 266728 135192 266780 135244
rect 272432 135235 272484 135244
rect 272432 135201 272441 135235
rect 272441 135201 272475 135235
rect 272475 135201 272484 135235
rect 272432 135192 272484 135201
rect 358728 135235 358780 135244
rect 358728 135201 358737 135235
rect 358737 135201 358771 135235
rect 358771 135201 358780 135235
rect 358728 135192 358780 135201
rect 470416 135192 470468 135244
rect 470600 135192 470652 135244
rect 232320 133943 232372 133952
rect 232320 133909 232329 133943
rect 232329 133909 232363 133943
rect 232363 133909 232372 133943
rect 232320 133900 232372 133909
rect 307024 133900 307076 133952
rect 323308 133943 323360 133952
rect 323308 133909 323317 133943
rect 323317 133909 323351 133943
rect 323351 133909 323360 133943
rect 323308 133900 323360 133909
rect 421196 133943 421248 133952
rect 421196 133909 421205 133943
rect 421205 133909 421239 133943
rect 421239 133909 421248 133943
rect 421196 133900 421248 133909
rect 265256 133875 265308 133884
rect 265256 133841 265265 133875
rect 265265 133841 265299 133875
rect 265299 133841 265308 133875
rect 265256 133832 265308 133841
rect 307024 133764 307076 133816
rect 324688 132472 324740 132524
rect 460204 132472 460256 132524
rect 463700 132472 463752 132524
rect 463884 132472 463936 132524
rect 289912 132447 289964 132456
rect 289912 132413 289921 132447
rect 289921 132413 289955 132447
rect 289955 132413 289964 132447
rect 289912 132404 289964 132413
rect 337200 132447 337252 132456
rect 337200 132413 337209 132447
rect 337209 132413 337243 132447
rect 337243 132413 337252 132447
rect 337200 132404 337252 132413
rect 288624 131155 288676 131164
rect 288624 131121 288633 131155
rect 288633 131121 288667 131155
rect 288667 131121 288676 131155
rect 288624 131112 288676 131121
rect 295616 131112 295668 131164
rect 291476 131087 291528 131096
rect 291476 131053 291485 131087
rect 291485 131053 291519 131087
rect 291519 131053 291528 131087
rect 291476 131044 291528 131053
rect 297180 131044 297232 131096
rect 270500 130364 270552 130416
rect 270684 130364 270736 130416
rect 294420 129795 294472 129804
rect 294420 129761 294429 129795
rect 294429 129761 294463 129795
rect 294463 129761 294472 129795
rect 294420 129752 294472 129761
rect 250076 128324 250128 128376
rect 284668 128324 284720 128376
rect 302608 128324 302660 128376
rect 250168 128256 250220 128308
rect 284760 128256 284812 128308
rect 325976 128392 326028 128444
rect 327264 128392 327316 128444
rect 341248 128392 341300 128444
rect 339684 128324 339736 128376
rect 339868 128324 339920 128376
rect 325884 128256 325936 128308
rect 327172 128256 327224 128308
rect 341248 128256 341300 128308
rect 302608 128188 302660 128240
rect 272156 125808 272208 125860
rect 272432 125808 272484 125860
rect 358728 125647 358780 125656
rect 358728 125613 358737 125647
rect 358737 125613 358771 125647
rect 358771 125613 358780 125647
rect 358728 125604 358780 125613
rect 239128 125579 239180 125588
rect 239128 125545 239137 125579
rect 239137 125545 239171 125579
rect 239171 125545 239180 125579
rect 239128 125536 239180 125545
rect 251456 125579 251508 125588
rect 251456 125545 251465 125579
rect 251465 125545 251499 125579
rect 251499 125545 251508 125579
rect 251456 125536 251508 125545
rect 262588 125536 262640 125588
rect 262772 125536 262824 125588
rect 267740 125536 267792 125588
rect 267924 125536 267976 125588
rect 270684 125579 270736 125588
rect 270684 125545 270693 125579
rect 270693 125545 270727 125579
rect 270727 125545 270736 125579
rect 270684 125536 270736 125545
rect 272156 125536 272208 125588
rect 272432 125536 272484 125588
rect 317696 125536 317748 125588
rect 317972 125536 318024 125588
rect 325884 125536 325936 125588
rect 326068 125536 326120 125588
rect 327172 125536 327224 125588
rect 327356 125536 327408 125588
rect 336740 125536 336792 125588
rect 336924 125536 336976 125588
rect 339776 125579 339828 125588
rect 339776 125545 339785 125579
rect 339785 125545 339819 125579
rect 339819 125545 339828 125579
rect 339776 125536 339828 125545
rect 341248 125536 341300 125588
rect 259828 124219 259880 124228
rect 259828 124185 259837 124219
rect 259837 124185 259871 124219
rect 259871 124185 259880 124219
rect 259828 124176 259880 124185
rect 265256 124219 265308 124228
rect 265256 124185 265265 124219
rect 265265 124185 265299 124219
rect 265299 124185 265308 124219
rect 265256 124176 265308 124185
rect 360200 124176 360252 124228
rect 360384 124176 360436 124228
rect 232320 124151 232372 124160
rect 232320 124117 232329 124151
rect 232329 124117 232363 124151
rect 232363 124117 232372 124151
rect 232320 124108 232372 124117
rect 250168 124108 250220 124160
rect 272432 124151 272484 124160
rect 272432 124117 272441 124151
rect 272441 124117 272475 124151
rect 272475 124117 272484 124151
rect 272432 124108 272484 124117
rect 299848 124151 299900 124160
rect 299848 124117 299857 124151
rect 299857 124117 299891 124151
rect 299891 124117 299900 124151
rect 299848 124108 299900 124117
rect 306840 124151 306892 124160
rect 306840 124117 306849 124151
rect 306849 124117 306883 124151
rect 306883 124117 306892 124151
rect 306840 124108 306892 124117
rect 359096 124108 359148 124160
rect 359188 124108 359240 124160
rect 421196 124151 421248 124160
rect 421196 124117 421205 124151
rect 421205 124117 421239 124151
rect 421239 124117 421248 124151
rect 421196 124108 421248 124117
rect 460020 124040 460072 124092
rect 460204 124040 460256 124092
rect 284760 122748 284812 122800
rect 324688 122791 324740 122800
rect 324688 122757 324697 122791
rect 324697 122757 324731 122791
rect 324731 122757 324740 122791
rect 324688 122748 324740 122757
rect 291568 122680 291620 122732
rect 284760 122612 284812 122664
rect 2780 122272 2832 122324
rect 4988 122272 5040 122324
rect 288624 121456 288676 121508
rect 288900 121456 288952 121508
rect 294328 121456 294380 121508
rect 294420 121456 294472 121508
rect 296904 121499 296956 121508
rect 296904 121465 296913 121499
rect 296913 121465 296947 121499
rect 296947 121465 296956 121499
rect 296904 121456 296956 121465
rect 270684 120683 270736 120692
rect 270684 120649 270693 120683
rect 270693 120649 270727 120683
rect 270727 120649 270736 120683
rect 270684 120640 270736 120649
rect 273536 118668 273588 118720
rect 372712 118668 372764 118720
rect 377128 118668 377180 118720
rect 273628 118600 273680 118652
rect 339776 118643 339828 118652
rect 339776 118609 339785 118643
rect 339785 118609 339819 118643
rect 339819 118609 339828 118643
rect 339776 118600 339828 118609
rect 341156 118643 341208 118652
rect 341156 118609 341165 118643
rect 341165 118609 341199 118643
rect 341199 118609 341208 118643
rect 341156 118600 341208 118609
rect 372712 118532 372764 118584
rect 377128 118532 377180 118584
rect 327264 118464 327316 118516
rect 327356 118464 327408 118516
rect 262588 117988 262640 118040
rect 262772 117988 262824 118040
rect 239128 115991 239180 116000
rect 239128 115957 239137 115991
rect 239137 115957 239171 115991
rect 239171 115957 239180 115991
rect 239128 115948 239180 115957
rect 251456 115991 251508 116000
rect 251456 115957 251465 115991
rect 251465 115957 251499 115991
rect 251499 115957 251508 115991
rect 251456 115948 251508 115957
rect 341248 115880 341300 115932
rect 367008 115923 367060 115932
rect 367008 115889 367017 115923
rect 367017 115889 367051 115923
rect 367051 115889 367060 115923
rect 367008 115880 367060 115889
rect 376944 115880 376996 115932
rect 377128 115880 377180 115932
rect 470600 115923 470652 115932
rect 470600 115889 470609 115923
rect 470609 115889 470643 115923
rect 470643 115889 470652 115923
rect 470600 115880 470652 115889
rect 259828 115404 259880 115456
rect 259828 115268 259880 115320
rect 232320 114563 232372 114572
rect 232320 114529 232329 114563
rect 232329 114529 232363 114563
rect 232363 114529 232372 114563
rect 232320 114520 232372 114529
rect 249984 114563 250036 114572
rect 249984 114529 249993 114563
rect 249993 114529 250027 114563
rect 250027 114529 250036 114563
rect 249984 114520 250036 114529
rect 272432 114563 272484 114572
rect 272432 114529 272441 114563
rect 272441 114529 272475 114563
rect 272475 114529 272484 114563
rect 272432 114520 272484 114529
rect 296904 114588 296956 114640
rect 357532 114588 357584 114640
rect 299848 114563 299900 114572
rect 299848 114529 299857 114563
rect 299857 114529 299891 114563
rect 299891 114529 299900 114563
rect 299848 114520 299900 114529
rect 337200 114563 337252 114572
rect 337200 114529 337209 114563
rect 337209 114529 337243 114563
rect 337243 114529 337252 114563
rect 337200 114520 337252 114529
rect 357440 114520 357492 114572
rect 358636 114520 358688 114572
rect 358728 114520 358780 114572
rect 421196 114563 421248 114572
rect 421196 114529 421205 114563
rect 421205 114529 421239 114563
rect 421239 114529 421248 114563
rect 421196 114520 421248 114529
rect 296812 114452 296864 114504
rect 327264 114452 327316 114504
rect 306748 113228 306800 113280
rect 286048 113160 286100 113212
rect 286232 113160 286284 113212
rect 324688 113203 324740 113212
rect 324688 113169 324697 113203
rect 324697 113169 324731 113203
rect 324731 113169 324740 113203
rect 324688 113160 324740 113169
rect 265256 113135 265308 113144
rect 265256 113101 265265 113135
rect 265265 113101 265299 113135
rect 265299 113101 265308 113135
rect 265256 113092 265308 113101
rect 284668 113135 284720 113144
rect 284668 113101 284677 113135
rect 284677 113101 284711 113135
rect 284711 113101 284720 113135
rect 284668 113092 284720 113101
rect 291568 113135 291620 113144
rect 291568 113101 291577 113135
rect 291577 113101 291611 113135
rect 291611 113101 291620 113135
rect 291568 113092 291620 113101
rect 296812 113135 296864 113144
rect 296812 113101 296821 113135
rect 296821 113101 296855 113135
rect 296855 113101 296864 113135
rect 296812 113092 296864 113101
rect 306840 113092 306892 113144
rect 307024 113092 307076 113144
rect 329932 113092 329984 113144
rect 330208 113092 330260 113144
rect 286048 113024 286100 113076
rect 286232 113024 286284 113076
rect 270684 111052 270736 111104
rect 270868 111052 270920 111104
rect 463884 111052 463936 111104
rect 464068 111052 464120 111104
rect 294328 109735 294380 109744
rect 294328 109701 294337 109735
rect 294337 109701 294371 109735
rect 294371 109701 294380 109735
rect 294328 109692 294380 109701
rect 247224 109055 247276 109064
rect 247224 109021 247233 109055
rect 247233 109021 247267 109055
rect 247267 109021 247276 109055
rect 247224 109012 247276 109021
rect 310796 109012 310848 109064
rect 375656 109012 375708 109064
rect 310888 108944 310940 108996
rect 375564 108944 375616 108996
rect 272156 106496 272208 106548
rect 272432 106496 272484 106548
rect 247224 106335 247276 106344
rect 247224 106301 247233 106335
rect 247233 106301 247267 106335
rect 247267 106301 247276 106335
rect 247224 106292 247276 106301
rect 325976 106335 326028 106344
rect 325976 106301 325985 106335
rect 325985 106301 326019 106335
rect 326019 106301 326028 106335
rect 325976 106292 326028 106301
rect 341156 106335 341208 106344
rect 341156 106301 341165 106335
rect 341165 106301 341199 106335
rect 341199 106301 341208 106335
rect 341156 106292 341208 106301
rect 358636 106292 358688 106344
rect 367008 106335 367060 106344
rect 367008 106301 367017 106335
rect 367017 106301 367051 106335
rect 367051 106301 367060 106335
rect 367008 106292 367060 106301
rect 470600 106335 470652 106344
rect 470600 106301 470609 106335
rect 470609 106301 470643 106335
rect 470643 106301 470652 106335
rect 470600 106292 470652 106301
rect 236460 106224 236512 106276
rect 236644 106224 236696 106276
rect 239128 106224 239180 106276
rect 239312 106224 239364 106276
rect 251456 106267 251508 106276
rect 251456 106233 251465 106267
rect 251465 106233 251499 106267
rect 251499 106233 251508 106267
rect 251456 106224 251508 106233
rect 259736 106224 259788 106276
rect 259828 106224 259880 106276
rect 266728 106224 266780 106276
rect 266820 106224 266872 106276
rect 267832 106224 267884 106276
rect 267924 106224 267976 106276
rect 270684 106267 270736 106276
rect 270684 106233 270693 106267
rect 270693 106233 270727 106267
rect 270727 106233 270736 106267
rect 270684 106224 270736 106233
rect 272156 106224 272208 106276
rect 272432 106224 272484 106276
rect 360384 106224 360436 106276
rect 360568 106224 360620 106276
rect 372712 106224 372764 106276
rect 372804 106224 372856 106276
rect 386512 106267 386564 106276
rect 386512 106233 386521 106267
rect 386521 106233 386555 106267
rect 386555 106233 386564 106267
rect 386512 106224 386564 106233
rect 358728 106156 358780 106208
rect 289912 104864 289964 104916
rect 290004 104864 290056 104916
rect 317788 104864 317840 104916
rect 317972 104864 318024 104916
rect 325976 104907 326028 104916
rect 325976 104873 325985 104907
rect 325985 104873 326019 104907
rect 326019 104873 326028 104907
rect 325976 104864 326028 104873
rect 327172 104907 327224 104916
rect 327172 104873 327181 104907
rect 327181 104873 327215 104907
rect 327215 104873 327224 104907
rect 327172 104864 327224 104873
rect 339776 104864 339828 104916
rect 339868 104864 339920 104916
rect 357532 104864 357584 104916
rect 357716 104864 357768 104916
rect 232320 104839 232372 104848
rect 232320 104805 232329 104839
rect 232329 104805 232363 104839
rect 232363 104805 232372 104839
rect 232320 104796 232372 104805
rect 324596 104796 324648 104848
rect 324688 104796 324740 104848
rect 341156 104839 341208 104848
rect 341156 104805 341165 104839
rect 341165 104805 341199 104839
rect 341199 104805 341208 104839
rect 341156 104796 341208 104805
rect 421196 104839 421248 104848
rect 421196 104805 421205 104839
rect 421205 104805 421239 104839
rect 421239 104805 421248 104839
rect 421196 104796 421248 104805
rect 339776 104771 339828 104780
rect 339776 104737 339785 104771
rect 339785 104737 339819 104771
rect 339819 104737 339828 104771
rect 339776 104728 339828 104737
rect 358728 104728 358780 104780
rect 359004 104728 359056 104780
rect 291660 103572 291712 103624
rect 265256 103547 265308 103556
rect 265256 103513 265265 103547
rect 265265 103513 265299 103547
rect 265299 103513 265308 103547
rect 265256 103504 265308 103513
rect 284668 103547 284720 103556
rect 284668 103513 284677 103547
rect 284677 103513 284711 103547
rect 284711 103513 284720 103547
rect 284668 103504 284720 103513
rect 288808 103504 288860 103556
rect 288900 103504 288952 103556
rect 296812 103547 296864 103556
rect 296812 103513 296821 103547
rect 296821 103513 296855 103547
rect 296855 103513 296864 103547
rect 296812 103504 296864 103513
rect 262588 103436 262640 103488
rect 262772 103436 262824 103488
rect 266820 103479 266872 103488
rect 266820 103445 266829 103479
rect 266829 103445 266863 103479
rect 266863 103445 266872 103479
rect 266820 103436 266872 103445
rect 267924 103479 267976 103488
rect 267924 103445 267933 103479
rect 267933 103445 267967 103479
rect 267967 103445 267976 103479
rect 267924 103436 267976 103445
rect 290004 103436 290056 103488
rect 295616 103479 295668 103488
rect 295616 103445 295625 103479
rect 295625 103445 295659 103479
rect 295659 103445 295668 103479
rect 295616 103436 295668 103445
rect 301228 103436 301280 103488
rect 306840 103479 306892 103488
rect 306840 103445 306849 103479
rect 306849 103445 306883 103479
rect 306883 103445 306892 103479
rect 306840 103436 306892 103445
rect 324688 103436 324740 103488
rect 330116 103436 330168 103488
rect 330208 103436 330260 103488
rect 290096 103368 290148 103420
rect 296904 103368 296956 103420
rect 297088 103368 297140 103420
rect 294328 102187 294380 102196
rect 294328 102153 294337 102187
rect 294337 102153 294371 102187
rect 294371 102153 294380 102187
rect 294328 102144 294380 102153
rect 262772 102119 262824 102128
rect 262772 102085 262781 102119
rect 262781 102085 262815 102119
rect 262815 102085 262824 102119
rect 262772 102076 262824 102085
rect 291660 102119 291712 102128
rect 291660 102085 291669 102119
rect 291669 102085 291703 102119
rect 291703 102085 291712 102119
rect 291660 102076 291712 102085
rect 330208 102076 330260 102128
rect 270684 101371 270736 101380
rect 270684 101337 270693 101371
rect 270693 101337 270727 101371
rect 270727 101337 270736 101371
rect 270684 101328 270736 101337
rect 337108 99424 337160 99476
rect 460112 99424 460164 99476
rect 244372 99356 244424 99408
rect 377036 99356 377088 99408
rect 244464 99288 244516 99340
rect 337108 99288 337160 99340
rect 375564 99288 375616 99340
rect 375748 99288 375800 99340
rect 377128 99288 377180 99340
rect 386512 99331 386564 99340
rect 386512 99297 386521 99331
rect 386521 99297 386555 99331
rect 386555 99297 386564 99331
rect 386512 99288 386564 99297
rect 460112 99288 460164 99340
rect 463700 98948 463752 99000
rect 463884 98948 463936 99000
rect 310888 96772 310940 96824
rect 247132 96636 247184 96688
rect 247224 96636 247276 96688
rect 250076 96636 250128 96688
rect 250168 96636 250220 96688
rect 251456 96679 251508 96688
rect 251456 96645 251465 96679
rect 251465 96645 251499 96679
rect 251499 96645 251508 96679
rect 251456 96636 251508 96645
rect 310796 96636 310848 96688
rect 270684 96568 270736 96620
rect 270868 96568 270920 96620
rect 360292 96611 360344 96620
rect 360292 96577 360301 96611
rect 360301 96577 360335 96611
rect 360335 96577 360344 96611
rect 360292 96568 360344 96577
rect 367008 96611 367060 96620
rect 367008 96577 367017 96611
rect 367017 96577 367051 96611
rect 367051 96577 367060 96611
rect 367008 96568 367060 96577
rect 375380 96568 375432 96620
rect 375564 96568 375616 96620
rect 470600 96611 470652 96620
rect 470600 96577 470609 96611
rect 470609 96577 470643 96611
rect 470643 96577 470652 96611
rect 470600 96568 470652 96577
rect 266820 96475 266872 96484
rect 266820 96441 266829 96475
rect 266829 96441 266863 96475
rect 266863 96441 266872 96475
rect 266820 96432 266872 96441
rect 273536 95276 273588 95328
rect 273628 95276 273680 95328
rect 232320 95251 232372 95260
rect 232320 95217 232329 95251
rect 232329 95217 232363 95251
rect 232363 95217 232372 95251
rect 232320 95208 232372 95217
rect 339960 95208 340012 95260
rect 341156 95251 341208 95260
rect 341156 95217 341165 95251
rect 341165 95217 341199 95251
rect 341199 95217 341208 95251
rect 341156 95208 341208 95217
rect 247132 95183 247184 95192
rect 247132 95149 247141 95183
rect 247141 95149 247175 95183
rect 247175 95149 247184 95183
rect 247132 95140 247184 95149
rect 284668 95140 284720 95192
rect 310796 95183 310848 95192
rect 310796 95149 310805 95183
rect 310805 95149 310839 95183
rect 310839 95149 310848 95183
rect 310796 95140 310848 95149
rect 284760 95072 284812 95124
rect 317972 93916 318024 93968
rect 265164 93848 265216 93900
rect 265256 93848 265308 93900
rect 267740 93848 267792 93900
rect 295616 93891 295668 93900
rect 295616 93857 295625 93891
rect 295625 93857 295659 93891
rect 295659 93857 295668 93891
rect 295616 93848 295668 93857
rect 301136 93891 301188 93900
rect 301136 93857 301145 93891
rect 301145 93857 301179 93891
rect 301179 93857 301188 93891
rect 301136 93848 301188 93857
rect 306840 93891 306892 93900
rect 306840 93857 306849 93891
rect 306849 93857 306883 93891
rect 306883 93857 306892 93891
rect 306840 93848 306892 93857
rect 317696 93848 317748 93900
rect 324596 93891 324648 93900
rect 324596 93857 324605 93891
rect 324605 93857 324639 93891
rect 324639 93857 324648 93891
rect 324596 93848 324648 93857
rect 262772 92531 262824 92540
rect 262772 92497 262781 92531
rect 262781 92497 262815 92531
rect 262815 92497 262824 92531
rect 262772 92488 262824 92497
rect 291660 92531 291712 92540
rect 291660 92497 291669 92531
rect 291669 92497 291703 92531
rect 291703 92497 291712 92531
rect 291660 92488 291712 92497
rect 341156 90380 341208 90432
rect 386420 89700 386472 89752
rect 386604 89700 386656 89752
rect 360292 89675 360344 89684
rect 360292 89641 360301 89675
rect 360301 89641 360335 89675
rect 360335 89641 360344 89675
rect 360292 89632 360344 89641
rect 262772 88952 262824 89004
rect 265164 88995 265216 89004
rect 265164 88961 265173 88995
rect 265173 88961 265207 88995
rect 265207 88961 265216 88995
rect 265164 88952 265216 88961
rect 317696 88383 317748 88392
rect 317696 88349 317705 88383
rect 317705 88349 317739 88383
rect 317739 88349 317748 88383
rect 317696 88340 317748 88349
rect 454040 87252 454092 87304
rect 456984 87252 457036 87304
rect 437204 87116 437256 87168
rect 437480 87116 437532 87168
rect 494612 87116 494664 87168
rect 502248 87116 502300 87168
rect 251180 87048 251232 87100
rect 260656 87048 260708 87100
rect 347780 86980 347832 87032
rect 357348 86980 357400 87032
rect 367008 87023 367060 87032
rect 367008 86989 367017 87023
rect 367017 86989 367051 87023
rect 367051 86989 367060 87023
rect 367008 86980 367060 86989
rect 421196 87023 421248 87032
rect 421196 86989 421205 87023
rect 421205 86989 421239 87023
rect 421239 86989 421248 87023
rect 421196 86980 421248 86989
rect 470600 87023 470652 87032
rect 470600 86989 470609 87023
rect 470609 86989 470643 87023
rect 470643 86989 470652 87023
rect 470600 86980 470652 86989
rect 236460 86912 236512 86964
rect 251456 86955 251508 86964
rect 251456 86921 251465 86955
rect 251465 86921 251499 86955
rect 251499 86921 251508 86955
rect 251456 86912 251508 86921
rect 323308 86912 323360 86964
rect 323400 86912 323452 86964
rect 324596 86912 324648 86964
rect 325884 86912 325936 86964
rect 327172 86912 327224 86964
rect 327264 86912 327316 86964
rect 336924 86955 336976 86964
rect 336924 86921 336933 86955
rect 336933 86921 336967 86955
rect 336967 86921 336976 86955
rect 336924 86912 336976 86921
rect 337200 86955 337252 86964
rect 337200 86921 337209 86955
rect 337209 86921 337243 86955
rect 337243 86921 337252 86955
rect 337200 86912 337252 86921
rect 324688 86844 324740 86896
rect 325976 86844 326028 86896
rect 360200 86844 360252 86896
rect 360384 86844 360436 86896
rect 375564 86844 375616 86896
rect 375656 86844 375708 86896
rect 286232 85620 286284 85672
rect 247224 85552 247276 85604
rect 285956 85552 286008 85604
rect 291660 85552 291712 85604
rect 294236 85552 294288 85604
rect 294328 85552 294380 85604
rect 310796 85595 310848 85604
rect 310796 85561 310805 85595
rect 310805 85561 310839 85595
rect 310839 85561 310848 85595
rect 310796 85552 310848 85561
rect 232320 85527 232372 85536
rect 232320 85493 232329 85527
rect 232329 85493 232363 85527
rect 232363 85493 232372 85527
rect 232320 85484 232372 85493
rect 267740 85484 267792 85536
rect 267832 85484 267884 85536
rect 273536 85484 273588 85536
rect 273628 85484 273680 85536
rect 299848 85527 299900 85536
rect 299848 85493 299857 85527
rect 299857 85493 299891 85527
rect 299891 85493 299900 85527
rect 299848 85484 299900 85493
rect 301044 85484 301096 85536
rect 301228 85484 301280 85536
rect 306656 85484 306708 85536
rect 306840 85484 306892 85536
rect 324688 85527 324740 85536
rect 324688 85493 324697 85527
rect 324697 85493 324731 85527
rect 324731 85493 324740 85527
rect 324688 85484 324740 85493
rect 358728 85527 358780 85536
rect 358728 85493 358737 85527
rect 358737 85493 358771 85527
rect 358771 85493 358780 85527
rect 358728 85484 358780 85493
rect 421196 85527 421248 85536
rect 421196 85493 421205 85527
rect 421205 85493 421239 85527
rect 421239 85493 421248 85527
rect 421196 85484 421248 85493
rect 296996 84260 297048 84312
rect 291568 84235 291620 84244
rect 291568 84201 291577 84235
rect 291577 84201 291611 84235
rect 291611 84201 291620 84235
rect 291568 84192 291620 84201
rect 297088 84192 297140 84244
rect 272340 84124 272392 84176
rect 284760 84124 284812 84176
rect 285956 84167 286008 84176
rect 285956 84133 285965 84167
rect 285965 84133 285999 84167
rect 285999 84133 286008 84167
rect 285956 84124 286008 84133
rect 288716 82807 288768 82816
rect 288716 82773 288725 82807
rect 288725 82773 288759 82807
rect 288759 82773 288768 82807
rect 288716 82764 288768 82773
rect 270776 80767 270828 80776
rect 270776 80733 270785 80767
rect 270785 80733 270819 80767
rect 270819 80733 270828 80767
rect 270776 80724 270828 80733
rect 357716 80112 357768 80164
rect 359188 80112 359240 80164
rect 372804 80112 372856 80164
rect 303896 80044 303948 80096
rect 357624 80044 357676 80096
rect 359096 80044 359148 80096
rect 372712 80044 372764 80096
rect 303896 79908 303948 79960
rect 2780 79772 2832 79824
rect 4896 79772 4948 79824
rect 236276 77435 236328 77444
rect 236276 77401 236285 77435
rect 236285 77401 236319 77435
rect 236319 77401 236328 77435
rect 236276 77392 236328 77401
rect 358820 77324 358872 77376
rect 358912 77324 358964 77376
rect 251456 77299 251508 77308
rect 251456 77265 251465 77299
rect 251465 77265 251499 77299
rect 251499 77265 251508 77299
rect 251456 77256 251508 77265
rect 330208 77256 330260 77308
rect 337200 77299 337252 77308
rect 337200 77265 337209 77299
rect 337209 77265 337243 77299
rect 337243 77265 337252 77299
rect 337200 77256 337252 77265
rect 339776 77256 339828 77308
rect 339960 77256 340012 77308
rect 341064 77299 341116 77308
rect 341064 77265 341073 77299
rect 341073 77265 341107 77299
rect 341107 77265 341116 77299
rect 341064 77256 341116 77265
rect 303896 77188 303948 77240
rect 303988 77188 304040 77240
rect 358820 77188 358872 77240
rect 358912 77188 358964 77240
rect 386696 77188 386748 77240
rect 470600 77231 470652 77240
rect 470600 77197 470609 77231
rect 470609 77197 470643 77231
rect 470643 77197 470652 77231
rect 470600 77188 470652 77197
rect 310796 76100 310848 76152
rect 328920 76100 328972 76152
rect 338028 76100 338080 76152
rect 369860 76100 369912 76152
rect 376668 76100 376720 76152
rect 396080 76032 396132 76084
rect 399392 76032 399444 76084
rect 414020 76032 414072 76084
rect 423404 76032 423456 76084
rect 437204 76032 437256 76084
rect 437480 76032 437532 76084
rect 310796 75964 310848 76016
rect 324688 76007 324740 76016
rect 324688 75973 324697 76007
rect 324697 75973 324731 76007
rect 324731 75973 324740 76007
rect 324688 75964 324740 75973
rect 232320 75939 232372 75948
rect 232320 75905 232329 75939
rect 232329 75905 232363 75939
rect 232363 75905 232372 75939
rect 232320 75896 232372 75905
rect 262680 75939 262732 75948
rect 262680 75905 262689 75939
rect 262689 75905 262723 75939
rect 262723 75905 262732 75939
rect 262680 75896 262732 75905
rect 289912 75896 289964 75948
rect 290096 75896 290148 75948
rect 291384 75896 291436 75948
rect 291568 75896 291620 75948
rect 295524 75896 295576 75948
rect 295708 75896 295760 75948
rect 299848 75939 299900 75948
rect 299848 75905 299857 75939
rect 299857 75905 299891 75939
rect 299891 75905 299900 75939
rect 299848 75896 299900 75905
rect 302516 75896 302568 75948
rect 302608 75896 302660 75948
rect 317696 75939 317748 75948
rect 317696 75905 317705 75939
rect 317705 75905 317739 75939
rect 317739 75905 317748 75939
rect 317696 75896 317748 75905
rect 336924 75939 336976 75948
rect 336924 75905 336933 75939
rect 336933 75905 336967 75939
rect 336967 75905 336976 75939
rect 336924 75896 336976 75905
rect 359004 75896 359056 75948
rect 421196 75939 421248 75948
rect 421196 75905 421205 75939
rect 421205 75905 421239 75939
rect 421239 75905 421248 75939
rect 421196 75896 421248 75905
rect 310796 75871 310848 75880
rect 310796 75837 310805 75871
rect 310805 75837 310839 75871
rect 310839 75837 310848 75871
rect 310796 75828 310848 75837
rect 324688 75828 324740 75880
rect 296812 74604 296864 74656
rect 297088 74604 297140 74656
rect 265440 74536 265492 74588
rect 272248 74579 272300 74588
rect 272248 74545 272257 74579
rect 272257 74545 272291 74579
rect 272291 74545 272300 74579
rect 272248 74536 272300 74545
rect 239128 70499 239180 70508
rect 239128 70465 239137 70499
rect 239137 70465 239171 70499
rect 239171 70465 239180 70499
rect 239128 70456 239180 70465
rect 244464 70499 244516 70508
rect 244464 70465 244473 70499
rect 244473 70465 244507 70499
rect 244507 70465 244516 70499
rect 244464 70456 244516 70465
rect 377128 70499 377180 70508
rect 377128 70465 377137 70499
rect 377137 70465 377171 70499
rect 377171 70465 377180 70499
rect 377128 70456 377180 70465
rect 367008 67736 367060 67788
rect 272248 67711 272300 67720
rect 272248 67677 272257 67711
rect 272257 67677 272291 67711
rect 272291 67677 272300 67711
rect 272248 67668 272300 67677
rect 323308 67668 323360 67720
rect 239128 67643 239180 67652
rect 239128 67609 239137 67643
rect 239137 67609 239171 67643
rect 239171 67609 239180 67643
rect 239128 67600 239180 67609
rect 244464 67643 244516 67652
rect 244464 67609 244473 67643
rect 244473 67609 244507 67643
rect 244507 67609 244516 67643
rect 244464 67600 244516 67609
rect 270776 67643 270828 67652
rect 270776 67609 270785 67643
rect 270785 67609 270819 67643
rect 270819 67609 270828 67643
rect 270776 67600 270828 67609
rect 299756 67600 299808 67652
rect 299848 67600 299900 67652
rect 323400 67600 323452 67652
rect 341064 67600 341116 67652
rect 341156 67600 341208 67652
rect 358728 67600 358780 67652
rect 359004 67600 359056 67652
rect 367008 67600 367060 67652
rect 377128 67643 377180 67652
rect 377128 67609 377137 67643
rect 377137 67609 377171 67643
rect 377171 67609 377180 67643
rect 377128 67600 377180 67609
rect 386604 67643 386656 67652
rect 386604 67609 386613 67643
rect 386613 67609 386647 67643
rect 386647 67609 386656 67643
rect 386604 67600 386656 67609
rect 470600 67643 470652 67652
rect 470600 67609 470609 67643
rect 470609 67609 470643 67643
rect 470643 67609 470652 67643
rect 470600 67600 470652 67609
rect 236276 67532 236328 67584
rect 236368 67532 236420 67584
rect 250076 67575 250128 67584
rect 250076 67541 250085 67575
rect 250085 67541 250119 67575
rect 250119 67541 250128 67575
rect 250076 67532 250128 67541
rect 375656 67575 375708 67584
rect 375656 67541 375665 67575
rect 375665 67541 375699 67575
rect 375699 67541 375708 67575
rect 375656 67532 375708 67541
rect 459928 67532 459980 67584
rect 460204 67532 460256 67584
rect 272248 67099 272300 67108
rect 272248 67065 272257 67099
rect 272257 67065 272291 67099
rect 272291 67065 272300 67099
rect 272248 67056 272300 67065
rect 310796 66351 310848 66360
rect 310796 66317 310805 66351
rect 310805 66317 310839 66351
rect 310839 66317 310848 66351
rect 310796 66308 310848 66317
rect 324596 66351 324648 66360
rect 324596 66317 324605 66351
rect 324605 66317 324639 66351
rect 324639 66317 324648 66351
rect 324596 66308 324648 66317
rect 267740 66240 267792 66292
rect 267832 66240 267884 66292
rect 284668 66283 284720 66292
rect 284668 66249 284677 66283
rect 284677 66249 284711 66283
rect 284711 66249 284720 66283
rect 284668 66240 284720 66249
rect 285956 66283 286008 66292
rect 285956 66249 285965 66283
rect 285965 66249 285999 66283
rect 285999 66249 286008 66283
rect 285956 66240 286008 66249
rect 296812 66240 296864 66292
rect 327264 66240 327316 66292
rect 232320 66215 232372 66224
rect 232320 66181 232329 66215
rect 232329 66181 232363 66215
rect 232363 66181 232372 66215
rect 232320 66172 232372 66181
rect 236368 66172 236420 66224
rect 270776 66215 270828 66224
rect 270776 66181 270785 66215
rect 270785 66181 270819 66215
rect 270819 66181 270828 66215
rect 270776 66172 270828 66181
rect 273444 66215 273496 66224
rect 273444 66181 273453 66215
rect 273453 66181 273487 66215
rect 273487 66181 273496 66215
rect 273444 66172 273496 66181
rect 310796 66215 310848 66224
rect 310796 66181 310805 66215
rect 310805 66181 310839 66215
rect 310839 66181 310848 66215
rect 310796 66172 310848 66181
rect 323400 66172 323452 66224
rect 324596 66215 324648 66224
rect 324596 66181 324605 66215
rect 324605 66181 324639 66215
rect 324639 66181 324648 66215
rect 324596 66172 324648 66181
rect 296904 66104 296956 66156
rect 330116 66215 330168 66224
rect 330116 66181 330125 66215
rect 330125 66181 330159 66215
rect 330159 66181 330168 66215
rect 330116 66172 330168 66181
rect 336924 66215 336976 66224
rect 336924 66181 336933 66215
rect 336933 66181 336967 66215
rect 336967 66181 336976 66215
rect 336924 66172 336976 66181
rect 358728 66172 358780 66224
rect 367008 66215 367060 66224
rect 367008 66181 367017 66215
rect 367017 66181 367051 66215
rect 367051 66181 367060 66215
rect 367008 66172 367060 66181
rect 421196 66215 421248 66224
rect 421196 66181 421205 66215
rect 421205 66181 421239 66215
rect 421239 66181 421248 66215
rect 421196 66172 421248 66181
rect 327356 66104 327408 66156
rect 306656 65764 306708 65816
rect 306840 65764 306892 65816
rect 288900 64880 288952 64932
rect 3332 64812 3384 64864
rect 24124 64812 24176 64864
rect 294236 64855 294288 64864
rect 294236 64821 294245 64855
rect 294245 64821 294279 64855
rect 294279 64821 294288 64855
rect 294236 64812 294288 64821
rect 378508 63860 378560 63912
rect 386328 63860 386380 63912
rect 367100 63724 367152 63776
rect 376668 63724 376720 63776
rect 417884 63656 417936 63708
rect 418160 63656 418212 63708
rect 437204 63656 437256 63708
rect 437480 63656 437532 63708
rect 456524 63656 456576 63708
rect 456892 63656 456944 63708
rect 262588 62772 262640 62824
rect 262772 62772 262824 62824
rect 259736 62636 259788 62688
rect 265348 62636 265400 62688
rect 259920 62568 259972 62620
rect 375656 61999 375708 62008
rect 375656 61965 375665 61999
rect 375665 61965 375699 61999
rect 375699 61965 375708 61999
rect 375656 61956 375708 61965
rect 324688 61344 324740 61396
rect 339684 60664 339736 60716
rect 339868 60664 339920 60716
rect 341156 60664 341208 60716
rect 341340 60664 341392 60716
rect 360292 60664 360344 60716
rect 360476 60664 360528 60716
rect 310888 59984 310940 60036
rect 239128 58012 239180 58064
rect 244464 57944 244516 57996
rect 250168 57944 250220 57996
rect 266728 57944 266780 57996
rect 266820 57944 266872 57996
rect 267740 57944 267792 57996
rect 267832 57944 267884 57996
rect 284668 57944 284720 57996
rect 284760 57944 284812 57996
rect 285956 57944 286008 57996
rect 286048 57944 286100 57996
rect 291476 58012 291528 58064
rect 303896 57944 303948 57996
rect 303988 57944 304040 57996
rect 265164 57919 265216 57928
rect 265164 57885 265173 57919
rect 265173 57885 265207 57919
rect 265207 57885 265216 57919
rect 265164 57876 265216 57885
rect 291384 57876 291436 57928
rect 339868 57876 339920 57928
rect 460112 57876 460164 57928
rect 470600 57919 470652 57928
rect 470600 57885 470609 57919
rect 470609 57885 470643 57919
rect 470643 57885 470652 57919
rect 470600 57876 470652 57885
rect 244556 57808 244608 57860
rect 301044 56652 301096 56704
rect 301228 56652 301280 56704
rect 232320 56627 232372 56636
rect 232320 56593 232329 56627
rect 232329 56593 232363 56627
rect 232363 56593 232372 56627
rect 232320 56584 232372 56593
rect 236276 56627 236328 56636
rect 236276 56593 236285 56627
rect 236285 56593 236319 56627
rect 236319 56593 236328 56627
rect 236276 56584 236328 56593
rect 239036 56627 239088 56636
rect 239036 56593 239045 56627
rect 239045 56593 239079 56627
rect 239079 56593 239088 56627
rect 239036 56584 239088 56593
rect 270776 56627 270828 56636
rect 270776 56593 270785 56627
rect 270785 56593 270819 56627
rect 270819 56593 270828 56627
rect 270776 56584 270828 56593
rect 330208 56584 330260 56636
rect 336924 56627 336976 56636
rect 336924 56593 336933 56627
rect 336933 56593 336967 56627
rect 336967 56593 336976 56627
rect 336924 56584 336976 56593
rect 357532 56584 357584 56636
rect 357716 56584 357768 56636
rect 358636 56627 358688 56636
rect 358636 56593 358645 56627
rect 358645 56593 358679 56627
rect 358679 56593 358688 56627
rect 358636 56584 358688 56593
rect 421196 56627 421248 56636
rect 421196 56593 421205 56627
rect 421205 56593 421239 56627
rect 421239 56593 421248 56627
rect 421196 56584 421248 56593
rect 244556 56559 244608 56568
rect 244556 56525 244565 56559
rect 244565 56525 244599 56559
rect 244599 56525 244608 56559
rect 244556 56516 244608 56525
rect 299664 56559 299716 56568
rect 299664 56525 299673 56559
rect 299673 56525 299707 56559
rect 299707 56525 299716 56559
rect 299664 56516 299716 56525
rect 301044 56559 301096 56568
rect 301044 56525 301053 56559
rect 301053 56525 301087 56559
rect 301087 56525 301096 56559
rect 301044 56516 301096 56525
rect 324780 56559 324832 56568
rect 324780 56525 324789 56559
rect 324789 56525 324823 56559
rect 324823 56525 324832 56559
rect 324780 56516 324832 56525
rect 337292 56559 337344 56568
rect 337292 56525 337301 56559
rect 337301 56525 337335 56559
rect 337335 56525 337344 56559
rect 337292 56516 337344 56525
rect 357532 56491 357584 56500
rect 357532 56457 357541 56491
rect 357541 56457 357575 56491
rect 357575 56457 357584 56491
rect 357532 56448 357584 56457
rect 288716 55292 288768 55344
rect 288900 55224 288952 55276
rect 317512 55224 317564 55276
rect 317696 55224 317748 55276
rect 310888 55156 310940 55208
rect 311072 55156 311124 55208
rect 239036 53184 239088 53236
rect 265164 53116 265216 53168
rect 265348 53116 265400 53168
rect 247224 51076 247276 51128
rect 247132 51008 247184 51060
rect 386420 51008 386472 51060
rect 386604 51008 386656 51060
rect 273536 50940 273588 50992
rect 2780 50464 2832 50516
rect 4804 50464 4856 50516
rect 286048 48356 286100 48408
rect 360476 48356 360528 48408
rect 239128 48331 239180 48340
rect 239128 48297 239137 48331
rect 239137 48297 239171 48331
rect 239171 48297 239180 48331
rect 239128 48288 239180 48297
rect 267832 48288 267884 48340
rect 236276 48263 236328 48272
rect 236276 48229 236285 48263
rect 236285 48229 236319 48263
rect 236319 48229 236328 48263
rect 236276 48220 236328 48229
rect 250168 48220 250220 48272
rect 250260 48220 250312 48272
rect 284668 48288 284720 48340
rect 284760 48288 284812 48340
rect 285956 48288 286008 48340
rect 323308 48331 323360 48340
rect 323308 48297 323317 48331
rect 323317 48297 323351 48331
rect 323351 48297 323360 48331
rect 323308 48288 323360 48297
rect 339776 48331 339828 48340
rect 339776 48297 339785 48331
rect 339785 48297 339819 48331
rect 339819 48297 339828 48331
rect 339776 48288 339828 48297
rect 341248 48288 341300 48340
rect 341432 48288 341484 48340
rect 358636 48288 358688 48340
rect 358728 48288 358780 48340
rect 360384 48288 360436 48340
rect 367008 48331 367060 48340
rect 367008 48297 367017 48331
rect 367017 48297 367051 48331
rect 367051 48297 367060 48331
rect 367008 48288 367060 48297
rect 460020 48331 460072 48340
rect 460020 48297 460029 48331
rect 460029 48297 460063 48331
rect 460063 48297 460072 48331
rect 460020 48288 460072 48297
rect 470600 48331 470652 48340
rect 470600 48297 470609 48331
rect 470609 48297 470643 48331
rect 470643 48297 470652 48331
rect 470600 48288 470652 48297
rect 273536 48263 273588 48272
rect 273536 48229 273545 48263
rect 273545 48229 273579 48263
rect 273579 48229 273588 48263
rect 273536 48220 273588 48229
rect 244556 48195 244608 48204
rect 244556 48161 244565 48195
rect 244565 48161 244599 48195
rect 244599 48161 244608 48195
rect 244556 48152 244608 48161
rect 267924 48152 267976 48204
rect 460020 48195 460072 48204
rect 460020 48161 460029 48195
rect 460029 48161 460063 48195
rect 460063 48161 460072 48195
rect 460020 48152 460072 48161
rect 291384 46996 291436 47048
rect 337200 46996 337252 47048
rect 266544 46928 266596 46980
rect 266728 46928 266780 46980
rect 288716 46928 288768 46980
rect 288900 46928 288952 46980
rect 291476 46928 291528 46980
rect 294236 46971 294288 46980
rect 294236 46937 294245 46971
rect 294245 46937 294279 46971
rect 294279 46937 294288 46971
rect 294236 46928 294288 46937
rect 301044 46971 301096 46980
rect 301044 46937 301053 46971
rect 301053 46937 301087 46971
rect 301087 46937 301096 46971
rect 301044 46928 301096 46937
rect 303804 46928 303856 46980
rect 303896 46928 303948 46980
rect 306748 46928 306800 46980
rect 306840 46928 306892 46980
rect 324596 46928 324648 46980
rect 357624 46928 357676 46980
rect 377220 46928 377272 46980
rect 377312 46928 377364 46980
rect 244556 46903 244608 46912
rect 244556 46869 244565 46903
rect 244565 46869 244599 46903
rect 244599 46869 244608 46903
rect 244556 46860 244608 46869
rect 262588 46860 262640 46912
rect 262772 46860 262824 46912
rect 323308 46903 323360 46912
rect 323308 46869 323317 46903
rect 323317 46869 323351 46903
rect 323351 46869 323360 46903
rect 323308 46860 323360 46869
rect 327264 46903 327316 46912
rect 327264 46869 327273 46903
rect 327273 46869 327307 46903
rect 327307 46869 327316 46903
rect 327264 46860 327316 46869
rect 330116 46903 330168 46912
rect 330116 46869 330125 46903
rect 330125 46869 330159 46903
rect 330159 46869 330168 46903
rect 330116 46860 330168 46869
rect 336924 46903 336976 46912
rect 336924 46869 336933 46903
rect 336933 46869 336967 46903
rect 336967 46869 336976 46903
rect 336924 46860 336976 46869
rect 337200 46903 337252 46912
rect 337200 46869 337209 46903
rect 337209 46869 337243 46903
rect 337243 46869 337252 46903
rect 337200 46860 337252 46869
rect 341432 46860 341484 46912
rect 358728 46860 358780 46912
rect 359096 46860 359148 46912
rect 367008 46903 367060 46912
rect 367008 46869 367017 46903
rect 367017 46869 367051 46903
rect 367051 46869 367060 46903
rect 367008 46860 367060 46869
rect 421196 46903 421248 46912
rect 421196 46869 421205 46903
rect 421205 46869 421239 46903
rect 421239 46869 421248 46903
rect 421196 46860 421248 46869
rect 357624 46835 357676 46844
rect 357624 46801 357633 46835
rect 357633 46801 357667 46835
rect 357667 46801 357676 46835
rect 357624 46792 357676 46801
rect 299756 45568 299808 45620
rect 262772 45543 262824 45552
rect 262772 45509 262781 45543
rect 262781 45509 262815 45543
rect 262815 45509 262824 45543
rect 262772 45500 262824 45509
rect 294236 45543 294288 45552
rect 294236 45509 294245 45543
rect 294245 45509 294279 45543
rect 294279 45509 294288 45543
rect 294236 45500 294288 45509
rect 310888 45500 310940 45552
rect 311072 45500 311124 45552
rect 317512 45500 317564 45552
rect 317696 45500 317748 45552
rect 299756 45432 299808 45484
rect 299848 45432 299900 45484
rect 284668 44684 284720 44736
rect 239128 42032 239180 42084
rect 360292 41352 360344 41404
rect 360476 41352 360528 41404
rect 460204 41352 460256 41404
rect 367100 40196 367152 40248
rect 376668 40196 376720 40248
rect 417884 40196 417936 40248
rect 420368 40196 420420 40248
rect 437204 40196 437256 40248
rect 437480 40196 437532 40248
rect 456524 40196 456576 40248
rect 456892 40196 456944 40248
rect 306380 40128 306432 40180
rect 315948 40128 316000 40180
rect 232320 38632 232372 38684
rect 236276 38675 236328 38684
rect 236276 38641 236285 38675
rect 236285 38641 236319 38675
rect 236319 38641 236328 38675
rect 236276 38632 236328 38641
rect 247132 38632 247184 38684
rect 247224 38632 247276 38684
rect 270776 38632 270828 38684
rect 270868 38632 270920 38684
rect 272156 38632 272208 38684
rect 272248 38632 272300 38684
rect 273536 38675 273588 38684
rect 273536 38641 273545 38675
rect 273545 38641 273579 38675
rect 273579 38641 273588 38675
rect 273536 38632 273588 38641
rect 296812 38632 296864 38684
rect 301044 38632 301096 38684
rect 302516 38632 302568 38684
rect 302608 38632 302660 38684
rect 232504 38496 232556 38548
rect 236276 38539 236328 38548
rect 236276 38505 236285 38539
rect 236285 38505 236319 38539
rect 236319 38505 236328 38539
rect 236276 38496 236328 38505
rect 301320 38564 301372 38616
rect 303804 38607 303856 38616
rect 303804 38573 303813 38607
rect 303813 38573 303847 38607
rect 303847 38573 303856 38607
rect 303804 38564 303856 38573
rect 306748 38564 306800 38616
rect 306840 38564 306892 38616
rect 377128 38564 377180 38616
rect 377312 38564 377364 38616
rect 296904 38496 296956 38548
rect 250260 38156 250312 38208
rect 250260 38020 250312 38072
rect 337200 37383 337252 37392
rect 337200 37349 337209 37383
rect 337209 37349 337243 37383
rect 337243 37349 337252 37383
rect 337200 37340 337252 37349
rect 244556 37315 244608 37324
rect 244556 37281 244565 37315
rect 244565 37281 244599 37315
rect 244599 37281 244608 37315
rect 244556 37272 244608 37281
rect 266544 37272 266596 37324
rect 266636 37272 266688 37324
rect 323400 37272 323452 37324
rect 327264 37315 327316 37324
rect 327264 37281 327273 37315
rect 327273 37281 327307 37315
rect 327307 37281 327316 37315
rect 327264 37272 327316 37281
rect 330116 37315 330168 37324
rect 330116 37281 330125 37315
rect 330125 37281 330159 37315
rect 330159 37281 330168 37315
rect 330116 37272 330168 37281
rect 336924 37315 336976 37324
rect 336924 37281 336933 37315
rect 336933 37281 336967 37315
rect 336967 37281 336976 37315
rect 336924 37272 336976 37281
rect 341248 37315 341300 37324
rect 341248 37281 341257 37315
rect 341257 37281 341291 37315
rect 341291 37281 341300 37315
rect 341248 37272 341300 37281
rect 357624 37315 357676 37324
rect 357624 37281 357633 37315
rect 357633 37281 357667 37315
rect 357667 37281 357676 37315
rect 357624 37272 357676 37281
rect 358636 37315 358688 37324
rect 358636 37281 358645 37315
rect 358645 37281 358679 37315
rect 358679 37281 358688 37315
rect 358636 37272 358688 37281
rect 359004 37315 359056 37324
rect 359004 37281 359013 37315
rect 359013 37281 359047 37315
rect 359047 37281 359056 37315
rect 359004 37272 359056 37281
rect 367008 37315 367060 37324
rect 367008 37281 367017 37315
rect 367017 37281 367051 37315
rect 367051 37281 367060 37315
rect 367008 37272 367060 37281
rect 421196 37315 421248 37324
rect 421196 37281 421205 37315
rect 421205 37281 421239 37315
rect 421239 37281 421248 37315
rect 421196 37272 421248 37281
rect 251180 37204 251232 37256
rect 251456 37204 251508 37256
rect 259736 37247 259788 37256
rect 259736 37213 259745 37247
rect 259745 37213 259779 37247
rect 259779 37213 259788 37247
rect 259736 37204 259788 37213
rect 267924 37204 267976 37256
rect 272248 37204 272300 37256
rect 272340 37204 272392 37256
rect 288716 37204 288768 37256
rect 337200 37204 337252 37256
rect 337292 37204 337344 37256
rect 288808 37136 288860 37188
rect 262772 35955 262824 35964
rect 262772 35921 262781 35955
rect 262781 35921 262815 35955
rect 262815 35921 262824 35955
rect 262772 35912 262824 35921
rect 3148 35844 3200 35896
rect 6184 35844 6236 35896
rect 272340 35844 272392 35896
rect 301320 35844 301372 35896
rect 311072 35844 311124 35896
rect 359004 34076 359056 34128
rect 359096 34008 359148 34060
rect 336740 33804 336792 33856
rect 336924 33804 336976 33856
rect 303896 32376 303948 32428
rect 357624 32376 357676 32428
rect 357808 32376 357860 32428
rect 341248 32283 341300 32292
rect 341248 32249 341257 32283
rect 341257 32249 341291 32283
rect 341291 32249 341300 32283
rect 341248 32240 341300 32249
rect 317512 31764 317564 31816
rect 317696 31764 317748 31816
rect 327264 31764 327316 31816
rect 377128 31764 377180 31816
rect 386512 31764 386564 31816
rect 236368 31628 236420 31680
rect 377128 31628 377180 31680
rect 386604 31628 386656 31680
rect 327264 31560 327316 31612
rect 278780 29248 278832 29300
rect 281264 29248 281316 29300
rect 367100 29180 367152 29232
rect 376668 29180 376720 29232
rect 240140 29112 240192 29164
rect 249708 29112 249760 29164
rect 367008 29112 367060 29164
rect 437204 29112 437256 29164
rect 437480 29112 437532 29164
rect 456524 29112 456576 29164
rect 456800 29112 456852 29164
rect 302516 29044 302568 29096
rect 341248 29087 341300 29096
rect 341248 29053 341257 29087
rect 341257 29053 341291 29087
rect 341291 29053 341300 29087
rect 341248 29044 341300 29053
rect 347780 29044 347832 29096
rect 357348 29044 357400 29096
rect 239036 29019 239088 29028
rect 239036 28985 239045 29019
rect 239045 28985 239079 29019
rect 239079 28985 239088 29019
rect 239036 28976 239088 28985
rect 284760 29019 284812 29028
rect 284760 28985 284769 29019
rect 284769 28985 284803 29019
rect 284803 28985 284812 29019
rect 284760 28976 284812 28985
rect 285956 28976 286008 29028
rect 286048 28976 286100 29028
rect 492772 29044 492824 29096
rect 502248 29044 502300 29096
rect 325976 28976 326028 29028
rect 326068 28976 326120 29028
rect 358636 28976 358688 29028
rect 358728 28976 358780 29028
rect 367008 28976 367060 29028
rect 232228 28908 232280 28960
rect 232412 28908 232464 28960
rect 236368 28951 236420 28960
rect 236368 28917 236377 28951
rect 236377 28917 236411 28951
rect 236411 28917 236420 28951
rect 236368 28908 236420 28917
rect 291476 28908 291528 28960
rect 291660 28908 291712 28960
rect 295524 28908 295576 28960
rect 295616 28908 295668 28960
rect 302516 28908 302568 28960
rect 323308 28908 323360 28960
rect 323400 28908 323452 28960
rect 324596 28908 324648 28960
rect 324688 28908 324740 28960
rect 306380 28840 306432 28892
rect 315948 28840 316000 28892
rect 267832 28611 267884 28620
rect 267832 28577 267841 28611
rect 267841 28577 267875 28611
rect 267875 28577 267884 28611
rect 267832 28568 267884 28577
rect 259736 27659 259788 27668
rect 259736 27625 259745 27659
rect 259745 27625 259779 27659
rect 259779 27625 259788 27659
rect 259736 27616 259788 27625
rect 247132 27591 247184 27600
rect 247132 27557 247141 27591
rect 247141 27557 247175 27591
rect 247175 27557 247184 27591
rect 247132 27548 247184 27557
rect 250168 27548 250220 27600
rect 251364 27591 251416 27600
rect 251364 27557 251373 27591
rect 251373 27557 251407 27591
rect 251407 27557 251416 27591
rect 251364 27548 251416 27557
rect 262588 27548 262640 27600
rect 262680 27548 262732 27600
rect 265256 27548 265308 27600
rect 284760 27591 284812 27600
rect 284760 27557 284769 27591
rect 284769 27557 284803 27591
rect 284803 27557 284812 27591
rect 284760 27548 284812 27557
rect 286048 27548 286100 27600
rect 341156 27548 341208 27600
rect 357624 27591 357676 27600
rect 357624 27557 357633 27591
rect 357633 27557 357667 27591
rect 357667 27557 357676 27591
rect 357624 27548 357676 27557
rect 358728 27548 358780 27600
rect 359096 27548 359148 27600
rect 359188 27548 359240 27600
rect 367008 27548 367060 27600
rect 421196 27591 421248 27600
rect 421196 27557 421205 27591
rect 421205 27557 421239 27591
rect 421239 27557 421248 27591
rect 421196 27548 421248 27557
rect 272248 26299 272300 26308
rect 272248 26265 272257 26299
rect 272257 26265 272291 26299
rect 272291 26265 272300 26299
rect 272248 26256 272300 26265
rect 294420 26256 294472 26308
rect 301136 26299 301188 26308
rect 301136 26265 301145 26299
rect 301145 26265 301179 26299
rect 301179 26265 301188 26299
rect 301136 26256 301188 26265
rect 310888 26299 310940 26308
rect 310888 26265 310897 26299
rect 310897 26265 310931 26299
rect 310931 26265 310940 26299
rect 310888 26256 310940 26265
rect 386604 26188 386656 26240
rect 271880 26120 271932 26172
rect 272248 26120 272300 26172
rect 236460 22720 236512 22772
rect 270776 22108 270828 22160
rect 310796 22108 310848 22160
rect 377128 22108 377180 22160
rect 377036 22040 377088 22092
rect 291568 19932 291620 19984
rect 291568 19796 291620 19848
rect 306748 19320 306800 19372
rect 306840 19320 306892 19372
rect 336740 19320 336792 19372
rect 336924 19320 336976 19372
rect 251364 19295 251416 19304
rect 251364 19261 251373 19295
rect 251373 19261 251407 19295
rect 251407 19261 251416 19295
rect 251364 19252 251416 19261
rect 325976 19252 326028 19304
rect 327264 19252 327316 19304
rect 470600 19295 470652 19304
rect 470600 19261 470609 19295
rect 470609 19261 470643 19295
rect 470643 19261 470652 19295
rect 470600 19252 470652 19261
rect 325976 19116 326028 19168
rect 327264 19116 327316 19168
rect 337292 18436 337344 18488
rect 247132 18003 247184 18012
rect 247132 17969 247141 18003
rect 247141 17969 247175 18003
rect 247175 17969 247184 18003
rect 247132 17960 247184 17969
rect 249984 18003 250036 18012
rect 249984 17969 249993 18003
rect 249993 17969 250027 18003
rect 250027 17969 250036 18003
rect 249984 17960 250036 17969
rect 265164 18003 265216 18012
rect 265164 17969 265173 18003
rect 265173 17969 265207 18003
rect 265207 17969 265216 18003
rect 265164 17960 265216 17969
rect 270592 17960 270644 18012
rect 271972 17960 272024 18012
rect 284760 18003 284812 18012
rect 284760 17969 284769 18003
rect 284769 17969 284803 18003
rect 284803 17969 284812 18003
rect 284760 17960 284812 17969
rect 285956 18003 286008 18012
rect 285956 17969 285965 18003
rect 285965 17969 285999 18003
rect 285999 17969 286008 18003
rect 285956 17960 286008 17969
rect 337108 18003 337160 18012
rect 337108 17969 337117 18003
rect 337117 17969 337151 18003
rect 337151 17969 337160 18003
rect 337108 17960 337160 17969
rect 357716 17960 357768 18012
rect 236460 17892 236512 17944
rect 244556 17892 244608 17944
rect 270500 17935 270552 17944
rect 270500 17901 270509 17935
rect 270509 17901 270543 17935
rect 270543 17901 270552 17935
rect 270500 17892 270552 17901
rect 273444 17935 273496 17944
rect 273444 17901 273453 17935
rect 273453 17901 273487 17935
rect 273487 17901 273496 17935
rect 273444 17892 273496 17901
rect 270592 17824 270644 17876
rect 271972 17824 272024 17876
rect 347780 16872 347832 16924
rect 352656 16872 352708 16924
rect 456524 16872 456576 16924
rect 457444 16872 457496 16924
rect 369676 16804 369728 16856
rect 376668 16804 376720 16856
rect 475568 16804 475620 16856
rect 482928 16804 482980 16856
rect 437204 16736 437256 16788
rect 437480 16736 437532 16788
rect 320824 16668 320876 16720
rect 325608 16668 325660 16720
rect 386236 16643 386288 16652
rect 386236 16609 386245 16643
rect 386245 16609 386279 16643
rect 386279 16609 386288 16643
rect 386236 16600 386288 16609
rect 278780 16532 278832 16584
rect 290556 16532 290608 16584
rect 310888 15215 310940 15224
rect 310888 15181 310897 15215
rect 310897 15181 310931 15215
rect 310931 15181 310940 15215
rect 310888 15172 310940 15181
rect 110328 15104 110380 15156
rect 274732 15104 274784 15156
rect 107476 15036 107528 15088
rect 273352 15036 273404 15088
rect 103428 14968 103480 15020
rect 271972 14968 272024 15020
rect 99288 14900 99340 14952
rect 270592 14900 270644 14952
rect 96528 14832 96580 14884
rect 269212 14832 269264 14884
rect 92388 14764 92440 14816
rect 266452 14764 266504 14816
rect 89628 14696 89680 14748
rect 265072 14696 265124 14748
rect 85488 14628 85540 14680
rect 263692 14628 263744 14680
rect 82728 14560 82780 14612
rect 262588 14560 262640 14612
rect 78588 14492 78640 14544
rect 260932 14492 260984 14544
rect 74448 14424 74500 14476
rect 259644 14424 259696 14476
rect 114468 14356 114520 14408
rect 276112 14356 276164 14408
rect 117228 14288 117280 14340
rect 277676 14288 277728 14340
rect 121368 14220 121420 14272
rect 278872 14220 278924 14272
rect 125416 14152 125468 14204
rect 280252 14152 280304 14204
rect 186228 13744 186280 13796
rect 306564 13744 306616 13796
rect 183468 13676 183520 13728
rect 303896 13676 303948 13728
rect 179328 13608 179380 13660
rect 302608 13608 302660 13660
rect 176568 13540 176620 13592
rect 301136 13540 301188 13592
rect 172428 13472 172480 13524
rect 299756 13472 299808 13524
rect 168288 13404 168340 13456
rect 298284 13404 298336 13456
rect 165528 13336 165580 13388
rect 296904 13336 296956 13388
rect 160008 13268 160060 13320
rect 294328 13268 294380 13320
rect 155868 13200 155920 13252
rect 292764 13200 292816 13252
rect 71688 13132 71740 13184
rect 258172 13132 258224 13184
rect 31668 13064 31720 13116
rect 241612 13064 241664 13116
rect 190368 12996 190420 13048
rect 307944 12996 307996 13048
rect 206928 12928 206980 12980
rect 314844 12928 314896 12980
rect 211068 12860 211120 12912
rect 316224 12860 316276 12912
rect 213828 12792 213880 12844
rect 317604 12792 317656 12844
rect 217968 12724 218020 12776
rect 318984 12724 319036 12776
rect 220728 12656 220780 12708
rect 320272 12656 320324 12708
rect 224868 12588 224920 12640
rect 321744 12588 321796 12640
rect 229008 12520 229060 12572
rect 323124 12520 323176 12572
rect 295616 12495 295668 12504
rect 295616 12461 295625 12495
rect 295625 12461 295659 12495
rect 295659 12461 295668 12495
rect 295616 12452 295668 12461
rect 366916 12452 366968 12504
rect 173808 12384 173860 12436
rect 300952 12384 301004 12436
rect 426440 12384 426492 12436
rect 427544 12384 427596 12436
rect 169668 12316 169720 12368
rect 299572 12316 299624 12368
rect 366916 12316 366968 12368
rect 386236 12316 386288 12368
rect 386604 12316 386656 12368
rect 166908 12248 166960 12300
rect 298192 12248 298244 12300
rect 162768 12180 162820 12232
rect 151728 12112 151780 12164
rect 291568 12112 291620 12164
rect 148968 12044 149020 12096
rect 290004 12044 290056 12096
rect 144828 11976 144880 12028
rect 288808 11976 288860 12028
rect 142068 11908 142120 11960
rect 287336 11908 287388 11960
rect 128268 11840 128320 11892
rect 281540 11840 281592 11892
rect 284576 11840 284628 11892
rect 284760 11840 284812 11892
rect 126888 11772 126940 11824
rect 281632 11772 281684 11824
rect 23388 11704 23440 11756
rect 238944 11704 238996 11756
rect 176476 11636 176528 11688
rect 302332 11636 302384 11688
rect 180708 11568 180760 11620
rect 303712 11568 303764 11620
rect 184848 11500 184900 11552
rect 305092 11500 305144 11552
rect 187608 11432 187660 11484
rect 306472 11432 306524 11484
rect 191748 11364 191800 11416
rect 308036 11364 308088 11416
rect 194508 11296 194560 11348
rect 309416 11296 309468 11348
rect 198648 11228 198700 11280
rect 310888 11228 310940 11280
rect 113088 10956 113140 11008
rect 276020 10956 276072 11008
rect 108948 10888 109000 10940
rect 106188 10820 106240 10872
rect 271880 10820 271932 10872
rect 102048 10752 102100 10804
rect 270500 10752 270552 10804
rect 99196 10684 99248 10736
rect 269304 10684 269356 10736
rect 95148 10616 95200 10668
rect 267740 10616 267792 10668
rect 91008 10548 91060 10600
rect 266544 10548 266596 10600
rect 64788 10480 64840 10532
rect 255596 10480 255648 10532
rect 60648 10412 60700 10464
rect 254032 10412 254084 10464
rect 56508 10344 56560 10396
rect 252652 10344 252704 10396
rect 53748 10276 53800 10328
rect 251272 10276 251324 10328
rect 117136 10208 117188 10260
rect 277584 10208 277636 10260
rect 119988 10140 120040 10192
rect 278964 10140 279016 10192
rect 124128 10072 124180 10124
rect 280344 10072 280396 10124
rect 143448 10004 143500 10056
rect 288532 10004 288584 10056
rect 147588 9936 147640 9988
rect 289820 9936 289872 9988
rect 151636 9868 151688 9920
rect 291292 9868 291344 9920
rect 154488 9800 154540 9852
rect 292856 9800 292908 9852
rect 158628 9732 158680 9784
rect 294052 9732 294104 9784
rect 306748 9732 306800 9784
rect 161388 9664 161440 9716
rect 295432 9664 295484 9716
rect 306656 9664 306708 9716
rect 341248 9707 341300 9716
rect 341248 9673 341257 9707
rect 341257 9673 341291 9707
rect 341291 9673 341300 9707
rect 341248 9664 341300 9673
rect 358544 9707 358596 9716
rect 358544 9673 358553 9707
rect 358553 9673 358587 9707
rect 358587 9673 358596 9707
rect 358544 9664 358596 9673
rect 366824 9707 366876 9716
rect 366824 9673 366833 9707
rect 366833 9673 366867 9707
rect 366867 9673 366876 9707
rect 366824 9664 366876 9673
rect 421380 9664 421432 9716
rect 470600 9707 470652 9716
rect 470600 9673 470609 9707
rect 470609 9673 470643 9707
rect 470643 9673 470652 9707
rect 470600 9664 470652 9673
rect 203892 9596 203944 9648
rect 313372 9596 313424 9648
rect 200396 9528 200448 9580
rect 311992 9528 312044 9580
rect 196808 9460 196860 9512
rect 310612 9460 310664 9512
rect 193220 9392 193272 9444
rect 309232 9392 309284 9444
rect 139676 9324 139728 9376
rect 287152 9324 287204 9376
rect 136088 9256 136140 9308
rect 285864 9256 285916 9308
rect 49332 9188 49384 9240
rect 249892 9188 249944 9240
rect 253848 9188 253900 9240
rect 334164 9188 334216 9240
rect 44548 9120 44600 9172
rect 247132 9120 247184 9172
rect 250352 9120 250404 9172
rect 332784 9120 332836 9172
rect 27896 9052 27948 9104
rect 233884 9052 233936 9104
rect 243176 9052 243228 9104
rect 330024 9052 330076 9104
rect 18328 8984 18380 9036
rect 236184 8984 236236 9036
rect 239588 8984 239640 9036
rect 328644 8984 328696 9036
rect 13636 8916 13688 8968
rect 234804 8916 234856 8968
rect 236000 8916 236052 8968
rect 325976 8916 326028 8968
rect 207480 8848 207532 8900
rect 314936 8848 314988 8900
rect 210976 8780 211028 8832
rect 316132 8780 316184 8832
rect 214656 8712 214708 8764
rect 317512 8712 317564 8764
rect 218152 8644 218204 8696
rect 318892 8644 318944 8696
rect 221740 8576 221792 8628
rect 320180 8576 320232 8628
rect 225328 8508 225380 8560
rect 321652 8508 321704 8560
rect 228916 8440 228968 8492
rect 323308 8440 323360 8492
rect 232504 8372 232556 8424
rect 324596 8372 324648 8424
rect 236276 8347 236328 8356
rect 236276 8313 236285 8347
rect 236285 8313 236319 8347
rect 236319 8313 236328 8347
rect 236276 8304 236328 8313
rect 238944 8304 238996 8356
rect 239036 8304 239088 8356
rect 244372 8347 244424 8356
rect 244372 8313 244381 8347
rect 244381 8313 244415 8347
rect 244415 8313 244424 8347
rect 244372 8304 244424 8313
rect 246764 8304 246816 8356
rect 331404 8304 331456 8356
rect 468760 8304 468812 8356
rect 469036 8304 469088 8356
rect 87328 8236 87380 8288
rect 265164 8236 265216 8288
rect 270500 8236 270552 8288
rect 340972 8236 341024 8288
rect 445484 8236 445536 8288
rect 523868 8236 523920 8288
rect 83832 8168 83884 8220
rect 263876 8168 263928 8220
rect 267004 8168 267056 8220
rect 339592 8168 339644 8220
rect 446956 8168 447008 8220
rect 527456 8168 527508 8220
rect 80244 8100 80296 8152
rect 262404 8100 262456 8152
rect 263416 8100 263468 8152
rect 338304 8100 338356 8152
rect 448244 8100 448296 8152
rect 531044 8100 531096 8152
rect 40960 8032 41012 8084
rect 245844 8032 245896 8084
rect 259828 8032 259880 8084
rect 336924 8032 336976 8084
rect 451004 8032 451056 8084
rect 534540 8032 534592 8084
rect 37372 7964 37424 8016
rect 244372 7964 244424 8016
rect 256240 7964 256292 8016
rect 334072 7964 334124 8016
rect 452476 7964 452528 8016
rect 538128 7964 538180 8016
rect 33876 7896 33928 7948
rect 242992 7896 243044 7948
rect 252652 7896 252704 7948
rect 332692 7896 332744 7948
rect 453764 7896 453816 7948
rect 541716 7896 541768 7948
rect 30288 7828 30340 7880
rect 241796 7828 241848 7880
rect 249156 7828 249208 7880
rect 331312 7828 331364 7880
rect 455236 7828 455288 7880
rect 545304 7828 545356 7880
rect 26700 7760 26752 7812
rect 240416 7760 240468 7812
rect 245568 7760 245620 7812
rect 330208 7760 330260 7812
rect 456616 7760 456668 7812
rect 548892 7760 548944 7812
rect 21916 7692 21968 7744
rect 238852 7692 238904 7744
rect 241980 7692 242032 7744
rect 328552 7692 328604 7744
rect 457996 7692 458048 7744
rect 552388 7692 552440 7744
rect 8852 7624 8904 7676
rect 4068 7556 4120 7608
rect 230664 7624 230716 7676
rect 234804 7624 234856 7676
rect 325792 7624 325844 7676
rect 459376 7624 459428 7676
rect 555976 7624 556028 7676
rect 227720 7556 227772 7608
rect 229008 7556 229060 7608
rect 231308 7556 231360 7608
rect 324412 7556 324464 7608
rect 460756 7556 460808 7608
rect 559564 7556 559616 7608
rect 134892 7488 134944 7540
rect 284576 7488 284628 7540
rect 444196 7488 444248 7540
rect 520280 7488 520332 7540
rect 138480 7420 138532 7472
rect 285956 7420 286008 7472
rect 442816 7420 442868 7472
rect 516784 7420 516836 7472
rect 141976 7352 142028 7404
rect 287060 7352 287112 7404
rect 441436 7352 441488 7404
rect 513196 7352 513248 7404
rect 145656 7284 145708 7336
rect 288440 7284 288492 7336
rect 440056 7284 440108 7336
rect 509608 7284 509660 7336
rect 149244 7216 149296 7268
rect 291200 7216 291252 7268
rect 152740 7148 152792 7200
rect 292580 7148 292632 7200
rect 156328 7080 156380 7132
rect 293960 7080 294012 7132
rect 159916 7012 159968 7064
rect 295340 7012 295392 7064
rect 233424 6944 233476 6996
rect 238392 6944 238444 6996
rect 327264 6944 327316 6996
rect 516692 6876 516744 6928
rect 516876 6876 516928 6928
rect 170588 6808 170640 6860
rect 299480 6808 299532 6860
rect 431776 6808 431828 6860
rect 490564 6808 490616 6860
rect 167092 6740 167144 6792
rect 298376 6740 298428 6792
rect 433156 6740 433208 6792
rect 491760 6740 491812 6792
rect 163504 6672 163556 6724
rect 296720 6672 296772 6724
rect 298100 6672 298152 6724
rect 338396 6672 338448 6724
rect 434628 6672 434680 6724
rect 495348 6672 495400 6724
rect 131396 6604 131448 6656
rect 283012 6604 283064 6656
rect 297364 6604 297416 6656
rect 336832 6604 336884 6656
rect 436008 6604 436060 6656
rect 497740 6604 497792 6656
rect 76656 6536 76708 6588
rect 261024 6536 261076 6588
rect 295892 6536 295944 6588
rect 335452 6536 335504 6588
rect 433248 6536 433300 6588
rect 494152 6536 494204 6588
rect 73068 6468 73120 6520
rect 259460 6468 259512 6520
rect 289820 6468 289872 6520
rect 339684 6468 339736 6520
rect 433524 6468 433576 6520
rect 434628 6468 434680 6520
rect 435916 6468 435968 6520
rect 498936 6468 498988 6520
rect 69480 6400 69532 6452
rect 258264 6400 258316 6452
rect 288440 6400 288492 6452
rect 341248 6400 341300 6452
rect 437296 6400 437348 6452
rect 501236 6400 501288 6452
rect 65984 6332 66036 6384
rect 256792 6332 256844 6384
rect 288532 6332 288584 6384
rect 343640 6332 343692 6384
rect 437388 6332 437440 6384
rect 502432 6332 502484 6384
rect 62396 6264 62448 6316
rect 255504 6264 255556 6316
rect 294328 6264 294380 6316
rect 350632 6264 350684 6316
rect 438676 6264 438728 6316
rect 504824 6264 504876 6316
rect 58808 6196 58860 6248
rect 253940 6196 253992 6248
rect 280068 6196 280120 6248
rect 345204 6196 345256 6248
rect 438768 6196 438820 6248
rect 506020 6196 506072 6248
rect 55220 6128 55272 6180
rect 251364 6128 251416 6180
rect 274088 6128 274140 6180
rect 342352 6128 342404 6180
rect 440148 6128 440200 6180
rect 508412 6128 508464 6180
rect 174176 6060 174228 6112
rect 300860 6060 300912 6112
rect 337108 6103 337160 6112
rect 337108 6069 337117 6103
rect 337117 6069 337151 6103
rect 337151 6069 337160 6103
rect 337108 6060 337160 6069
rect 430396 6060 430448 6112
rect 486976 6060 487028 6112
rect 177764 5992 177816 6044
rect 302240 5992 302292 6044
rect 431868 5992 431920 6044
rect 488172 5992 488224 6044
rect 181352 5924 181404 5976
rect 303620 5924 303672 5976
rect 429108 5924 429160 5976
rect 483480 5924 483532 5976
rect 184848 5856 184900 5908
rect 305000 5856 305052 5908
rect 430488 5856 430540 5908
rect 484584 5856 484636 5908
rect 188436 5788 188488 5840
rect 306656 5788 306708 5840
rect 427728 5788 427780 5840
rect 479892 5788 479944 5840
rect 192024 5720 192076 5772
rect 307760 5720 307812 5772
rect 426348 5720 426400 5772
rect 476304 5720 476356 5772
rect 195612 5652 195664 5704
rect 309140 5652 309192 5704
rect 199200 5584 199252 5636
rect 310520 5584 310572 5636
rect 470600 5584 470652 5636
rect 202696 5516 202748 5568
rect 313280 5516 313332 5568
rect 468944 5516 468996 5568
rect 137284 5448 137336 5500
rect 285680 5448 285732 5500
rect 297824 5448 297876 5500
rect 352104 5448 352156 5500
rect 452568 5448 452620 5500
rect 540520 5448 540572 5500
rect 133788 5380 133840 5432
rect 284300 5380 284352 5432
rect 290740 5380 290792 5432
rect 349344 5380 349396 5432
rect 408408 5380 408460 5432
rect 433524 5380 433576 5432
rect 453856 5380 453908 5432
rect 544108 5380 544160 5432
rect 130200 5312 130252 5364
rect 283196 5312 283248 5364
rect 287152 5312 287204 5364
rect 347964 5312 348016 5364
rect 412364 5312 412416 5364
rect 440608 5312 440660 5364
rect 455328 5312 455380 5364
rect 547696 5312 547748 5364
rect 67180 5244 67232 5296
rect 256976 5244 257028 5296
rect 283656 5244 283708 5296
rect 346584 5244 346636 5296
rect 413836 5244 413888 5296
rect 444196 5244 444248 5296
rect 459468 5244 459520 5296
rect 48136 5176 48188 5228
rect 248512 5176 248564 5228
rect 251456 5176 251508 5228
rect 332600 5176 332652 5228
rect 415308 5176 415360 5228
rect 447784 5176 447836 5228
rect 460848 5176 460900 5228
rect 551192 5244 551244 5296
rect 17224 5108 17276 5160
rect 236092 5108 236144 5160
rect 247960 5108 248012 5160
rect 331220 5108 331272 5160
rect 416504 5108 416556 5160
rect 451280 5108 451332 5160
rect 12440 5040 12492 5092
rect 234712 5040 234764 5092
rect 244372 5040 244424 5092
rect 327080 5040 327132 5092
rect 329840 5040 329892 5092
rect 337108 5040 337160 5092
rect 368572 5040 368624 5092
rect 417976 5040 418028 5092
rect 454868 5040 454920 5092
rect 458088 5040 458140 5092
rect 7656 4972 7708 5024
rect 232136 4972 232188 5024
rect 240784 4972 240836 5024
rect 315948 4972 316000 5024
rect 325608 4972 325660 5024
rect 338120 4972 338172 5024
rect 419448 4972 419500 5024
rect 458456 4972 458508 5024
rect 2872 4904 2924 4956
rect 572 4836 624 4888
rect 229100 4904 229152 4956
rect 237196 4904 237248 4956
rect 230112 4836 230164 4888
rect 318708 4904 318760 4956
rect 1676 4768 1728 4820
rect 230756 4768 230808 4820
rect 233700 4768 233752 4820
rect 325700 4836 325752 4888
rect 212264 4700 212316 4752
rect 316040 4700 316092 4752
rect 324320 4768 324372 4820
rect 328736 4904 328788 4956
rect 333612 4904 333664 4956
rect 367192 4904 367244 4956
rect 420736 4904 420788 4956
rect 462044 4972 462096 5024
rect 463516 5108 463568 5160
rect 554780 5176 554832 5228
rect 464988 5040 465040 5092
rect 558368 5108 558420 5160
rect 465632 4972 465684 5024
rect 561956 5040 562008 5092
rect 466184 4904 466236 4956
rect 565544 4972 565596 5024
rect 327080 4836 327132 4888
rect 361672 4836 361724 4888
rect 422208 4836 422260 4888
rect 328460 4768 328512 4820
rect 363052 4768 363104 4820
rect 381544 4768 381596 4820
rect 423588 4768 423640 4820
rect 469128 4836 469180 4888
rect 569040 4904 569092 4956
rect 572628 4836 572680 4888
rect 462136 4768 462188 4820
rect 579804 4768 579856 4820
rect 324228 4700 324280 4752
rect 359188 4700 359240 4752
rect 451096 4700 451148 4752
rect 536932 4700 536984 4752
rect 215852 4632 215904 4684
rect 317420 4632 317472 4684
rect 322940 4632 322992 4684
rect 219348 4564 219400 4616
rect 318800 4564 318852 4616
rect 222936 4496 222988 4548
rect 321560 4564 321612 4616
rect 326528 4632 326580 4684
rect 360292 4632 360344 4684
rect 449808 4632 449860 4684
rect 533436 4632 533488 4684
rect 333980 4564 334032 4616
rect 448336 4564 448388 4616
rect 529848 4564 529900 4616
rect 320364 4496 320416 4548
rect 335360 4496 335412 4548
rect 447048 4496 447100 4548
rect 526260 4496 526312 4548
rect 226524 4428 226576 4480
rect 322572 4428 322624 4480
rect 445576 4428 445628 4480
rect 522672 4428 522724 4480
rect 201500 4360 201552 4412
rect 271144 4360 271196 4412
rect 301412 4360 301464 4412
rect 353484 4360 353536 4412
rect 380164 4360 380216 4412
rect 444288 4360 444340 4412
rect 519084 4360 519136 4412
rect 205088 4292 205140 4344
rect 272524 4292 272576 4344
rect 305000 4292 305052 4344
rect 354956 4292 355008 4344
rect 442908 4292 442960 4344
rect 515588 4292 515640 4344
rect 230572 4224 230624 4276
rect 308588 4224 308640 4276
rect 356152 4224 356204 4276
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 140872 4156 140924 4208
rect 142068 4156 142120 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 160008 4156 160060 4208
rect 175372 4156 175424 4208
rect 176568 4156 176620 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 312084 4156 312136 4208
rect 312176 4156 312228 4208
rect 357716 4156 357768 4208
rect 34980 4088 35032 4140
rect 50344 4088 50396 4140
rect 57612 4088 57664 4140
rect 250444 4088 250496 4140
rect 268108 4088 268160 4140
rect 269028 4088 269080 4140
rect 295892 4088 295944 4140
rect 296720 4088 296772 4140
rect 297916 4088 297968 4140
rect 300308 4088 300360 4140
rect 332416 4088 332468 4140
rect 333244 4088 333296 4140
rect 334716 4088 334768 4140
rect 335268 4088 335320 4140
rect 338764 4088 338816 4140
rect 339500 4088 339552 4140
rect 340788 4088 340840 4140
rect 345664 4088 345716 4140
rect 347872 4088 347924 4140
rect 349068 4088 349120 4140
rect 351184 4088 351236 4140
rect 351368 4088 351420 4140
rect 351828 4088 351880 4140
rect 351920 4088 351972 4140
rect 352564 4088 352616 4140
rect 20720 4020 20772 4072
rect 28264 4020 28316 4072
rect 50528 4020 50580 4072
rect 249064 4020 249116 4072
rect 261024 4020 261076 4072
rect 297364 4020 297416 4072
rect 302608 4020 302660 4072
rect 309784 4020 309836 4072
rect 314568 4020 314620 4072
rect 358912 4020 358964 4072
rect 365720 4020 365772 4072
rect 366916 4020 366968 4072
rect 369216 4020 369268 4072
rect 369768 4020 369820 4072
rect 370412 4088 370464 4140
rect 371148 4088 371200 4140
rect 377588 4088 377640 4140
rect 378048 4088 378100 4140
rect 378784 4088 378836 4140
rect 372620 4020 372672 4072
rect 376760 4020 376812 4072
rect 46940 3952 46992 4004
rect 248696 3952 248748 4004
rect 257436 3952 257488 4004
rect 298100 3952 298152 4004
rect 313372 3952 313424 4004
rect 358820 3952 358872 4004
rect 359740 3952 359792 4004
rect 45744 3884 45796 3936
rect 247684 3884 247736 3936
rect 264612 3884 264664 3936
rect 275284 3884 275336 3936
rect 275928 3884 275980 3936
rect 282460 3884 282512 3936
rect 325608 3884 325660 3936
rect 39764 3816 39816 3868
rect 245936 3816 245988 3868
rect 289544 3816 289596 3868
rect 365812 3884 365864 3936
rect 371608 3884 371660 3936
rect 379980 4088 380032 4140
rect 380808 4088 380860 4140
rect 381176 4088 381228 4140
rect 382188 4088 382240 4140
rect 383568 4088 383620 4140
rect 384304 4088 384356 4140
rect 388260 4088 388312 4140
rect 389088 4088 389140 4140
rect 385868 4020 385920 4072
rect 387064 4020 387116 4072
rect 411168 4020 411220 4072
rect 424968 4156 425020 4208
rect 437480 4088 437532 4140
rect 441528 4224 441580 4276
rect 512000 4224 512052 4276
rect 472716 4156 472768 4208
rect 521476 4088 521528 4140
rect 529204 4088 529256 4140
rect 575020 4088 575072 4140
rect 382372 3952 382424 4004
rect 386604 3952 386656 4004
rect 398104 3952 398156 4004
rect 404912 3952 404964 4004
rect 411076 3952 411128 4004
rect 439412 4020 439464 4072
rect 439596 4020 439648 4072
rect 448428 4020 448480 4072
rect 528652 4020 528704 4072
rect 530584 4020 530636 4072
rect 582196 4020 582248 4072
rect 420184 3952 420236 4004
rect 423956 3952 424008 4004
rect 424324 3952 424376 4004
rect 425152 3952 425204 4004
rect 427084 3952 427136 4004
rect 431132 3952 431184 4004
rect 433984 3952 434036 4004
rect 435824 3952 435876 4004
rect 535736 3952 535788 4004
rect 385316 3884 385368 3936
rect 404268 3884 404320 3936
rect 412548 3884 412600 3936
rect 441804 3884 441856 3936
rect 19524 3748 19576 3800
rect 32404 3748 32456 3800
rect 38568 3748 38620 3800
rect 245752 3748 245804 3800
rect 278872 3748 278924 3800
rect 285956 3748 286008 3800
rect 335544 3748 335596 3800
rect 342904 3816 342956 3868
rect 343088 3816 343140 3868
rect 369124 3816 369176 3868
rect 372804 3816 372856 3868
rect 373908 3816 373960 3868
rect 407028 3816 407080 3868
rect 341524 3748 341576 3800
rect 341892 3748 341944 3800
rect 370136 3748 370188 3800
rect 374000 3748 374052 3800
rect 375288 3748 375340 3800
rect 399484 3748 399536 3800
rect 408500 3748 408552 3800
rect 32680 3680 32732 3732
rect 243084 3680 243136 3732
rect 326436 3680 326488 3732
rect 328460 3680 328512 3732
rect 331220 3680 331272 3732
rect 338304 3680 338356 3732
rect 370504 3680 370556 3732
rect 375196 3680 375248 3732
rect 383844 3680 383896 3732
rect 393136 3680 393188 3732
rect 396632 3680 396684 3732
rect 400036 3680 400088 3732
rect 412088 3680 412140 3732
rect 413928 3816 413980 3868
rect 445392 3816 445444 3868
rect 412456 3748 412508 3800
rect 443000 3748 443052 3800
rect 25504 3612 25556 3664
rect 240324 3612 240376 3664
rect 262220 3612 262272 3664
rect 322572 3612 322624 3664
rect 325240 3612 325292 3664
rect 355324 3612 355376 3664
rect 358084 3612 358136 3664
rect 360936 3612 360988 3664
rect 377404 3612 377456 3664
rect 400128 3612 400180 3664
rect 413192 3612 413244 3664
rect 416688 3612 416740 3664
rect 418068 3612 418120 3664
rect 420736 3612 420788 3664
rect 420828 3612 420880 3664
rect 428464 3680 428516 3732
rect 453672 3884 453724 3936
rect 453948 3884 454000 3936
rect 542912 3884 542964 3936
rect 445668 3816 445720 3868
rect 456708 3816 456760 3868
rect 550088 3816 550140 3868
rect 459652 3748 459704 3800
rect 460020 3748 460072 3800
rect 463240 3748 463292 3800
rect 451188 3680 451240 3732
rect 442264 3612 442316 3664
rect 11244 3544 11296 3596
rect 19984 3544 20036 3596
rect 24308 3544 24360 3596
rect 239036 3544 239088 3596
rect 265808 3544 265860 3596
rect 322848 3544 322900 3596
rect 327080 3544 327132 3596
rect 363604 3544 363656 3596
rect 402244 3544 402296 3596
rect 415676 3544 415728 3596
rect 417424 3544 417476 3596
rect 434536 3587 434588 3596
rect 434536 3553 434545 3587
rect 434545 3553 434579 3587
rect 434579 3553 434588 3587
rect 434536 3544 434588 3553
rect 557172 3748 557224 3800
rect 16028 3476 16080 3528
rect 236276 3476 236328 3528
rect 258632 3476 258684 3528
rect 320364 3476 320416 3528
rect 320456 3476 320508 3528
rect 321468 3476 321520 3528
rect 324044 3476 324096 3528
rect 363144 3476 363196 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 14832 3408 14884 3460
rect 234896 3408 234948 3460
rect 255044 3408 255096 3460
rect 318708 3408 318760 3460
rect 321652 3408 321704 3460
rect 361856 3408 361908 3460
rect 368664 3476 368716 3528
rect 368020 3408 368072 3460
rect 390836 3476 390888 3528
rect 391848 3476 391900 3528
rect 394516 3476 394568 3528
rect 400220 3476 400272 3528
rect 402888 3476 402940 3528
rect 413284 3476 413336 3528
rect 414480 3476 414532 3528
rect 418068 3476 418120 3528
rect 29092 3340 29144 3392
rect 35164 3340 35216 3392
rect 36176 3340 36228 3392
rect 39304 3340 39356 3392
rect 10048 3272 10100 3324
rect 13084 3272 13136 3324
rect 42156 3272 42208 3324
rect 57244 3272 57296 3324
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 61384 3272 61436 3324
rect 52828 3204 52880 3256
rect 53748 3204 53800 3256
rect 54024 3204 54076 3256
rect 43352 3136 43404 3188
rect 64788 3204 64840 3256
rect 251824 3340 251876 3392
rect 289820 3340 289872 3392
rect 299112 3340 299164 3392
rect 302884 3340 302936 3392
rect 310980 3340 311032 3392
rect 353760 3340 353812 3392
rect 375472 3340 375524 3392
rect 71872 3272 71924 3324
rect 253204 3272 253256 3324
rect 61200 3136 61252 3188
rect 66904 3068 66956 3120
rect 68284 3136 68336 3188
rect 71044 3068 71096 3120
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 75460 3136 75512 3188
rect 79324 3136 79376 3188
rect 82636 3136 82688 3188
rect 84844 3204 84896 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 88524 3204 88576 3256
rect 89628 3204 89680 3256
rect 254584 3204 254636 3256
rect 269304 3204 269356 3256
rect 89720 3068 89772 3120
rect 255964 3136 256016 3188
rect 272892 3136 272944 3188
rect 276480 3204 276532 3256
rect 284760 3272 284812 3324
rect 285588 3272 285640 3324
rect 303804 3272 303856 3324
rect 344284 3272 344336 3324
rect 350264 3272 350316 3324
rect 374276 3272 374328 3324
rect 277676 3136 277728 3188
rect 288440 3204 288492 3256
rect 291936 3204 291988 3256
rect 316684 3204 316736 3256
rect 318064 3204 318116 3256
rect 348424 3204 348476 3256
rect 349068 3204 349120 3256
rect 356704 3204 356756 3256
rect 357348 3204 357400 3256
rect 376024 3204 376076 3256
rect 94504 3068 94556 3120
rect 95148 3068 95200 3120
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 98092 3068 98144 3120
rect 99196 3068 99248 3120
rect 101588 3068 101640 3120
rect 102048 3068 102100 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 105176 3068 105228 3120
rect 106188 3068 106240 3120
rect 106372 3068 106424 3120
rect 107476 3068 107528 3120
rect 77944 3000 77996 3052
rect 93308 3000 93360 3052
rect 102600 3000 102652 3052
rect 79048 2932 79100 2984
rect 86132 2932 86184 2984
rect 96896 2932 96948 2984
rect 257344 3068 257396 3120
rect 288532 3136 288584 3188
rect 309784 3136 309836 3188
rect 335912 3136 335964 3188
rect 340696 3136 340748 3188
rect 346676 3136 346728 3188
rect 362132 3136 362184 3188
rect 362868 3136 362920 3188
rect 363328 3136 363380 3188
rect 364248 3136 364300 3188
rect 364524 3136 364576 3188
rect 290464 3068 290516 3120
rect 295524 3068 295576 3120
rect 319444 3068 319496 3120
rect 327724 3068 327776 3120
rect 328828 3068 328880 3120
rect 362224 3068 362276 3120
rect 379704 3408 379756 3460
rect 406384 3408 406436 3460
rect 410892 3408 410944 3460
rect 422760 3408 422812 3460
rect 460848 3476 460900 3528
rect 462228 3476 462280 3528
rect 564348 3680 564400 3732
rect 463608 3612 463660 3664
rect 566740 3612 566792 3664
rect 466368 3544 466420 3596
rect 571432 3544 571484 3596
rect 466276 3476 466328 3528
rect 573824 3476 573876 3528
rect 429936 3408 429988 3460
rect 467932 3408 467984 3460
rect 469036 3408 469088 3460
rect 578608 3408 578660 3460
rect 403624 3340 403676 3392
rect 407304 3340 407356 3392
rect 409788 3340 409840 3392
rect 437020 3340 437072 3392
rect 437480 3340 437532 3392
rect 438216 3340 438268 3392
rect 443644 3340 443696 3392
rect 395988 3272 396040 3324
rect 402520 3272 402572 3324
rect 402796 3272 402848 3324
rect 419172 3272 419224 3324
rect 420276 3272 420328 3324
rect 446588 3272 446640 3324
rect 409144 3204 409196 3256
rect 431224 3204 431276 3256
rect 442356 3204 442408 3256
rect 503628 3272 503680 3324
rect 514024 3340 514076 3392
rect 517888 3340 517940 3392
rect 514392 3272 514444 3324
rect 516876 3272 516928 3324
rect 525064 3340 525116 3392
rect 527824 3340 527876 3392
rect 567844 3340 567896 3392
rect 496544 3204 496596 3256
rect 512644 3204 512696 3256
rect 577412 3272 577464 3324
rect 570236 3204 570288 3256
rect 405648 3136 405700 3188
rect 426348 3136 426400 3188
rect 432328 3136 432380 3188
rect 393228 3068 393280 3120
rect 395436 3068 395488 3120
rect 405004 3068 405056 3120
rect 416872 3068 416924 3120
rect 103980 2864 104032 2916
rect 258724 3000 258776 3052
rect 293132 3000 293184 3052
rect 312544 3000 312596 3052
rect 315764 3000 315816 3052
rect 324228 3000 324280 3052
rect 327632 3000 327684 3052
rect 335912 3000 335964 3052
rect 367284 3000 367336 3052
rect 376392 3000 376444 3052
rect 381636 3000 381688 3052
rect 394608 3000 394660 3052
rect 399024 3000 399076 3052
rect 112352 2932 112404 2984
rect 113088 2932 113140 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 115940 2932 115992 2984
rect 116952 2932 117004 2984
rect 119436 2932 119488 2984
rect 119988 2932 120040 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 111156 2864 111208 2916
rect 258816 2932 258868 2984
rect 316960 2932 317012 2984
rect 344192 2932 344244 2984
rect 351920 2932 351972 2984
rect 352564 2932 352616 2984
rect 374092 2932 374144 2984
rect 395896 2932 395948 2984
rect 401324 2932 401376 2984
rect 416596 2932 416648 2984
rect 431316 3068 431368 3120
rect 475108 3068 475160 3120
rect 475384 3068 475436 3120
rect 477500 3068 477552 3120
rect 505744 3136 505796 3188
rect 563152 3136 563204 3188
rect 482284 3068 482336 3120
rect 524972 3068 525024 3120
rect 560760 3068 560812 3120
rect 421564 3000 421616 3052
rect 450176 3000 450228 3052
rect 489368 3000 489420 3052
rect 509884 3000 509936 3052
rect 523684 3000 523736 3052
rect 553584 3000 553636 3052
rect 418068 2932 418120 2984
rect 428740 2932 428792 2984
rect 429844 2932 429896 2984
rect 448980 2932 449032 2984
rect 481088 2932 481140 2984
rect 520924 2932 520976 2984
rect 546500 2932 546552 2984
rect 95884 2796 95936 2848
rect 114744 2796 114796 2848
rect 260104 2864 260156 2916
rect 319260 2864 319312 2916
rect 326528 2864 326580 2916
rect 344284 2864 344336 2916
rect 121828 2796 121880 2848
rect 261484 2796 261536 2848
rect 330024 2796 330076 2848
rect 335544 2796 335596 2848
rect 354956 2864 355008 2916
rect 355968 2864 356020 2916
rect 359464 2864 359516 2916
rect 398196 2864 398248 2916
rect 403716 2864 403768 2916
rect 420368 2864 420420 2916
rect 356152 2796 356204 2848
rect 375564 2796 375616 2848
rect 388444 2796 388496 2848
rect 424416 2864 424468 2916
rect 438124 2864 438176 2916
rect 387064 2728 387116 2780
rect 439504 2796 439556 2848
rect 449164 2864 449216 2916
rect 460296 2864 460348 2916
rect 473912 2864 473964 2916
rect 521016 2864 521068 2916
rect 539324 2864 539376 2916
rect 466828 2796 466880 2848
rect 518164 2796 518216 2848
rect 532240 2796 532292 2848
rect 457260 2116 457312 2168
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 164700 552 164752 604
rect 165528 552 165580 604
rect 165896 552 165948 604
rect 166908 552 166960 604
rect 169392 552 169444 604
rect 169668 552 169720 604
rect 182548 552 182600 604
rect 183468 552 183520 604
rect 183744 552 183796 604
rect 184756 552 184808 604
rect 187240 552 187292 604
rect 187608 552 187660 604
rect 189632 552 189684 604
rect 190368 552 190420 604
rect 281264 552 281316 604
rect 281448 552 281500 604
rect 345480 595 345532 604
rect 345480 561 345489 595
rect 345489 561 345523 595
rect 345523 561 345532 595
rect 345480 552 345532 561
rect 384672 552 384724 604
rect 384948 552 385000 604
rect 392124 552 392176 604
rect 393044 552 393096 604
rect 405924 552 405976 604
rect 406108 552 406160 604
rect 452476 552 452528 604
rect 463700 552 463752 604
rect 464436 552 464488 604
rect 471520 595 471572 604
rect 471520 561 471529 595
rect 471529 561 471563 595
rect 471563 561 471572 595
rect 471520 552 471572 561
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700670 137876 703520
rect 154132 700738 154160 703520
rect 170324 700942 170352 703520
rect 202800 701010 202828 703520
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 170312 700936 170364 700942
rect 170312 700878 170364 700884
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 218992 700262 219020 703520
rect 218980 700256 219032 700262
rect 218980 700198 219032 700204
rect 235184 700058 235212 703520
rect 235172 700052 235224 700058
rect 235172 699994 235224 700000
rect 267660 699990 267688 703520
rect 267648 699984 267700 699990
rect 267648 699926 267700 699932
rect 283852 699922 283880 703520
rect 283840 699916 283892 699922
rect 283840 699858 283892 699864
rect 300136 699718 300164 703520
rect 328368 700868 328420 700874
rect 328368 700810 328420 700816
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 300780 584662 300808 699654
rect 321468 696992 321520 696998
rect 321468 696934 321520 696940
rect 320088 673532 320140 673538
rect 320088 673474 320140 673480
rect 315948 650072 316000 650078
rect 315948 650014 316000 650020
rect 313188 626612 313240 626618
rect 313188 626554 313240 626560
rect 309048 603152 309100 603158
rect 309048 603094 309100 603100
rect 300768 584656 300820 584662
rect 300768 584598 300820 584604
rect 304540 583704 304592 583710
rect 304540 583646 304592 583652
rect 298192 583636 298244 583642
rect 298192 583578 298244 583584
rect 256056 583568 256108 583574
rect 4802 583536 4858 583545
rect 256056 583510 256108 583516
rect 4802 583471 4858 583480
rect 245568 583500 245620 583506
rect 4712 583364 4764 583370
rect 4712 583306 4764 583312
rect 3148 583092 3200 583098
rect 3148 583034 3200 583040
rect 3056 567384 3108 567390
rect 3054 567352 3056 567361
rect 3108 567352 3110 567361
rect 3054 567287 3110 567296
rect 2780 553104 2832 553110
rect 2778 553072 2780 553081
rect 2832 553072 2834 553081
rect 2778 553007 2834 553016
rect 3056 538688 3108 538694
rect 3054 538656 3056 538665
rect 3108 538656 3110 538665
rect 3054 538591 3110 538600
rect 3056 510264 3108 510270
rect 3056 510206 3108 510212
rect 3068 509969 3096 510206
rect 3054 509960 3110 509969
rect 3054 509895 3110 509904
rect 2780 496732 2832 496738
rect 2780 496674 2832 496680
rect 2792 495553 2820 496674
rect 2778 495544 2834 495553
rect 2778 495479 2834 495488
rect 2964 481160 3016 481166
rect 2962 481128 2964 481137
rect 3016 481128 3018 481137
rect 2962 481063 3018 481072
rect 3160 452441 3188 583034
rect 3240 582888 3292 582894
rect 3240 582830 3292 582836
rect 3146 452432 3202 452441
rect 3146 452367 3202 452376
rect 3148 438864 3200 438870
rect 3148 438806 3200 438812
rect 3160 438025 3188 438806
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 3148 424108 3200 424114
rect 3148 424050 3200 424056
rect 3160 423745 3188 424050
rect 3146 423736 3202 423745
rect 3146 423671 3202 423680
rect 3252 395049 3280 582830
rect 4068 582684 4120 582690
rect 4068 582626 4120 582632
rect 3884 582548 3936 582554
rect 3884 582490 3936 582496
rect 3700 582412 3752 582418
rect 3700 582354 3752 582360
rect 3332 578536 3384 578542
rect 3332 578478 3384 578484
rect 3238 395040 3294 395049
rect 3238 394975 3294 394984
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 3344 366217 3372 578478
rect 3608 578400 3660 578406
rect 3608 578342 3660 578348
rect 3424 578332 3476 578338
rect 3424 578274 3476 578280
rect 3330 366208 3386 366217
rect 3330 366143 3386 366152
rect 3332 324284 3384 324290
rect 3332 324226 3384 324232
rect 3344 323105 3372 324226
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 2780 308848 2832 308854
rect 2778 308816 2780 308825
rect 2832 308816 2834 308825
rect 2778 308751 2834 308760
rect 2962 295216 3018 295225
rect 2962 295151 3018 295160
rect 2976 294409 3004 295151
rect 2962 294400 3018 294409
rect 2962 294335 3018 294344
rect 2780 252544 2832 252550
rect 2780 252486 2832 252492
rect 2792 251297 2820 252486
rect 2778 251288 2834 251297
rect 2778 251223 2834 251232
rect 3056 237380 3108 237386
rect 3056 237322 3108 237328
rect 3068 237017 3096 237322
rect 3054 237008 3110 237017
rect 3054 236943 3110 236952
rect 2780 165504 2832 165510
rect 2780 165446 2832 165452
rect 2792 165073 2820 165446
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 3332 151768 3384 151774
rect 3332 151710 3384 151716
rect 3344 150793 3372 151710
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2780 136536 2832 136542
rect 2780 136478 2832 136484
rect 2792 136377 2820 136478
rect 2778 136368 2834 136377
rect 2778 136303 2834 136312
rect 2780 122324 2832 122330
rect 2780 122266 2832 122272
rect 2792 122097 2820 122266
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3436 93265 3464 578274
rect 3516 578264 3568 578270
rect 3516 578206 3568 578212
rect 3528 107681 3556 578206
rect 3620 179489 3648 578342
rect 3712 193905 3740 582354
rect 3792 579896 3844 579902
rect 3792 579838 3844 579844
rect 3804 208185 3832 579838
rect 3896 222601 3924 582490
rect 3976 578468 4028 578474
rect 3976 578410 4028 578416
rect 3988 265713 4016 578410
rect 4080 280129 4108 582626
rect 4724 553110 4752 583306
rect 4712 553104 4764 553110
rect 4712 553046 4764 553052
rect 4066 280120 4122 280129
rect 4066 280055 4122 280064
rect 3974 265704 4030 265713
rect 3974 265639 4030 265648
rect 3882 222592 3938 222601
rect 3882 222527 3938 222536
rect 3790 208176 3846 208185
rect 3790 208111 3846 208120
rect 3698 193896 3754 193905
rect 3698 193831 3754 193840
rect 3606 179480 3662 179489
rect 3606 179415 3662 179424
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 2780 79824 2832 79830
rect 2780 79766 2832 79772
rect 2792 78985 2820 79766
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 4816 50522 4844 583471
rect 245568 583442 245620 583448
rect 243452 583432 243504 583438
rect 243452 583374 243504 583380
rect 5448 583296 5500 583302
rect 5448 583238 5500 583244
rect 5356 582820 5408 582826
rect 5356 582762 5408 582768
rect 5264 582616 5316 582622
rect 5078 582584 5134 582593
rect 5264 582558 5316 582564
rect 5078 582519 5134 582528
rect 4988 579828 5040 579834
rect 4988 579770 5040 579776
rect 4896 579760 4948 579766
rect 4896 579702 4948 579708
rect 4908 79830 4936 579702
rect 5000 122330 5028 579770
rect 5092 136542 5120 582519
rect 5172 582480 5224 582486
rect 5172 582422 5224 582428
rect 5184 165510 5212 582422
rect 5276 252550 5304 582558
rect 5368 308854 5396 582762
rect 5460 496738 5488 583238
rect 10324 583228 10376 583234
rect 10324 583170 10376 583176
rect 6276 583160 6328 583166
rect 6276 583102 6328 583108
rect 6184 579692 6236 579698
rect 6184 579634 6236 579640
rect 5448 496732 5500 496738
rect 5448 496674 5500 496680
rect 5356 308848 5408 308854
rect 5356 308790 5408 308796
rect 5264 252544 5316 252550
rect 5264 252486 5316 252492
rect 5172 165504 5224 165510
rect 5172 165446 5224 165452
rect 5080 136536 5132 136542
rect 5080 136478 5132 136484
rect 4988 122324 5040 122330
rect 4988 122266 5040 122272
rect 4896 79824 4948 79830
rect 4896 79766 4948 79772
rect 2780 50516 2832 50522
rect 2780 50458 2832 50464
rect 4804 50516 4856 50522
rect 4804 50458 4856 50464
rect 2792 50153 2820 50458
rect 2778 50144 2834 50153
rect 2778 50079 2834 50088
rect 6196 35902 6224 579634
rect 6288 424114 6316 583102
rect 6644 580168 6696 580174
rect 6644 580110 6696 580116
rect 6552 580100 6604 580106
rect 6552 580042 6604 580048
rect 6460 580032 6512 580038
rect 6460 579974 6512 579980
rect 6368 579964 6420 579970
rect 6368 579906 6420 579912
rect 6380 481166 6408 579906
rect 6472 510270 6500 579974
rect 6564 538694 6592 580042
rect 6656 567390 6684 580110
rect 6644 567384 6696 567390
rect 6644 567326 6696 567332
rect 6552 538688 6604 538694
rect 6552 538630 6604 538636
rect 6460 510264 6512 510270
rect 6460 510206 6512 510212
rect 6368 481160 6420 481166
rect 6368 481102 6420 481108
rect 10336 438870 10364 583170
rect 13084 583024 13136 583030
rect 13084 582966 13136 582972
rect 10324 438864 10376 438870
rect 10324 438806 10376 438812
rect 6276 424108 6328 424114
rect 6276 424050 6328 424056
rect 13096 380866 13124 582966
rect 14464 582956 14516 582962
rect 14464 582898 14516 582904
rect 13084 380860 13136 380866
rect 13084 380802 13136 380808
rect 13084 337408 13136 337414
rect 10322 337376 10378 337385
rect 13084 337350 13136 337356
rect 10322 337311 10378 337320
rect 3148 35896 3200 35902
rect 3146 35864 3148 35873
rect 6184 35896 6236 35902
rect 3200 35864 3202 35873
rect 6184 35838 6236 35844
rect 3146 35799 3202 35808
rect 3146 11656 3202 11665
rect 3146 11591 3202 11600
rect 3160 7177 3188 11591
rect 8852 7676 8904 7682
rect 8852 7618 8904 7624
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 3146 7168 3202 7177
rect 3146 7103 3202 7112
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8864 480 8892 7618
rect 10336 3466 10364 337311
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10048 3324 10100 3330
rect 10048 3266 10100 3272
rect 10060 480 10088 3266
rect 11256 480 11284 3538
rect 12452 480 12480 5034
rect 13096 3330 13124 337350
rect 14476 324290 14504 582898
rect 17222 582856 17278 582865
rect 17222 582791 17278 582800
rect 15844 582752 15896 582758
rect 15844 582694 15896 582700
rect 14464 324284 14516 324290
rect 14464 324226 14516 324232
rect 15856 237386 15884 582694
rect 15844 237380 15896 237386
rect 15844 237322 15896 237328
rect 17236 151774 17264 582791
rect 24122 582720 24178 582729
rect 24122 582655 24178 582664
rect 19984 337476 20036 337482
rect 19984 337418 20036 337424
rect 17224 151768 17276 151774
rect 17224 151710 17276 151716
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13084 3324 13136 3330
rect 13084 3266 13136 3272
rect 13648 480 13676 8910
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 480 14872 3402
rect 16040 480 16068 3470
rect 17236 480 17264 5102
rect 18340 480 18368 8978
rect 19524 3800 19576 3806
rect 19524 3742 19576 3748
rect 19536 480 19564 3742
rect 19996 3602 20024 337418
rect 24136 64870 24164 582655
rect 243464 579972 243492 583374
rect 245580 579972 245608 583442
rect 251824 581120 251876 581126
rect 251824 581062 251876 581068
rect 251836 579972 251864 581062
rect 256068 579972 256096 583510
rect 293958 583264 294014 583273
rect 293958 583199 294014 583208
rect 289728 581528 289780 581534
rect 289728 581470 289780 581476
rect 287612 581460 287664 581466
rect 287612 581402 287664 581408
rect 283472 581392 283524 581398
rect 283472 581334 283524 581340
rect 281356 581324 281408 581330
rect 281356 581266 281408 581272
rect 275008 581256 275060 581262
rect 275008 581198 275060 581204
rect 268660 581188 268712 581194
rect 268660 581130 268712 581136
rect 264520 581052 264572 581058
rect 264520 580994 264572 581000
rect 262404 580304 262456 580310
rect 262404 580246 262456 580252
rect 262416 579972 262444 580246
rect 264532 579972 264560 580994
rect 268672 579972 268700 581130
rect 275020 579972 275048 581198
rect 281368 579972 281396 581266
rect 283484 579972 283512 581334
rect 287624 579972 287652 581402
rect 289740 579972 289768 581470
rect 293972 579972 294000 583199
rect 296076 581596 296128 581602
rect 296076 581538 296128 581544
rect 296088 579972 296116 581538
rect 298204 579972 298232 583578
rect 300306 583400 300362 583409
rect 300306 583335 300362 583344
rect 300320 579972 300348 583335
rect 302424 581664 302476 581670
rect 302424 581606 302476 581612
rect 302436 579972 302464 581606
rect 304552 579972 304580 583646
rect 306564 580236 306616 580242
rect 306564 580178 306616 580184
rect 306576 579972 306604 580178
rect 309060 579986 309088 603094
rect 311808 592068 311860 592074
rect 311808 592010 311860 592016
rect 311820 580122 311848 592010
rect 308706 579958 309088 579986
rect 311268 580094 311848 580122
rect 311268 579850 311296 580094
rect 313200 579986 313228 626554
rect 312938 579958 313228 579986
rect 315960 579850 315988 650014
rect 317328 638988 317380 638994
rect 317328 638930 317380 638936
rect 317340 579986 317368 638930
rect 320100 580122 320128 673474
rect 317170 579958 317368 579986
rect 319732 580094 320128 580122
rect 319732 579850 319760 580094
rect 321480 579986 321508 696934
rect 324228 685908 324280 685914
rect 324228 685850 324280 685856
rect 321402 579958 321508 579986
rect 324240 579850 324268 685850
rect 325516 584452 325568 584458
rect 325516 584394 325568 584400
rect 325528 579972 325556 584394
rect 328380 579850 328408 700810
rect 329748 700800 329800 700806
rect 329748 700742 329800 700748
rect 329760 579972 329788 700742
rect 332520 699718 332548 703520
rect 336648 700188 336700 700194
rect 336648 700130 336700 700136
rect 335268 700120 335320 700126
rect 335268 700062 335320 700068
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 331864 584520 331916 584526
rect 331864 584462 331916 584468
rect 331876 579972 331904 584462
rect 335280 580122 335308 700062
rect 334452 580094 335308 580122
rect 334452 579850 334480 580094
rect 336660 579850 336688 700130
rect 343548 699848 343600 699854
rect 343548 699790 343600 699796
rect 340788 699780 340840 699786
rect 340788 699722 340840 699728
rect 338212 584588 338264 584594
rect 338212 584530 338264 584536
rect 338224 579972 338252 584530
rect 340800 579986 340828 699722
rect 340354 579958 340828 579986
rect 343560 579850 343588 699790
rect 348804 699718 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365208 703474
rect 358820 701004 358872 701010
rect 358820 700946 358872 700952
rect 356060 700052 356112 700058
rect 356060 699994 356112 700000
rect 351920 699984 351972 699990
rect 351920 699926 351972 699932
rect 346400 699712 346452 699718
rect 346400 699654 346452 699660
rect 347780 699712 347832 699718
rect 347780 699654 347832 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 344468 584724 344520 584730
rect 344468 584666 344520 584672
rect 344480 579972 344508 584666
rect 346412 579986 346440 699654
rect 346412 579958 346610 579986
rect 310822 579822 311296 579850
rect 315054 579822 315988 579850
rect 319286 579822 319760 579850
rect 323426 579822 324268 579850
rect 327658 579822 328408 579850
rect 334006 579822 334480 579850
rect 336122 579822 336688 579850
rect 342378 579822 343588 579850
rect 347792 579850 347820 699654
rect 350816 584656 350868 584662
rect 350816 584598 350868 584604
rect 350828 579972 350856 584598
rect 351932 579850 351960 699926
rect 354680 699916 354732 699922
rect 354680 699858 354732 699864
rect 354692 579986 354720 699858
rect 354692 579958 355074 579986
rect 356072 579850 356100 699994
rect 358832 579850 358860 700946
rect 362960 700936 363012 700942
rect 362960 700878 363012 700884
rect 360200 700256 360252 700262
rect 360200 700198 360252 700204
rect 360212 580122 360240 700198
rect 360212 580094 360884 580122
rect 360856 579850 360884 580094
rect 362972 579986 363000 700878
rect 364340 700664 364392 700670
rect 364340 700606 364392 700612
rect 364352 580122 364380 700606
rect 365180 687818 365208 703446
rect 367100 700732 367152 700738
rect 367100 700674 367152 700680
rect 364616 687812 364668 687818
rect 364616 687754 364668 687760
rect 365168 687812 365220 687818
rect 365168 687754 365220 687760
rect 364628 685846 364656 687754
rect 364616 685840 364668 685846
rect 364616 685782 364668 685788
rect 364524 676252 364576 676258
rect 364524 676194 364576 676200
rect 364536 669338 364564 676194
rect 364536 669310 364748 669338
rect 364720 650026 364748 669310
rect 364536 649998 364748 650026
rect 364536 630714 364564 649998
rect 364536 630686 364656 630714
rect 364628 618254 364656 630686
rect 364616 618248 364668 618254
rect 364616 618190 364668 618196
rect 364524 608660 364576 608666
rect 364524 608602 364576 608608
rect 364536 601746 364564 608602
rect 364536 601718 364656 601746
rect 364628 598942 364656 601718
rect 364616 598936 364668 598942
rect 364616 598878 364668 598884
rect 364708 589348 364760 589354
rect 364708 589290 364760 589296
rect 364720 584730 364748 589290
rect 364708 584724 364760 584730
rect 364708 584666 364760 584672
rect 364352 580094 365208 580122
rect 365180 579986 365208 580094
rect 362972 579958 363446 579986
rect 365180 579958 365562 579986
rect 367112 579850 367140 700674
rect 368480 700596 368532 700602
rect 368480 700538 368532 700544
rect 368492 580122 368520 700538
rect 374000 700528 374052 700534
rect 374000 700470 374052 700476
rect 371240 700460 371292 700466
rect 371240 700402 371292 700408
rect 368492 580094 369348 580122
rect 369320 579850 369348 580094
rect 371252 579850 371280 700402
rect 374012 579972 374040 700470
rect 375380 700392 375432 700398
rect 375380 700334 375432 700340
rect 378138 700360 378194 700369
rect 375392 579850 375420 700334
rect 378138 700295 378194 700304
rect 379520 700324 379572 700330
rect 378152 579986 378180 700295
rect 379520 700266 379572 700272
rect 378152 579958 378258 579986
rect 379532 579850 379560 700266
rect 397472 699786 397500 703520
rect 413664 699854 413692 703520
rect 413652 699848 413704 699854
rect 413652 699790 413704 699796
rect 397460 699780 397512 699786
rect 397460 699722 397512 699728
rect 429856 688634 429884 703520
rect 462332 700126 462360 703520
rect 478524 700194 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 462320 700120 462372 700126
rect 462320 700062 462372 700068
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700874 527220 703520
rect 527180 700868 527232 700874
rect 527180 700810 527232 700816
rect 543476 700806 543504 703520
rect 543464 700800 543516 700806
rect 543464 700742 543516 700748
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 382280 681760 382332 681766
rect 382280 681702 382332 681708
rect 382292 579986 382320 681702
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 386420 667956 386472 667962
rect 386420 667898 386472 667904
rect 383660 652792 383712 652798
rect 383660 652734 383712 652740
rect 382292 579958 382398 579986
rect 383672 579850 383700 652734
rect 386432 579986 386460 667898
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 429672 659682 429700 666538
rect 429488 659654 429700 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 429488 647290 429516 659654
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 494072 644450 494100 654094
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 387800 623824 387852 623830
rect 387800 623766 387852 623772
rect 386432 579958 386630 579986
rect 387812 579850 387840 623766
rect 429396 621058 429424 630550
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 429396 621030 429516 621058
rect 429488 611386 429516 621030
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 391940 610020 391992 610026
rect 391940 609962 391992 609968
rect 390560 594856 390612 594862
rect 390560 594798 390612 594804
rect 390572 579986 390600 594798
rect 390572 579958 390862 579986
rect 391952 579850 391980 609962
rect 429396 608598 429424 611238
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 494256 596222 494284 605798
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 429672 584594 429700 589290
rect 429660 584588 429712 584594
rect 429660 584530 429712 584536
rect 494256 584526 494284 596006
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 494244 584520 494296 584526
rect 494244 584462 494296 584468
rect 559392 584458 559420 589290
rect 559380 584452 559432 584458
rect 559380 584394 559432 584400
rect 471428 583704 471480 583710
rect 471428 583646 471480 583652
rect 471336 583636 471388 583642
rect 471336 583578 471388 583584
rect 460294 583536 460350 583545
rect 460294 583471 460350 583480
rect 399208 583364 399260 583370
rect 399208 583306 399260 583312
rect 395068 580168 395120 580174
rect 395068 580110 395120 580116
rect 395080 579972 395108 580110
rect 397092 580100 397144 580106
rect 397092 580042 397144 580048
rect 397104 579972 397132 580042
rect 399220 579972 399248 583306
rect 405556 583296 405608 583302
rect 405556 583238 405608 583244
rect 400956 580032 401008 580038
rect 401008 579980 401350 579986
rect 400956 579974 401350 579980
rect 400968 579958 401350 579974
rect 403176 579970 403466 579986
rect 405568 579972 405596 583238
rect 411904 583228 411956 583234
rect 411904 583170 411956 583176
rect 409788 583160 409840 583166
rect 409788 583102 409840 583108
rect 407672 583092 407724 583098
rect 407672 583034 407724 583040
rect 407684 579972 407712 583034
rect 409800 579972 409828 583102
rect 411916 579972 411944 583170
rect 420274 583128 420330 583137
rect 420274 583063 420330 583072
rect 418160 583024 418212 583030
rect 418160 582966 418212 582972
rect 414020 582888 414072 582894
rect 414020 582830 414072 582836
rect 414032 579972 414060 582830
rect 418172 579972 418200 582966
rect 420288 579972 420316 583063
rect 426622 582992 426678 583001
rect 424508 582956 424560 582962
rect 426622 582927 426678 582936
rect 424508 582898 424560 582904
rect 422392 582820 422444 582826
rect 422392 582762 422444 582768
rect 422404 579972 422432 582762
rect 424520 579972 424548 582898
rect 426636 579972 426664 582927
rect 449806 582856 449862 582865
rect 449806 582791 449862 582800
rect 437112 582752 437164 582758
rect 437112 582694 437164 582700
rect 430856 582684 430908 582690
rect 430856 582626 430908 582632
rect 430868 579972 430896 582626
rect 432972 582616 433024 582622
rect 432972 582558 433024 582564
rect 432984 579972 433012 582558
rect 434996 582548 435048 582554
rect 434996 582490 435048 582496
rect 435008 579972 435036 582490
rect 437124 579972 437152 582694
rect 447690 582584 447746 582593
rect 447690 582519 447746 582528
rect 445576 582480 445628 582486
rect 445576 582422 445628 582428
rect 443460 582412 443512 582418
rect 443460 582354 443512 582360
rect 443472 579972 443500 582354
rect 445588 579972 445616 582422
rect 447704 579972 447732 582519
rect 449820 579972 449848 582791
rect 460308 579972 460336 583471
rect 462410 582720 462466 582729
rect 462410 582655 462466 582664
rect 462424 579972 462452 582655
rect 469588 581664 469640 581670
rect 469588 581606 469640 581612
rect 403164 579964 403466 579970
rect 403216 579958 403466 579964
rect 403164 579906 403216 579912
rect 438860 579896 438912 579902
rect 347792 579822 348726 579850
rect 351932 579822 352958 579850
rect 356072 579822 357190 579850
rect 358832 579822 359306 579850
rect 360856 579822 361330 579850
rect 367112 579822 367678 579850
rect 369320 579822 369794 579850
rect 371252 579822 371910 579850
rect 375392 579822 376142 579850
rect 379532 579822 380282 579850
rect 383672 579822 384514 579850
rect 387812 579822 388746 579850
rect 391952 579822 392978 579850
rect 438912 579844 439254 579850
rect 438860 579838 439254 579844
rect 438872 579822 439254 579838
rect 451568 579834 451950 579850
rect 451556 579828 451950 579834
rect 451608 579822 451950 579828
rect 451556 579770 451608 579776
rect 458272 579760 458324 579766
rect 458206 579708 458272 579714
rect 468482 579728 468538 579737
rect 458206 579702 458324 579708
rect 458206 579686 458312 579702
rect 464264 579698 464554 579714
rect 464252 579692 464554 579698
rect 464304 579686 464554 579692
rect 468538 579686 468786 579714
rect 468482 579663 468538 579672
rect 464252 579634 464304 579640
rect 270802 579426 271184 579442
rect 270802 579420 271196 579426
rect 270802 579414 271144 579420
rect 271144 579362 271196 579368
rect 247960 579352 248012 579358
rect 231122 579320 231178 579329
rect 230874 579278 231122 579306
rect 232962 579320 233018 579329
rect 232898 579278 232962 579306
rect 231122 579255 231178 579264
rect 235262 579320 235318 579329
rect 235014 579278 235262 579306
rect 232962 579255 233018 579264
rect 237194 579320 237250 579329
rect 237130 579278 237194 579306
rect 235262 579255 235318 579264
rect 239402 579320 239458 579329
rect 239246 579278 239402 579306
rect 237194 579255 237250 579264
rect 241426 579320 241482 579329
rect 241362 579278 241426 579306
rect 239402 579255 239458 579264
rect 247710 579300 247960 579306
rect 254216 579352 254268 579358
rect 247710 579294 248012 579300
rect 249522 579320 249578 579329
rect 247710 579278 248000 579294
rect 241426 579255 241482 579264
rect 249578 579278 249734 579306
rect 253966 579300 254216 579306
rect 258448 579352 258500 579358
rect 253966 579294 254268 579300
rect 258198 579300 258448 579306
rect 260656 579352 260708 579358
rect 258198 579294 258500 579300
rect 260314 579300 260656 579306
rect 266912 579352 266964 579358
rect 260314 579294 260708 579300
rect 266662 579300 266912 579306
rect 273168 579352 273220 579358
rect 266662 579294 266964 579300
rect 272918 579300 273168 579306
rect 277308 579352 277360 579358
rect 272918 579294 273220 579300
rect 277150 579300 277308 579306
rect 279608 579352 279660 579358
rect 277150 579294 277360 579300
rect 279266 579300 279608 579306
rect 285772 579352 285824 579358
rect 279266 579294 279660 579300
rect 285614 579300 285772 579306
rect 292120 579352 292172 579358
rect 285614 579294 285824 579300
rect 291870 579300 292120 579306
rect 291870 579294 292172 579300
rect 415676 579352 415728 579358
rect 428372 579352 428424 579358
rect 415728 579300 416070 579306
rect 415676 579294 416070 579300
rect 441068 579352 441120 579358
rect 428424 579300 428766 579306
rect 428372 579294 428766 579300
rect 453580 579352 453632 579358
rect 441120 579300 441370 579306
rect 441068 579294 441370 579300
rect 455788 579352 455840 579358
rect 453632 579300 453974 579306
rect 453580 579294 453974 579300
rect 466458 579320 466514 579329
rect 455840 579300 456090 579306
rect 455788 579294 456090 579300
rect 253966 579278 254256 579294
rect 258198 579278 258488 579294
rect 260314 579278 260696 579294
rect 266662 579278 266952 579294
rect 272918 579278 273208 579294
rect 277150 579278 277348 579294
rect 279266 579278 279648 579294
rect 285614 579278 285812 579294
rect 291870 579278 292160 579294
rect 415688 579278 416070 579294
rect 428384 579278 428766 579294
rect 441080 579278 441370 579294
rect 453592 579278 453974 579294
rect 455800 579278 456090 579294
rect 249522 579255 249578 579264
rect 466514 579278 466670 579306
rect 466458 579255 466514 579264
rect 469600 557530 469628 581606
rect 469680 581596 469732 581602
rect 469680 581538 469732 581544
rect 469588 557524 469640 557530
rect 469588 557466 469640 557472
rect 469692 510610 469720 581538
rect 469772 581528 469824 581534
rect 469772 581470 469824 581476
rect 469680 510604 469732 510610
rect 469680 510546 469732 510552
rect 469784 463690 469812 581470
rect 470508 581460 470560 581466
rect 470508 581402 470560 581408
rect 470416 581392 470468 581398
rect 470416 581334 470468 581340
rect 470324 581324 470376 581330
rect 470324 581266 470376 581272
rect 470232 581256 470284 581262
rect 470232 581198 470284 581204
rect 470048 581188 470100 581194
rect 470048 581130 470100 581136
rect 469864 581120 469916 581126
rect 469864 581062 469916 581068
rect 469772 463684 469824 463690
rect 469772 463626 469824 463632
rect 232516 340190 232898 340218
rect 244752 340190 245226 340218
rect 290292 340190 290766 340218
rect 291764 340190 292238 340218
rect 294708 340190 295182 340218
rect 326540 340190 327014 340218
rect 386800 340190 387274 340218
rect 399510 340190 399892 340218
rect 422970 340190 423444 340218
rect 424442 340190 424916 340218
rect 460230 340190 460612 340218
rect 229112 340054 230046 340082
rect 230506 340054 230612 340082
rect 71044 338088 71096 338094
rect 71044 338030 71096 338036
rect 66904 338020 66956 338026
rect 66904 337962 66956 337968
rect 61384 337952 61436 337958
rect 61384 337894 61436 337900
rect 57244 337884 57296 337890
rect 57244 337826 57296 337832
rect 50344 337816 50396 337822
rect 50344 337758 50396 337764
rect 39304 337748 39356 337754
rect 39304 337690 39356 337696
rect 32404 337680 32456 337686
rect 32404 337622 32456 337628
rect 28264 337544 28316 337550
rect 28264 337486 28316 337492
rect 24124 64864 24176 64870
rect 24124 64806 24176 64812
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20732 480 20760 4014
rect 21928 480 21956 7686
rect 23400 610 23428 11698
rect 27896 9104 27948 9110
rect 27896 9046 27948 9052
rect 26700 7812 26752 7818
rect 26700 7754 26752 7760
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3538
rect 25516 480 25544 3606
rect 26712 480 26740 7754
rect 27908 480 27936 9046
rect 28276 4078 28304 337486
rect 31668 13116 31720 13122
rect 31668 13058 31720 13064
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 480 29132 3334
rect 30300 480 30328 7822
rect 31680 626 31708 13058
rect 32416 3806 32444 337622
rect 35164 337612 35216 337618
rect 35164 337554 35216 337560
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3674
rect 33888 480 33916 7890
rect 34980 4140 35032 4146
rect 34980 4082 35032 4088
rect 34992 480 35020 4082
rect 35176 3398 35204 337554
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36188 480 36216 3334
rect 37384 480 37412 7958
rect 38568 3800 38620 3806
rect 38568 3742 38620 3748
rect 38580 480 38608 3742
rect 39316 3398 39344 337690
rect 49332 9240 49384 9246
rect 49332 9182 49384 9188
rect 44548 9172 44600 9178
rect 44548 9114 44600 9120
rect 40960 8084 41012 8090
rect 40960 8026 41012 8032
rect 39764 3868 39816 3874
rect 39764 3810 39816 3816
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39776 480 39804 3810
rect 40972 480 41000 8026
rect 42156 3324 42208 3330
rect 42156 3266 42208 3272
rect 42168 480 42196 3266
rect 43352 3188 43404 3194
rect 43352 3130 43404 3136
rect 43364 480 43392 3130
rect 44560 480 44588 9114
rect 48136 5228 48188 5234
rect 48136 5170 48188 5176
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45756 480 45784 3878
rect 46952 480 46980 3946
rect 48148 480 48176 5170
rect 49344 480 49372 9182
rect 50356 4146 50384 337758
rect 56508 10396 56560 10402
rect 56508 10338 56560 10344
rect 53748 10328 53800 10334
rect 53748 10270 53800 10276
rect 51630 6216 51686 6225
rect 51630 6151 51686 6160
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50540 480 50568 4014
rect 51644 480 51672 6151
rect 53760 3262 53788 10270
rect 55220 6180 55272 6186
rect 55220 6122 55272 6128
rect 52828 3256 52880 3262
rect 52828 3198 52880 3204
rect 53748 3256 53800 3262
rect 53748 3198 53800 3204
rect 54024 3256 54076 3262
rect 54024 3198 54076 3204
rect 52840 480 52868 3198
rect 54036 480 54064 3198
rect 55232 480 55260 6122
rect 56520 3482 56548 10338
rect 56428 3454 56548 3482
rect 56428 480 56456 3454
rect 57256 3330 57284 337826
rect 57978 337784 58034 337793
rect 57978 337719 57980 337728
rect 58032 337719 58034 337728
rect 57980 337690 58032 337696
rect 60648 10464 60700 10470
rect 60648 10406 60700 10412
rect 58808 6248 58860 6254
rect 58808 6190 58860 6196
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57624 480 57652 4082
rect 58820 480 58848 6190
rect 60660 3398 60688 10406
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61396 3330 61424 337894
rect 64788 10532 64840 10538
rect 64788 10474 64840 10480
rect 62396 6316 62448 6322
rect 62396 6258 62448 6264
rect 61384 3324 61436 3330
rect 61384 3266 61436 3272
rect 61200 3188 61252 3194
rect 61200 3130 61252 3136
rect 61212 480 61240 3130
rect 62408 480 62436 6258
rect 64800 3398 64828 10474
rect 65984 6384 66036 6390
rect 65984 6326 66036 6332
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 63604 480 63632 3334
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64800 480 64828 3198
rect 65996 480 66024 6326
rect 66916 3126 66944 337962
rect 67546 337784 67602 337793
rect 67546 337719 67548 337728
rect 67600 337719 67602 337728
rect 67548 337690 67600 337696
rect 69480 6452 69532 6458
rect 69480 6394 69532 6400
rect 67180 5296 67232 5302
rect 67180 5238 67232 5244
rect 66904 3120 66956 3126
rect 66904 3062 66956 3068
rect 67192 480 67220 5238
rect 68284 3188 68336 3194
rect 68284 3130 68336 3136
rect 68296 480 68324 3130
rect 69492 480 69520 6394
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 70688 480 70716 3334
rect 71056 3126 71084 338030
rect 79324 337340 79376 337346
rect 79324 337282 79376 337288
rect 77944 337204 77996 337210
rect 77944 337146 77996 337152
rect 74448 14476 74500 14482
rect 74448 14418 74500 14424
rect 71688 13184 71740 13190
rect 71688 13126 71740 13132
rect 71700 3398 71728 13126
rect 73068 6520 73120 6526
rect 73068 6462 73120 6468
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71044 3120 71096 3126
rect 71044 3062 71096 3068
rect 71884 480 71912 3266
rect 73080 480 73108 6462
rect 74460 3380 74488 14418
rect 76656 6588 76708 6594
rect 76656 6530 76708 6536
rect 74276 3352 74488 3380
rect 74276 480 74304 3352
rect 75460 3188 75512 3194
rect 75460 3130 75512 3136
rect 75472 480 75500 3130
rect 76668 480 76696 6530
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 77864 480 77892 3198
rect 77956 3058 77984 337146
rect 78588 14544 78640 14550
rect 78588 14486 78640 14492
rect 78600 3262 78628 14486
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 79336 3194 79364 337282
rect 84844 337272 84896 337278
rect 84844 337214 84896 337220
rect 82728 14612 82780 14618
rect 82728 14554 82780 14560
rect 80244 8152 80296 8158
rect 80244 8094 80296 8100
rect 79324 3188 79376 3194
rect 79324 3130 79376 3136
rect 77944 3052 77996 3058
rect 77944 2994 77996 3000
rect 79048 2984 79100 2990
rect 79048 2926 79100 2932
rect 79060 480 79088 2926
rect 80256 480 80284 8094
rect 82740 3262 82768 14554
rect 83832 8220 83884 8226
rect 83832 8162 83884 8168
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 81452 480 81480 3198
rect 82636 3188 82688 3194
rect 82636 3130 82688 3136
rect 82648 480 82676 3130
rect 83844 480 83872 8162
rect 84856 3262 84884 337214
rect 100668 337136 100720 337142
rect 100668 337078 100720 337084
rect 95884 337068 95936 337074
rect 95884 337010 95936 337016
rect 92388 14816 92440 14822
rect 92388 14758 92440 14764
rect 89628 14748 89680 14754
rect 89628 14690 89680 14696
rect 85488 14680 85540 14686
rect 85488 14622 85540 14628
rect 85500 3262 85528 14622
rect 87328 8288 87380 8294
rect 87328 8230 87380 8236
rect 84844 3256 84896 3262
rect 84844 3198 84896 3204
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84948 480 84976 3198
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 86144 480 86172 2926
rect 87340 480 87368 8230
rect 89640 3262 89668 14690
rect 91008 10600 91060 10606
rect 91008 10542 91060 10548
rect 91020 3482 91048 10542
rect 92400 3482 92428 14758
rect 95148 10668 95200 10674
rect 95148 10610 95200 10616
rect 90928 3454 91048 3482
rect 92124 3454 92428 3482
rect 88524 3256 88576 3262
rect 88524 3198 88576 3204
rect 89628 3256 89680 3262
rect 89628 3198 89680 3204
rect 88536 480 88564 3198
rect 89720 3120 89772 3126
rect 89720 3062 89772 3068
rect 89732 480 89760 3062
rect 90928 480 90956 3454
rect 92124 480 92152 3454
rect 95160 3126 95188 10610
rect 94504 3120 94556 3126
rect 94504 3062 94556 3068
rect 95148 3120 95200 3126
rect 95148 3062 95200 3068
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 93308 3052 93360 3058
rect 93308 2994 93360 3000
rect 93320 480 93348 2994
rect 94516 480 94544 3062
rect 95712 480 95740 3062
rect 95896 2854 95924 337010
rect 99288 14952 99340 14958
rect 99288 14894 99340 14900
rect 96528 14884 96580 14890
rect 96528 14826 96580 14832
rect 96540 3126 96568 14826
rect 99196 10736 99248 10742
rect 99196 10678 99248 10684
rect 99208 3126 99236 10678
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 98092 3120 98144 3126
rect 98092 3062 98144 3068
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 96896 2984 96948 2990
rect 96896 2926 96948 2932
rect 95884 2848 95936 2854
rect 95884 2790 95936 2796
rect 96908 480 96936 2926
rect 98104 480 98132 3062
rect 99300 480 99328 14894
rect 100680 3482 100708 337078
rect 107568 337000 107620 337006
rect 107568 336942 107620 336948
rect 102784 336932 102836 336938
rect 102784 336874 102836 336880
rect 102048 10804 102100 10810
rect 102048 10746 102100 10752
rect 100496 3454 100708 3482
rect 100496 480 100524 3454
rect 102060 3126 102088 10746
rect 102796 3210 102824 336874
rect 107476 15088 107528 15094
rect 107476 15030 107528 15036
rect 103428 15020 103480 15026
rect 103428 14962 103480 14968
rect 102612 3182 102824 3210
rect 101588 3120 101640 3126
rect 101588 3062 101640 3068
rect 102048 3120 102100 3126
rect 102048 3062 102100 3068
rect 101600 480 101628 3062
rect 102612 3058 102640 3182
rect 103440 3126 103468 14962
rect 106188 10872 106240 10878
rect 106188 10814 106240 10820
rect 106200 3126 106228 10814
rect 107488 3126 107516 15030
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 105176 3120 105228 3126
rect 105176 3062 105228 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 102600 3052 102652 3058
rect 102600 2994 102652 3000
rect 102796 480 102824 3062
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 103992 480 104020 2858
rect 105188 480 105216 3062
rect 106384 480 106412 3062
rect 107580 480 107608 336942
rect 118608 336864 118660 336870
rect 118608 336806 118660 336812
rect 110328 15156 110380 15162
rect 110328 15098 110380 15104
rect 108948 10940 109000 10946
rect 108948 10882 109000 10888
rect 108960 3482 108988 10882
rect 110340 3482 110368 15098
rect 114468 14408 114520 14414
rect 114468 14350 114520 14356
rect 113088 11008 113140 11014
rect 113088 10950 113140 10956
rect 108776 3454 108988 3482
rect 109972 3454 110368 3482
rect 108776 480 108804 3454
rect 109972 480 110000 3454
rect 113100 2990 113128 10950
rect 114480 2990 114508 14350
rect 117228 14340 117280 14346
rect 117228 14282 117280 14288
rect 117136 10260 117188 10266
rect 117136 10202 117188 10208
rect 117148 3618 117176 10202
rect 116964 3590 117176 3618
rect 116964 2990 116992 3590
rect 117240 3482 117268 14282
rect 117148 3454 117268 3482
rect 112352 2984 112404 2990
rect 112352 2926 112404 2932
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 115940 2984 115992 2990
rect 115940 2926 115992 2932
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 111168 480 111196 2858
rect 112364 480 112392 2926
rect 113560 480 113588 2926
rect 114744 2848 114796 2854
rect 114744 2790 114796 2796
rect 114756 480 114784 2790
rect 115952 480 115980 2926
rect 117148 480 117176 3454
rect 118620 3346 118648 336806
rect 125508 336796 125560 336802
rect 125508 336738 125560 336744
rect 121368 14272 121420 14278
rect 121368 14214 121420 14220
rect 119988 10192 120040 10198
rect 119988 10134 120040 10140
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 120000 2990 120028 10134
rect 121380 2990 121408 14214
rect 125416 14204 125468 14210
rect 125416 14146 125468 14152
rect 124128 10124 124180 10130
rect 124128 10066 124180 10072
rect 124140 3482 124168 10066
rect 125428 4214 125456 14146
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 123036 3454 124168 3482
rect 119436 2984 119488 2990
rect 119436 2926 119488 2932
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 119448 480 119476 2926
rect 120644 480 120672 2926
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 3454
rect 124232 480 124260 4150
rect 125520 3482 125548 336738
rect 186228 13796 186280 13802
rect 186228 13738 186280 13744
rect 183468 13728 183520 13734
rect 183468 13670 183520 13676
rect 179328 13660 179380 13666
rect 179328 13602 179380 13608
rect 176568 13592 176620 13598
rect 176568 13534 176620 13540
rect 172428 13524 172480 13530
rect 172428 13466 172480 13472
rect 168288 13456 168340 13462
rect 168288 13398 168340 13404
rect 165528 13388 165580 13394
rect 165528 13330 165580 13336
rect 160008 13320 160060 13326
rect 160008 13262 160060 13268
rect 155868 13252 155920 13258
rect 155868 13194 155920 13200
rect 151728 12164 151780 12170
rect 151728 12106 151780 12112
rect 148968 12096 149020 12102
rect 148968 12038 149020 12044
rect 144828 12028 144880 12034
rect 144828 11970 144880 11976
rect 142068 11960 142120 11966
rect 142068 11902 142120 11908
rect 128268 11892 128320 11898
rect 128268 11834 128320 11840
rect 126888 11824 126940 11830
rect 126888 11766 126940 11772
rect 126900 3482 126928 11766
rect 128280 3482 128308 11834
rect 139676 9376 139728 9382
rect 139676 9318 139728 9324
rect 136088 9308 136140 9314
rect 136088 9250 136140 9256
rect 132590 8936 132646 8945
rect 132590 8871 132646 8880
rect 129002 7576 129058 7585
rect 129002 7511 129058 7520
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 7511
rect 131396 6656 131448 6662
rect 131396 6598 131448 6604
rect 130200 5364 130252 5370
rect 130200 5306 130252 5312
rect 130212 480 130240 5306
rect 131408 480 131436 6598
rect 132604 480 132632 8871
rect 134892 7540 134944 7546
rect 134892 7482 134944 7488
rect 133788 5432 133840 5438
rect 133788 5374 133840 5380
rect 133800 480 133828 5374
rect 134904 480 134932 7482
rect 136100 480 136128 9250
rect 138480 7472 138532 7478
rect 138480 7414 138532 7420
rect 137284 5500 137336 5506
rect 137284 5442 137336 5448
rect 137296 480 137324 5442
rect 138492 480 138520 7414
rect 139688 480 139716 9318
rect 141976 7404 142028 7410
rect 141976 7346 142028 7352
rect 140872 4208 140924 4214
rect 140872 4150 140924 4156
rect 140884 480 140912 4150
rect 141988 3482 142016 7346
rect 142080 4214 142108 11902
rect 143448 10056 143500 10062
rect 143448 9998 143500 10004
rect 142068 4208 142120 4214
rect 142068 4150 142120 4156
rect 143460 3482 143488 9998
rect 144840 3482 144868 11970
rect 147588 9988 147640 9994
rect 147588 9930 147640 9936
rect 145656 7336 145708 7342
rect 145656 7278 145708 7284
rect 141988 3454 142108 3482
rect 142080 480 142108 3454
rect 143276 3454 143488 3482
rect 144472 3454 144868 3482
rect 143276 480 143304 3454
rect 144472 480 144500 3454
rect 145668 480 145696 7278
rect 147600 3482 147628 9930
rect 148980 3482 149008 12038
rect 151636 9920 151688 9926
rect 151636 9862 151688 9868
rect 149244 7268 149296 7274
rect 149244 7210 149296 7216
rect 146864 3454 147628 3482
rect 148060 3454 149008 3482
rect 146864 480 146892 3454
rect 148060 480 148088 3454
rect 149256 480 149284 7210
rect 151648 4214 151676 9862
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 150452 480 150480 4150
rect 151740 3482 151768 12106
rect 154488 9852 154540 9858
rect 154488 9794 154540 9800
rect 152740 7200 152792 7206
rect 152740 7142 152792 7148
rect 151556 3454 151768 3482
rect 151556 480 151584 3454
rect 152752 480 152780 7142
rect 154500 3482 154528 9794
rect 155880 3482 155908 13194
rect 158628 9784 158680 9790
rect 158628 9726 158680 9732
rect 156328 7132 156380 7138
rect 156328 7074 156380 7080
rect 153948 3454 154528 3482
rect 155144 3454 155908 3482
rect 153948 480 153976 3454
rect 155144 480 155172 3454
rect 156340 480 156368 7074
rect 158640 3482 158668 9726
rect 159916 7064 159968 7070
rect 159916 7006 159968 7012
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 157536 3454 158668 3482
rect 157536 480 157564 3454
rect 158732 480 158760 4150
rect 159928 480 159956 7006
rect 160020 4214 160048 13262
rect 162768 12232 162820 12238
rect 162768 12174 162820 12180
rect 161388 9716 161440 9722
rect 161388 9658 161440 9664
rect 160008 4208 160060 4214
rect 160008 4150 160060 4156
rect 161400 3482 161428 9658
rect 161124 3454 161428 3482
rect 161124 480 161152 3454
rect 162780 626 162808 12174
rect 163504 6724 163556 6730
rect 163504 6666 163556 6672
rect 162320 598 162808 626
rect 162320 480 162348 598
rect 163516 480 163544 6666
rect 165540 610 165568 13330
rect 166908 12300 166960 12306
rect 166908 12242 166960 12248
rect 166920 610 166948 12242
rect 167092 6792 167144 6798
rect 167092 6734 167144 6740
rect 164700 604 164752 610
rect 164700 546 164752 552
rect 165528 604 165580 610
rect 165528 546 165580 552
rect 165896 604 165948 610
rect 165896 546 165948 552
rect 166908 604 166960 610
rect 166908 546 166960 552
rect 164712 480 164740 546
rect 165908 480 165936 546
rect 167104 480 167132 6734
rect 168300 626 168328 13398
rect 169668 12368 169720 12374
rect 169668 12310 169720 12316
rect 168208 598 168328 626
rect 169680 610 169708 12310
rect 170588 6860 170640 6866
rect 170588 6802 170640 6808
rect 169392 604 169444 610
rect 168208 480 168236 598
rect 169392 546 169444 552
rect 169668 604 169720 610
rect 169668 546 169720 552
rect 169404 480 169432 546
rect 170600 480 170628 6802
rect 172440 3346 172468 13466
rect 173808 12436 173860 12442
rect 173808 12378 173860 12384
rect 173820 3346 173848 12378
rect 176476 11688 176528 11694
rect 176476 11630 176528 11636
rect 174176 6112 174228 6118
rect 174176 6054 174228 6060
rect 171796 3318 172468 3346
rect 172992 3318 173848 3346
rect 171796 480 171824 3318
rect 172992 480 173020 3318
rect 174188 480 174216 6054
rect 175372 4208 175424 4214
rect 175372 4150 175424 4156
rect 175384 480 175412 4150
rect 176488 3482 176516 11630
rect 176580 4214 176608 13534
rect 177764 6044 177816 6050
rect 177764 5986 177816 5992
rect 176568 4208 176620 4214
rect 176568 4150 176620 4156
rect 176488 3454 176608 3482
rect 176580 480 176608 3454
rect 177776 480 177804 5986
rect 179340 3346 179368 13602
rect 180708 11620 180760 11626
rect 180708 11562 180760 11568
rect 180720 3346 180748 11562
rect 181352 5976 181404 5982
rect 181352 5918 181404 5924
rect 178972 3318 179368 3346
rect 180168 3318 180748 3346
rect 178972 480 179000 3318
rect 180168 480 180196 3318
rect 181364 480 181392 5918
rect 183480 610 183508 13670
rect 184848 11552 184900 11558
rect 184848 11494 184900 11500
rect 184860 6066 184888 11494
rect 184768 6038 184888 6066
rect 184768 610 184796 6038
rect 184848 5908 184900 5914
rect 184848 5850 184900 5856
rect 182548 604 182600 610
rect 182548 546 182600 552
rect 183468 604 183520 610
rect 183468 546 183520 552
rect 183744 604 183796 610
rect 183744 546 183796 552
rect 184756 604 184808 610
rect 184756 546 184808 552
rect 182560 480 182588 546
rect 183756 480 183784 546
rect 184860 480 184888 5850
rect 186240 626 186268 13738
rect 190368 13048 190420 13054
rect 190368 12990 190420 12996
rect 187608 11484 187660 11490
rect 187608 11426 187660 11432
rect 186056 598 186268 626
rect 187620 610 187648 11426
rect 188436 5840 188488 5846
rect 188436 5782 188488 5788
rect 187240 604 187292 610
rect 186056 480 186084 598
rect 187240 546 187292 552
rect 187608 604 187660 610
rect 187608 546 187660 552
rect 187252 480 187280 546
rect 188448 480 188476 5782
rect 190380 610 190408 12990
rect 206928 12980 206980 12986
rect 206928 12922 206980 12928
rect 191748 11416 191800 11422
rect 191748 11358 191800 11364
rect 191760 3346 191788 11358
rect 194508 11348 194560 11354
rect 194508 11290 194560 11296
rect 193220 9444 193272 9450
rect 193220 9386 193272 9392
rect 192024 5772 192076 5778
rect 192024 5714 192076 5720
rect 190840 3318 191788 3346
rect 189632 604 189684 610
rect 189632 546 189684 552
rect 190368 604 190420 610
rect 190368 546 190420 552
rect 189644 480 189672 546
rect 190840 480 190868 3318
rect 192036 480 192064 5714
rect 193232 480 193260 9386
rect 194520 3482 194548 11290
rect 198648 11280 198700 11286
rect 198648 11222 198700 11228
rect 196808 9512 196860 9518
rect 196808 9454 196860 9460
rect 195612 5704 195664 5710
rect 195612 5646 195664 5652
rect 194428 3454 194548 3482
rect 194428 480 194456 3454
rect 195624 480 195652 5646
rect 196820 480 196848 9454
rect 198660 3346 198688 11222
rect 203892 9648 203944 9654
rect 203892 9590 203944 9596
rect 200396 9580 200448 9586
rect 200396 9522 200448 9528
rect 199200 5636 199252 5642
rect 199200 5578 199252 5584
rect 198016 3318 198688 3346
rect 198016 480 198044 3318
rect 199212 480 199240 5578
rect 200408 480 200436 9522
rect 202696 5568 202748 5574
rect 202696 5510 202748 5516
rect 201500 4412 201552 4418
rect 201500 4354 201552 4360
rect 201512 480 201540 4354
rect 202708 480 202736 5510
rect 203904 480 203932 9590
rect 205088 4344 205140 4350
rect 205088 4286 205140 4292
rect 205100 480 205128 4286
rect 206940 3346 206968 12922
rect 211068 12912 211120 12918
rect 211068 12854 211120 12860
rect 207480 8900 207532 8906
rect 207480 8842 207532 8848
rect 206296 3318 206968 3346
rect 206296 480 206324 3318
rect 207492 480 207520 8842
rect 210976 8832 211028 8838
rect 210976 8774 211028 8780
rect 208674 4856 208730 4865
rect 208674 4791 208730 4800
rect 208688 480 208716 4791
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 209884 480 209912 4150
rect 210988 3482 211016 8774
rect 211080 4214 211108 12854
rect 213828 12844 213880 12850
rect 213828 12786 213880 12792
rect 212264 4752 212316 4758
rect 212264 4694 212316 4700
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 4694
rect 213840 3346 213868 12786
rect 217968 12776 218020 12782
rect 217968 12718 218020 12724
rect 214656 8764 214708 8770
rect 214656 8706 214708 8712
rect 213472 3318 213868 3346
rect 213472 480 213500 3318
rect 214668 480 214696 8706
rect 215852 4684 215904 4690
rect 215852 4626 215904 4632
rect 215864 480 215892 4626
rect 217980 3346 218008 12718
rect 220728 12708 220780 12714
rect 220728 12650 220780 12656
rect 218152 8696 218204 8702
rect 218152 8638 218204 8644
rect 217060 3318 218008 3346
rect 217060 480 217088 3318
rect 218164 480 218192 8638
rect 219348 4616 219400 4622
rect 219348 4558 219400 4564
rect 219360 480 219388 4558
rect 220740 3346 220768 12650
rect 224868 12640 224920 12646
rect 224868 12582 224920 12588
rect 221740 8628 221792 8634
rect 221740 8570 221792 8576
rect 220556 3318 220768 3346
rect 220556 480 220584 3318
rect 221752 480 221780 8570
rect 222936 4548 222988 4554
rect 222936 4490 222988 4496
rect 222948 480 222976 4490
rect 224880 3346 224908 12582
rect 229008 12572 229060 12578
rect 229008 12514 229060 12520
rect 225328 8560 225380 8566
rect 225328 8502 225380 8508
rect 224144 3318 224908 3346
rect 224144 480 224172 3318
rect 225340 480 225368 8502
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 227720 7608 227772 7614
rect 227720 7550 227772 7556
rect 226524 4480 226576 4486
rect 226524 4422 226576 4428
rect 226536 480 226564 4422
rect 227732 480 227760 7550
rect 228928 480 228956 8434
rect 229020 7614 229048 12514
rect 229008 7608 229060 7614
rect 229008 7550 229060 7556
rect 229112 4962 229140 340054
rect 229100 4956 229152 4962
rect 229100 4898 229152 4904
rect 230112 4888 230164 4894
rect 230112 4830 230164 4836
rect 230124 480 230152 4830
rect 230584 4282 230612 340054
rect 230768 340054 230966 340082
rect 231136 340054 231426 340082
rect 230664 337680 230716 337686
rect 230664 337622 230716 337628
rect 230676 7682 230704 337622
rect 230664 7676 230716 7682
rect 230664 7618 230716 7624
rect 230768 4826 230796 340054
rect 231136 337686 231164 340054
rect 231124 337680 231176 337686
rect 231124 337622 231176 337628
rect 231964 337385 231992 340068
rect 232056 340054 232438 340082
rect 231950 337376 232006 337385
rect 231950 337311 232006 337320
rect 231308 7608 231360 7614
rect 231308 7550 231360 7556
rect 230756 4820 230808 4826
rect 230756 4762 230808 4768
rect 230572 4276 230624 4282
rect 230572 4218 230624 4224
rect 231320 480 231348 7550
rect 232056 3369 232084 340054
rect 232516 337770 232544 340190
rect 232240 337742 232544 337770
rect 232240 321570 232268 337742
rect 232228 321564 232280 321570
rect 232228 321506 232280 321512
rect 232412 321564 232464 321570
rect 232412 321506 232464 321512
rect 232424 311982 232452 321506
rect 232412 311976 232464 311982
rect 232412 311918 232464 311924
rect 232320 311840 232372 311846
rect 232320 311782 232372 311788
rect 232332 205578 232360 311782
rect 232240 205550 232360 205578
rect 232240 196042 232268 205550
rect 232228 196036 232280 196042
rect 232228 195978 232280 195984
rect 232320 195968 232372 195974
rect 232320 195910 232372 195916
rect 232332 186266 232360 195910
rect 232240 186238 232360 186266
rect 232240 176730 232268 186238
rect 232228 176724 232280 176730
rect 232228 176666 232280 176672
rect 232320 176656 232372 176662
rect 232320 176598 232372 176604
rect 232332 166954 232360 176598
rect 232240 166926 232360 166954
rect 232240 162858 232268 166926
rect 232136 162852 232188 162858
rect 232136 162794 232188 162800
rect 232228 162852 232280 162858
rect 232228 162794 232280 162800
rect 232148 153241 232176 162794
rect 232134 153232 232190 153241
rect 232134 153167 232190 153176
rect 232318 153232 232374 153241
rect 232318 153167 232374 153176
rect 232332 143546 232360 153167
rect 232320 143540 232372 143546
rect 232320 143482 232372 143488
rect 232320 133952 232372 133958
rect 232320 133894 232372 133900
rect 232332 124166 232360 133894
rect 232320 124160 232372 124166
rect 232320 124102 232372 124108
rect 232320 114572 232372 114578
rect 232320 114514 232372 114520
rect 232332 104854 232360 114514
rect 232320 104848 232372 104854
rect 232320 104790 232372 104796
rect 232320 95260 232372 95266
rect 232320 95202 232372 95208
rect 232332 85542 232360 95202
rect 232320 85536 232372 85542
rect 232320 85478 232372 85484
rect 232320 75948 232372 75954
rect 232320 75890 232372 75896
rect 232332 67810 232360 75890
rect 232240 67782 232360 67810
rect 232240 67674 232268 67782
rect 232240 67646 232360 67674
rect 232332 66230 232360 67646
rect 232320 66224 232372 66230
rect 232320 66166 232372 66172
rect 232320 56636 232372 56642
rect 232320 56578 232372 56584
rect 232332 48385 232360 56578
rect 232318 48376 232374 48385
rect 232318 48311 232374 48320
rect 232318 47968 232374 47977
rect 232318 47903 232374 47912
rect 232332 38690 232360 47903
rect 232320 38684 232372 38690
rect 232320 38626 232372 38632
rect 232504 38548 232556 38554
rect 232504 38490 232556 38496
rect 232516 31634 232544 38490
rect 232424 31606 232544 31634
rect 232424 28966 232452 31606
rect 232228 28960 232280 28966
rect 232228 28902 232280 28908
rect 232412 28960 232464 28966
rect 232412 28902 232464 28908
rect 232240 12458 232268 28902
rect 232240 12430 232360 12458
rect 232332 12322 232360 12430
rect 232148 12294 232360 12322
rect 232148 5030 232176 12294
rect 232504 8424 232556 8430
rect 232504 8366 232556 8372
rect 232136 5024 232188 5030
rect 232136 4966 232188 4972
rect 232042 3360 232098 3369
rect 232042 3295 232098 3304
rect 232516 480 232544 8366
rect 233436 7002 233464 340068
rect 233528 340054 233910 340082
rect 233528 337414 233556 340054
rect 234356 337482 234384 340068
rect 234724 340054 234922 340082
rect 235000 340054 235382 340082
rect 235644 340054 235842 340082
rect 236394 340054 236500 340082
rect 234344 337476 234396 337482
rect 234344 337418 234396 337424
rect 233516 337408 233568 337414
rect 233516 337350 233568 337356
rect 233884 337408 233936 337414
rect 233884 337350 233936 337356
rect 233896 9110 233924 337350
rect 233884 9104 233936 9110
rect 233884 9046 233936 9052
rect 233424 6996 233476 7002
rect 233424 6938 233476 6944
rect 234724 5098 234752 340054
rect 235000 334642 235028 340054
rect 234816 334614 235028 334642
rect 234816 8974 234844 334614
rect 235644 334558 235672 340054
rect 236184 335708 236236 335714
rect 236184 335650 236236 335656
rect 236092 335640 236144 335646
rect 236092 335582 236144 335588
rect 234988 334552 235040 334558
rect 234988 334494 235040 334500
rect 235632 334552 235684 334558
rect 235632 334494 235684 334500
rect 235000 41290 235028 334494
rect 235000 41262 235120 41290
rect 235092 19394 235120 41262
rect 235000 19366 235120 19394
rect 235000 14498 235028 19366
rect 234908 14470 235028 14498
rect 234804 8968 234856 8974
rect 234804 8910 234856 8916
rect 234804 7676 234856 7682
rect 234804 7618 234856 7624
rect 234712 5092 234764 5098
rect 234712 5034 234764 5040
rect 233700 4820 233752 4826
rect 233700 4762 233752 4768
rect 233712 480 233740 4762
rect 234816 480 234844 7618
rect 234908 3466 234936 14470
rect 236000 8968 236052 8974
rect 236000 8910 236052 8916
rect 234896 3460 234948 3466
rect 234896 3402 234948 3408
rect 236012 480 236040 8910
rect 236104 5166 236132 335582
rect 236196 9042 236224 335650
rect 236472 321586 236500 340054
rect 236564 340054 236854 340082
rect 237024 340054 237314 340082
rect 236564 335646 236592 340054
rect 237024 335714 237052 340054
rect 237852 337550 237880 340068
rect 237840 337544 237892 337550
rect 237840 337486 237892 337492
rect 238312 337482 238340 340068
rect 238786 340054 238892 340082
rect 238300 337476 238352 337482
rect 238300 337418 238352 337424
rect 237012 335708 237064 335714
rect 237012 335650 237064 335656
rect 236552 335640 236604 335646
rect 236552 335582 236604 335588
rect 236288 321558 236500 321586
rect 236288 309369 236316 321558
rect 236274 309360 236330 309369
rect 236274 309295 236330 309304
rect 236274 309224 236330 309233
rect 236274 309159 236330 309168
rect 236288 309126 236316 309159
rect 236276 309120 236328 309126
rect 236276 309062 236328 309068
rect 236460 299532 236512 299538
rect 236460 299474 236512 299480
rect 236472 292602 236500 299474
rect 236276 292596 236328 292602
rect 236276 292538 236328 292544
rect 236460 292596 236512 292602
rect 236460 292538 236512 292544
rect 236288 282946 236316 292538
rect 236276 282940 236328 282946
rect 236276 282882 236328 282888
rect 236460 282804 236512 282810
rect 236460 282746 236512 282752
rect 236472 280158 236500 282746
rect 236460 280152 236512 280158
rect 236460 280094 236512 280100
rect 236276 270564 236328 270570
rect 236276 270506 236328 270512
rect 236288 270473 236316 270506
rect 236274 270464 236330 270473
rect 236274 270399 236330 270408
rect 236458 260944 236514 260953
rect 236458 260879 236514 260888
rect 236472 260846 236500 260879
rect 236460 260840 236512 260846
rect 236460 260782 236512 260788
rect 236276 251252 236328 251258
rect 236276 251194 236328 251200
rect 236288 251161 236316 251194
rect 236274 251152 236330 251161
rect 236274 251087 236330 251096
rect 236550 251152 236606 251161
rect 236550 251087 236606 251096
rect 236564 241534 236592 251087
rect 236552 241528 236604 241534
rect 236552 241470 236604 241476
rect 236644 241528 236696 241534
rect 236644 241470 236696 241476
rect 236656 232121 236684 241470
rect 236642 232112 236698 232121
rect 236642 232047 236698 232056
rect 236274 231976 236330 231985
rect 236274 231911 236330 231920
rect 236288 225010 236316 231911
rect 236276 225004 236328 225010
rect 236276 224946 236328 224952
rect 236460 224868 236512 224874
rect 236460 224810 236512 224816
rect 236472 222193 236500 224810
rect 236458 222184 236514 222193
rect 236458 222119 236514 222128
rect 236274 212664 236330 212673
rect 236274 212599 236330 212608
rect 236288 212537 236316 212599
rect 236274 212528 236330 212537
rect 236274 212463 236330 212472
rect 236550 212528 236606 212537
rect 236550 212463 236606 212472
rect 236564 203017 236592 212463
rect 236550 203008 236606 203017
rect 236550 202943 236606 202952
rect 236274 193352 236330 193361
rect 236274 193287 236330 193296
rect 236288 193225 236316 193287
rect 236274 193216 236330 193225
rect 236274 193151 236330 193160
rect 236550 193216 236606 193225
rect 236550 193151 236606 193160
rect 236472 183598 236500 183629
rect 236564 183598 236592 193151
rect 236460 183592 236512 183598
rect 236552 183592 236604 183598
rect 236512 183540 236552 183546
rect 236604 183540 236684 183546
rect 236460 183534 236684 183540
rect 236472 183518 236684 183534
rect 236656 173942 236684 183518
rect 236276 173936 236328 173942
rect 236276 173878 236328 173884
rect 236644 173936 236696 173942
rect 236644 173878 236696 173884
rect 236288 166954 236316 173878
rect 236288 166926 236500 166954
rect 236472 154601 236500 166926
rect 236274 154592 236330 154601
rect 236274 154527 236330 154536
rect 236458 154592 236514 154601
rect 236458 154527 236514 154536
rect 236288 147642 236316 154527
rect 236288 147614 236500 147642
rect 236472 135289 236500 147614
rect 236274 135280 236330 135289
rect 236274 135215 236330 135224
rect 236458 135280 236514 135289
rect 236458 135215 236514 135224
rect 236288 128330 236316 135215
rect 236288 128302 236500 128330
rect 236472 115977 236500 128302
rect 236274 115968 236330 115977
rect 236274 115903 236330 115912
rect 236458 115968 236514 115977
rect 236458 115903 236514 115912
rect 236288 109018 236316 115903
rect 236288 108990 236500 109018
rect 236472 106282 236500 108990
rect 236460 106276 236512 106282
rect 236460 106218 236512 106224
rect 236644 106276 236696 106282
rect 236644 106218 236696 106224
rect 236656 96665 236684 106218
rect 236274 96656 236330 96665
rect 236274 96591 236330 96600
rect 236642 96656 236698 96665
rect 236642 96591 236698 96600
rect 236288 89706 236316 96591
rect 236288 89678 236500 89706
rect 236472 86970 236500 89678
rect 236460 86964 236512 86970
rect 236460 86906 236512 86912
rect 236276 77444 236328 77450
rect 236276 77386 236328 77392
rect 236288 67590 236316 77386
rect 236276 67584 236328 67590
rect 236276 67526 236328 67532
rect 236368 67584 236420 67590
rect 236368 67526 236420 67532
rect 236380 66230 236408 67526
rect 236368 66224 236420 66230
rect 236368 66166 236420 66172
rect 236276 56636 236328 56642
rect 236276 56578 236328 56584
rect 236288 48278 236316 56578
rect 236276 48272 236328 48278
rect 236276 48214 236328 48220
rect 236276 38684 236328 38690
rect 236276 38626 236328 38632
rect 236288 38554 236316 38626
rect 236276 38548 236328 38554
rect 236276 38490 236328 38496
rect 236368 31680 236420 31686
rect 236368 31622 236420 31628
rect 236380 28966 236408 31622
rect 236368 28960 236420 28966
rect 236368 28902 236420 28908
rect 236460 22772 236512 22778
rect 236460 22714 236512 22720
rect 236472 17950 236500 22714
rect 236460 17944 236512 17950
rect 236460 17886 236512 17892
rect 236184 9036 236236 9042
rect 236184 8978 236236 8984
rect 236276 8356 236328 8362
rect 236276 8298 236328 8304
rect 236092 5160 236144 5166
rect 236092 5102 236144 5108
rect 236288 3534 236316 8298
rect 238864 7750 238892 340054
rect 238956 340054 239338 340082
rect 239508 340054 239798 340082
rect 240258 340054 240364 340082
rect 238956 11762 238984 340054
rect 239508 331242 239536 340054
rect 239140 331214 239536 331242
rect 239140 313970 239168 331214
rect 239140 313942 239352 313970
rect 239324 299538 239352 313942
rect 239128 299532 239180 299538
rect 239128 299474 239180 299480
rect 239312 299532 239364 299538
rect 239312 299474 239364 299480
rect 239140 292618 239168 299474
rect 239048 292590 239168 292618
rect 239048 292534 239076 292590
rect 239036 292528 239088 292534
rect 239036 292470 239088 292476
rect 239220 292528 239272 292534
rect 239220 292470 239272 292476
rect 239232 280242 239260 292470
rect 239140 280214 239260 280242
rect 239140 280158 239168 280214
rect 239128 280152 239180 280158
rect 239128 280094 239180 280100
rect 239220 270564 239272 270570
rect 239220 270506 239272 270512
rect 239232 263514 239260 270506
rect 239140 263486 239260 263514
rect 239140 260846 239168 263486
rect 239128 260840 239180 260846
rect 239128 260782 239180 260788
rect 239220 251252 239272 251258
rect 239220 251194 239272 251200
rect 239232 244202 239260 251194
rect 239140 244174 239260 244202
rect 239140 236722 239168 244174
rect 239140 236694 239260 236722
rect 239232 224890 239260 236694
rect 239140 224862 239260 224890
rect 239140 217410 239168 224862
rect 239140 217382 239260 217410
rect 239232 205578 239260 217382
rect 239140 205550 239260 205578
rect 239140 202842 239168 205550
rect 239128 202836 239180 202842
rect 239128 202778 239180 202784
rect 239220 202836 239272 202842
rect 239220 202778 239272 202784
rect 239232 186266 239260 202778
rect 239140 186238 239260 186266
rect 239140 183530 239168 186238
rect 239128 183524 239180 183530
rect 239128 183466 239180 183472
rect 239220 183524 239272 183530
rect 239220 183466 239272 183472
rect 239232 166954 239260 183466
rect 239140 166926 239260 166954
rect 239140 164218 239168 166926
rect 239128 164212 239180 164218
rect 239128 164154 239180 164160
rect 239220 164212 239272 164218
rect 239220 164154 239272 164160
rect 239232 147642 239260 164154
rect 239140 147614 239260 147642
rect 239140 138038 239168 147614
rect 239128 138032 239180 138038
rect 239128 137974 239180 137980
rect 239036 137964 239088 137970
rect 239036 137906 239088 137912
rect 239048 135289 239076 137906
rect 239034 135280 239090 135289
rect 239034 135215 239090 135224
rect 239218 135280 239274 135289
rect 239218 135215 239274 135224
rect 239232 128330 239260 135215
rect 239140 128302 239260 128330
rect 239140 125594 239168 128302
rect 239128 125588 239180 125594
rect 239128 125530 239180 125536
rect 239128 116000 239180 116006
rect 239128 115942 239180 115948
rect 239140 106282 239168 115942
rect 239128 106276 239180 106282
rect 239128 106218 239180 106224
rect 239312 106276 239364 106282
rect 239312 106218 239364 106224
rect 239324 96665 239352 106218
rect 239126 96656 239182 96665
rect 239126 96591 239182 96600
rect 239310 96656 239366 96665
rect 239310 96591 239366 96600
rect 239140 70514 239168 96591
rect 239128 70508 239180 70514
rect 239128 70450 239180 70456
rect 239128 67652 239180 67658
rect 239128 67594 239180 67600
rect 239140 58070 239168 67594
rect 239128 58064 239180 58070
rect 239128 58006 239180 58012
rect 239036 56636 239088 56642
rect 239036 56578 239088 56584
rect 239048 53242 239076 56578
rect 239036 53236 239088 53242
rect 239036 53178 239088 53184
rect 239128 48340 239180 48346
rect 239128 48282 239180 48288
rect 239140 42090 239168 48282
rect 239128 42084 239180 42090
rect 239128 42026 239180 42032
rect 240138 29200 240194 29209
rect 240138 29135 240140 29144
rect 240192 29135 240194 29144
rect 240140 29106 240192 29112
rect 239036 29028 239088 29034
rect 239036 28970 239088 28976
rect 238944 11756 238996 11762
rect 238944 11698 238996 11704
rect 239048 9738 239076 28970
rect 238956 9710 239076 9738
rect 238956 8362 238984 9710
rect 239588 9036 239640 9042
rect 239588 8978 239640 8984
rect 238944 8356 238996 8362
rect 238944 8298 238996 8304
rect 239036 8356 239088 8362
rect 239036 8298 239088 8304
rect 238852 7744 238904 7750
rect 238852 7686 238904 7692
rect 238392 6996 238444 7002
rect 238392 6938 238444 6944
rect 237196 4956 237248 4962
rect 237196 4898 237248 4904
rect 236276 3528 236328 3534
rect 236276 3470 236328 3476
rect 237208 480 237236 4898
rect 238404 480 238432 6938
rect 239048 3602 239076 8298
rect 239036 3596 239088 3602
rect 239036 3538 239088 3544
rect 239600 480 239628 8978
rect 240336 3670 240364 340054
rect 240428 340054 240810 340082
rect 240428 7818 240456 340054
rect 241256 337414 241284 340068
rect 241716 337618 241744 340068
rect 241808 340054 242282 340082
rect 242360 340054 242742 340082
rect 243096 340054 243202 340082
rect 243464 340054 243754 340082
rect 241704 337612 241756 337618
rect 241704 337554 241756 337560
rect 241244 337408 241296 337414
rect 241244 337350 241296 337356
rect 241612 335640 241664 335646
rect 241612 335582 241664 335588
rect 241624 13122 241652 335582
rect 241612 13116 241664 13122
rect 241612 13058 241664 13064
rect 241808 7886 241836 340054
rect 242360 335646 242388 340054
rect 242348 335640 242400 335646
rect 242348 335582 242400 335588
rect 242992 332104 243044 332110
rect 242992 332046 243044 332052
rect 243004 7954 243032 332046
rect 242992 7948 243044 7954
rect 242992 7890 243044 7896
rect 241796 7880 241848 7886
rect 241796 7822 241848 7828
rect 240416 7812 240468 7818
rect 240416 7754 240468 7760
rect 241980 7744 242032 7750
rect 241980 7686 242032 7692
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 240324 3664 240376 3670
rect 240324 3606 240376 3612
rect 240796 480 240824 4966
rect 241992 480 242020 7686
rect 243096 3738 243124 340054
rect 243464 332110 243492 340054
rect 244200 337822 244228 340068
rect 244188 337816 244240 337822
rect 244188 337758 244240 337764
rect 244660 337550 244688 340068
rect 244648 337544 244700 337550
rect 244648 337486 244700 337492
rect 244752 335594 244780 340190
rect 245686 340054 245792 340082
rect 244476 335566 244780 335594
rect 243452 332104 243504 332110
rect 243452 332046 243504 332052
rect 244476 311846 244504 335566
rect 244464 311840 244516 311846
rect 244464 311782 244516 311788
rect 244464 309188 244516 309194
rect 244464 309130 244516 309136
rect 244476 292618 244504 309130
rect 244384 292590 244504 292618
rect 244384 292482 244412 292590
rect 244384 292454 244504 292482
rect 244476 273306 244504 292454
rect 244384 273278 244504 273306
rect 244384 273170 244412 273278
rect 244384 273142 244504 273170
rect 244476 259457 244504 273142
rect 244462 259448 244518 259457
rect 244462 259383 244518 259392
rect 244646 259448 244702 259457
rect 244646 259383 244702 259392
rect 244660 254538 244688 259383
rect 244476 254510 244688 254538
rect 244476 241505 244504 254510
rect 244278 241496 244334 241505
rect 244278 241431 244334 241440
rect 244462 241496 244518 241505
rect 244462 241431 244518 241440
rect 244292 231878 244320 241431
rect 244280 231872 244332 231878
rect 244280 231814 244332 231820
rect 244464 231872 244516 231878
rect 244464 231814 244516 231820
rect 244476 222193 244504 231814
rect 244278 222184 244334 222193
rect 244278 222119 244334 222128
rect 244462 222184 244518 222193
rect 244462 222119 244518 222128
rect 244292 212566 244320 222119
rect 244280 212560 244332 212566
rect 244280 212502 244332 212508
rect 244464 212560 244516 212566
rect 244464 212502 244516 212508
rect 244476 202881 244504 212502
rect 244278 202872 244334 202881
rect 244278 202807 244334 202816
rect 244462 202872 244518 202881
rect 244462 202807 244518 202816
rect 244292 193254 244320 202807
rect 244280 193248 244332 193254
rect 244280 193190 244332 193196
rect 244464 193248 244516 193254
rect 244464 193190 244516 193196
rect 244476 176746 244504 193190
rect 244384 176718 244504 176746
rect 244384 176610 244412 176718
rect 244384 176582 244504 176610
rect 244476 164218 244504 176582
rect 244280 164212 244332 164218
rect 244280 164154 244332 164160
rect 244464 164212 244516 164218
rect 244464 164154 244516 164160
rect 244292 154601 244320 164154
rect 244278 154592 244334 154601
rect 244278 154527 244334 154536
rect 244462 154592 244518 154601
rect 244462 154527 244518 154536
rect 244476 144906 244504 154527
rect 244280 144900 244332 144906
rect 244280 144842 244332 144848
rect 244464 144900 244516 144906
rect 244464 144842 244516 144848
rect 244292 135289 244320 144842
rect 244278 135280 244334 135289
rect 244278 135215 244334 135224
rect 244462 135280 244518 135289
rect 244462 135215 244518 135224
rect 244476 118810 244504 135215
rect 244384 118782 244504 118810
rect 244384 118674 244412 118782
rect 244384 118646 244504 118674
rect 244476 106264 244504 118646
rect 244384 106236 244504 106264
rect 244384 99414 244412 106236
rect 244372 99408 244424 99414
rect 244372 99350 244424 99356
rect 244464 99340 244516 99346
rect 244464 99282 244516 99288
rect 244476 70514 244504 99282
rect 244464 70508 244516 70514
rect 244464 70450 244516 70456
rect 244464 67652 244516 67658
rect 244464 67594 244516 67600
rect 244476 58002 244504 67594
rect 244464 57996 244516 58002
rect 244464 57938 244516 57944
rect 244556 57860 244608 57866
rect 244556 57802 244608 57808
rect 244568 56574 244596 57802
rect 244556 56568 244608 56574
rect 244556 56510 244608 56516
rect 244556 48204 244608 48210
rect 244556 48146 244608 48152
rect 244568 46918 244596 48146
rect 244556 46912 244608 46918
rect 244556 46854 244608 46860
rect 244556 37324 244608 37330
rect 244556 37266 244608 37272
rect 244568 29050 244596 37266
rect 244476 29022 244596 29050
rect 244476 22658 244504 29022
rect 244384 22630 244504 22658
rect 244384 18034 244412 22630
rect 244384 18006 244596 18034
rect 244568 17950 244596 18006
rect 244556 17944 244608 17950
rect 244556 17886 244608 17892
rect 243176 9104 243228 9110
rect 243176 9046 243228 9052
rect 243084 3732 243136 3738
rect 243084 3674 243136 3680
rect 243188 480 243216 9046
rect 244372 8356 244424 8362
rect 244372 8298 244424 8304
rect 244384 8022 244412 8298
rect 244372 8016 244424 8022
rect 244372 7958 244424 7964
rect 245568 7812 245620 7818
rect 245568 7754 245620 7760
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 244384 480 244412 5034
rect 245580 480 245608 7754
rect 245764 3806 245792 340054
rect 245948 340054 246146 340082
rect 245844 335504 245896 335510
rect 245844 335446 245896 335452
rect 245856 8090 245884 335446
rect 245844 8084 245896 8090
rect 245844 8026 245896 8032
rect 245948 3874 245976 340054
rect 246684 335510 246712 340068
rect 247144 337890 247172 340068
rect 247604 337958 247632 340068
rect 247592 337952 247644 337958
rect 247592 337894 247644 337900
rect 247132 337884 247184 337890
rect 247132 337826 247184 337832
rect 247684 336524 247736 336530
rect 247684 336466 247736 336472
rect 246672 335504 246724 335510
rect 246672 335446 246724 335452
rect 247132 334212 247184 334218
rect 247132 334154 247184 334160
rect 247144 331106 247172 334154
rect 247144 331078 247264 331106
rect 247236 302274 247264 331078
rect 247144 302246 247264 302274
rect 247144 302138 247172 302246
rect 247144 302110 247264 302138
rect 247236 282962 247264 302110
rect 247144 282934 247264 282962
rect 247144 282826 247172 282934
rect 247144 282798 247264 282826
rect 247236 263650 247264 282798
rect 247144 263622 247264 263650
rect 247144 263514 247172 263622
rect 247144 263486 247264 263514
rect 247236 244338 247264 263486
rect 247144 244310 247264 244338
rect 247144 244202 247172 244310
rect 247144 244174 247264 244202
rect 247236 225026 247264 244174
rect 247144 224998 247264 225026
rect 247144 224890 247172 224998
rect 247144 224862 247264 224890
rect 247236 205714 247264 224862
rect 247144 205686 247264 205714
rect 247144 205578 247172 205686
rect 247144 205550 247264 205578
rect 247236 186402 247264 205550
rect 247144 186374 247264 186402
rect 247144 186266 247172 186374
rect 247144 186238 247264 186266
rect 247236 167090 247264 186238
rect 247144 167062 247264 167090
rect 247144 166954 247172 167062
rect 247144 166926 247264 166954
rect 247236 164200 247264 166926
rect 247236 164172 247356 164200
rect 247328 154630 247356 164172
rect 247224 154624 247276 154630
rect 247224 154566 247276 154572
rect 247316 154624 247368 154630
rect 247316 154566 247368 154572
rect 247236 147778 247264 154566
rect 247236 147750 247356 147778
rect 247328 144945 247356 147750
rect 247130 144936 247186 144945
rect 247314 144936 247370 144945
rect 247130 144871 247132 144880
rect 247184 144871 247186 144880
rect 247224 144900 247276 144906
rect 247132 144842 247184 144848
rect 247314 144871 247370 144880
rect 247224 144842 247276 144848
rect 247236 128466 247264 144842
rect 247144 128438 247264 128466
rect 247144 128330 247172 128438
rect 247144 128302 247264 128330
rect 247236 109070 247264 128302
rect 247224 109064 247276 109070
rect 247224 109006 247276 109012
rect 247224 106344 247276 106350
rect 247224 106286 247276 106292
rect 247236 96694 247264 106286
rect 247132 96688 247184 96694
rect 247132 96630 247184 96636
rect 247224 96688 247276 96694
rect 247224 96630 247276 96636
rect 247144 95198 247172 96630
rect 247132 95192 247184 95198
rect 247132 95134 247184 95140
rect 247224 85604 247276 85610
rect 247224 85546 247276 85552
rect 247236 60636 247264 85546
rect 247144 60608 247264 60636
rect 247144 60466 247172 60608
rect 247144 60438 247264 60466
rect 247236 51134 247264 60438
rect 247224 51128 247276 51134
rect 247224 51070 247276 51076
rect 247132 51060 247184 51066
rect 247132 51002 247184 51008
rect 247144 38690 247172 51002
rect 247132 38684 247184 38690
rect 247132 38626 247184 38632
rect 247224 38684 247276 38690
rect 247224 38626 247276 38632
rect 247236 29050 247264 38626
rect 247144 29022 247264 29050
rect 247144 27606 247172 29022
rect 247132 27600 247184 27606
rect 247132 27542 247184 27548
rect 247132 18012 247184 18018
rect 247132 17954 247184 17960
rect 247144 9178 247172 17954
rect 247132 9172 247184 9178
rect 247132 9114 247184 9120
rect 246764 8356 246816 8362
rect 246764 8298 246816 8304
rect 245936 3868 245988 3874
rect 245936 3810 245988 3816
rect 245752 3800 245804 3806
rect 245752 3742 245804 3748
rect 246776 480 246804 8298
rect 247696 3942 247724 336466
rect 248156 334218 248184 340068
rect 248616 336530 248644 340068
rect 248708 340054 249090 340082
rect 248604 336524 248656 336530
rect 248604 336466 248656 336472
rect 248512 336116 248564 336122
rect 248512 336058 248564 336064
rect 248144 334212 248196 334218
rect 248144 334154 248196 334160
rect 248524 5234 248552 336058
rect 248512 5228 248564 5234
rect 248512 5170 248564 5176
rect 247960 5160 248012 5166
rect 247960 5102 248012 5108
rect 247684 3936 247736 3942
rect 247684 3878 247736 3884
rect 247972 480 248000 5102
rect 248708 4010 248736 340054
rect 249064 337748 249116 337754
rect 249064 337690 249116 337696
rect 249076 4078 249104 337690
rect 249536 336122 249564 340068
rect 249904 340054 250102 340082
rect 249524 336116 249576 336122
rect 249524 336058 249576 336064
rect 249154 334248 249210 334257
rect 249154 334183 249210 334192
rect 249168 328545 249196 334183
rect 249154 328536 249210 328545
rect 249154 328471 249210 328480
rect 249154 322280 249210 322289
rect 249154 322215 249210 322224
rect 249168 317665 249196 322215
rect 249154 317656 249210 317665
rect 249154 317591 249210 317600
rect 249246 298072 249302 298081
rect 249246 298007 249302 298016
rect 249260 288561 249288 298007
rect 249246 288552 249302 288561
rect 249246 288487 249302 288496
rect 249246 288416 249302 288425
rect 249246 288351 249302 288360
rect 249260 279041 249288 288351
rect 249246 279032 249302 279041
rect 249246 278967 249302 278976
rect 249430 277400 249486 277409
rect 249430 277335 249486 277344
rect 249444 267889 249472 277335
rect 249430 267880 249486 267889
rect 249430 267815 249486 267824
rect 249246 212528 249302 212537
rect 249246 212463 249302 212472
rect 249260 205465 249288 212463
rect 249246 205456 249302 205465
rect 249246 205391 249302 205400
rect 249614 202872 249670 202881
rect 249614 202807 249670 202816
rect 249628 196625 249656 202807
rect 249614 196616 249670 196625
rect 249614 196551 249670 196560
rect 249246 191584 249302 191593
rect 249246 191519 249302 191528
rect 249260 182209 249288 191519
rect 249246 182200 249302 182209
rect 249246 182135 249302 182144
rect 249430 180568 249486 180577
rect 249430 180503 249486 180512
rect 249444 173913 249472 180503
rect 249430 173904 249486 173913
rect 249430 173839 249486 173848
rect 249708 29164 249760 29170
rect 249708 29106 249760 29112
rect 249720 29073 249748 29106
rect 249706 29064 249762 29073
rect 249706 28999 249762 29008
rect 249904 9246 249932 340054
rect 250548 337754 250576 340068
rect 250640 340054 251022 340082
rect 251284 340054 251574 340082
rect 250536 337748 250588 337754
rect 250536 337690 250588 337696
rect 250444 337408 250496 337414
rect 250444 337350 250496 337356
rect 250168 328500 250220 328506
rect 250168 328442 250220 328448
rect 250180 314022 250208 328442
rect 250168 314016 250220 314022
rect 250168 313958 250220 313964
rect 250168 313880 250220 313886
rect 250168 313822 250220 313828
rect 250180 292618 250208 313822
rect 250088 292590 250208 292618
rect 250088 289814 250116 292590
rect 250076 289808 250128 289814
rect 250076 289750 250128 289756
rect 250352 289808 250404 289814
rect 250352 289750 250404 289756
rect 250364 288425 250392 289750
rect 250074 288416 250130 288425
rect 250074 288351 250130 288360
rect 250350 288416 250406 288425
rect 250350 288351 250406 288360
rect 250088 278798 250116 288351
rect 250076 278792 250128 278798
rect 250076 278734 250128 278740
rect 250168 278792 250220 278798
rect 250168 278734 250220 278740
rect 250180 273358 250208 278734
rect 250168 273352 250220 273358
rect 250168 273294 250220 273300
rect 250076 273216 250128 273222
rect 250076 273158 250128 273164
rect 250088 269074 250116 273158
rect 250076 269068 250128 269074
rect 250076 269010 250128 269016
rect 250168 259480 250220 259486
rect 250168 259422 250220 259428
rect 250180 259350 250208 259422
rect 250168 259344 250220 259350
rect 250168 259286 250220 259292
rect 250352 251116 250404 251122
rect 250352 251058 250404 251064
rect 250364 231878 250392 251058
rect 250076 231872 250128 231878
rect 250076 231814 250128 231820
rect 250352 231872 250404 231878
rect 250352 231814 250404 231820
rect 250088 227202 250116 231814
rect 250088 227174 250392 227202
rect 250364 212566 250392 227174
rect 250076 212560 250128 212566
rect 250076 212502 250128 212508
rect 250352 212560 250404 212566
rect 250352 212502 250404 212508
rect 250088 211138 250116 212502
rect 250076 211132 250128 211138
rect 250076 211074 250128 211080
rect 250260 211132 250312 211138
rect 250260 211074 250312 211080
rect 250272 201498 250300 211074
rect 250272 201482 250392 201498
rect 250076 201476 250128 201482
rect 250272 201476 250404 201482
rect 250272 201470 250352 201476
rect 250076 201418 250128 201424
rect 250352 201418 250404 201424
rect 250088 200122 250116 201418
rect 250076 200116 250128 200122
rect 250076 200058 250128 200064
rect 250076 186312 250128 186318
rect 250076 186254 250128 186260
rect 250088 177342 250116 186254
rect 250076 177336 250128 177342
rect 250076 177278 250128 177284
rect 250352 177336 250404 177342
rect 250352 177278 250404 177284
rect 250364 154737 250392 177278
rect 250350 154728 250406 154737
rect 250350 154663 250406 154672
rect 250074 154592 250130 154601
rect 250074 154527 250130 154536
rect 250088 149682 250116 154527
rect 249996 149654 250116 149682
rect 249996 144922 250024 149654
rect 249996 144894 250300 144922
rect 250272 135425 250300 144894
rect 250258 135416 250314 135425
rect 250258 135351 250314 135360
rect 250074 135280 250130 135289
rect 250074 135215 250130 135224
rect 250088 128382 250116 135215
rect 250076 128376 250128 128382
rect 250076 128318 250128 128324
rect 250168 128308 250220 128314
rect 250168 128250 250220 128256
rect 250180 124166 250208 128250
rect 250168 124160 250220 124166
rect 250168 124102 250220 124108
rect 249984 114572 250036 114578
rect 249984 114514 250036 114520
rect 249996 109018 250024 114514
rect 249996 108990 250208 109018
rect 250180 96694 250208 108990
rect 250076 96688 250128 96694
rect 250076 96630 250128 96636
rect 250168 96688 250220 96694
rect 250168 96630 250220 96636
rect 250088 91746 250116 96630
rect 250088 91718 250208 91746
rect 250180 86952 250208 91718
rect 250088 86924 250208 86952
rect 250088 67590 250116 86924
rect 250076 67584 250128 67590
rect 250076 67526 250128 67532
rect 250168 57996 250220 58002
rect 250168 57938 250220 57944
rect 250180 48278 250208 57938
rect 250168 48272 250220 48278
rect 250168 48214 250220 48220
rect 250260 48272 250312 48278
rect 250260 48214 250312 48220
rect 250272 38214 250300 48214
rect 250260 38208 250312 38214
rect 250260 38150 250312 38156
rect 250260 38072 250312 38078
rect 250260 38014 250312 38020
rect 250272 29050 250300 38014
rect 250180 29022 250300 29050
rect 250180 27606 250208 29022
rect 250168 27600 250220 27606
rect 250168 27542 250220 27548
rect 249984 18012 250036 18018
rect 249984 17954 250036 17960
rect 249892 9240 249944 9246
rect 249892 9182 249944 9188
rect 249156 7880 249208 7886
rect 249156 7822 249208 7828
rect 249064 4072 249116 4078
rect 249064 4014 249116 4020
rect 248696 4004 248748 4010
rect 248696 3946 248748 3952
rect 249168 480 249196 7822
rect 249996 6225 250024 17954
rect 250352 9172 250404 9178
rect 250352 9114 250404 9120
rect 249982 6216 250038 6225
rect 249982 6151 250038 6160
rect 250364 480 250392 9114
rect 250456 4146 250484 337350
rect 250640 334490 250668 340054
rect 250628 334484 250680 334490
rect 250628 334426 250680 334432
rect 251178 87136 251234 87145
rect 251178 87071 251180 87080
rect 251232 87071 251234 87080
rect 251180 87042 251232 87048
rect 251180 37256 251232 37262
rect 251180 37198 251232 37204
rect 251192 27713 251220 37198
rect 251178 27704 251234 27713
rect 251178 27639 251234 27648
rect 251284 10334 251312 340054
rect 252020 338026 252048 340068
rect 252008 338020 252060 338026
rect 252008 337962 252060 337968
rect 252480 337754 252508 340068
rect 252664 340054 253046 340082
rect 251456 337748 251508 337754
rect 251456 337690 251508 337696
rect 252468 337748 252520 337754
rect 252468 337690 252520 337696
rect 251468 321638 251496 337690
rect 251824 336728 251876 336734
rect 251824 336670 251876 336676
rect 251456 321632 251508 321638
rect 251456 321574 251508 321580
rect 251548 321428 251600 321434
rect 251548 321370 251600 321376
rect 251560 294710 251588 321370
rect 251548 294704 251600 294710
rect 251548 294646 251600 294652
rect 251456 289876 251508 289882
rect 251456 289818 251508 289824
rect 251468 280158 251496 289818
rect 251456 280152 251508 280158
rect 251456 280094 251508 280100
rect 251456 270564 251508 270570
rect 251456 270506 251508 270512
rect 251468 260846 251496 270506
rect 251456 260840 251508 260846
rect 251456 260782 251508 260788
rect 251456 251252 251508 251258
rect 251456 251194 251508 251200
rect 251468 241505 251496 251194
rect 251454 241496 251510 241505
rect 251454 241431 251510 241440
rect 251638 241496 251694 241505
rect 251638 241431 251694 241440
rect 251652 231878 251680 241431
rect 251456 231872 251508 231878
rect 251456 231814 251508 231820
rect 251640 231872 251692 231878
rect 251640 231814 251692 231820
rect 251468 222193 251496 231814
rect 251454 222184 251510 222193
rect 251454 222119 251510 222128
rect 251638 222184 251694 222193
rect 251638 222119 251694 222128
rect 251652 212566 251680 222119
rect 251456 212560 251508 212566
rect 251456 212502 251508 212508
rect 251640 212560 251692 212566
rect 251640 212502 251692 212508
rect 251468 202881 251496 212502
rect 251454 202872 251510 202881
rect 251454 202807 251510 202816
rect 251638 202872 251694 202881
rect 251638 202807 251694 202816
rect 251652 193254 251680 202807
rect 251456 193248 251508 193254
rect 251456 193190 251508 193196
rect 251640 193248 251692 193254
rect 251640 193190 251692 193196
rect 251468 183569 251496 193190
rect 251454 183560 251510 183569
rect 251454 183495 251510 183504
rect 251638 183560 251694 183569
rect 251638 183495 251694 183504
rect 251652 173942 251680 183495
rect 251456 173936 251508 173942
rect 251456 173878 251508 173884
rect 251640 173936 251692 173942
rect 251640 173878 251692 173884
rect 251468 164218 251496 173878
rect 251456 164212 251508 164218
rect 251456 164154 251508 164160
rect 251640 164212 251692 164218
rect 251640 164154 251692 164160
rect 251652 154601 251680 164154
rect 251454 154592 251510 154601
rect 251454 154527 251510 154536
rect 251638 154592 251694 154601
rect 251638 154527 251694 154536
rect 251468 138122 251496 154527
rect 251376 138094 251496 138122
rect 251376 137986 251404 138094
rect 251376 137958 251496 137986
rect 251468 125594 251496 137958
rect 251456 125588 251508 125594
rect 251456 125530 251508 125536
rect 251456 116000 251508 116006
rect 251456 115942 251508 115948
rect 251468 106282 251496 115942
rect 251456 106276 251508 106282
rect 251456 106218 251508 106224
rect 251456 96688 251508 96694
rect 251456 96630 251508 96636
rect 251468 86970 251496 96630
rect 251456 86964 251508 86970
rect 251456 86906 251508 86912
rect 251456 77308 251508 77314
rect 251456 77250 251508 77256
rect 251468 48521 251496 77250
rect 251454 48512 251510 48521
rect 251454 48447 251510 48456
rect 251362 48376 251418 48385
rect 251362 48311 251418 48320
rect 251376 37346 251404 48311
rect 251376 37318 251496 37346
rect 251468 37262 251496 37318
rect 251456 37256 251508 37262
rect 251456 37198 251508 37204
rect 251362 27704 251418 27713
rect 251362 27639 251418 27648
rect 251376 27606 251404 27639
rect 251364 27600 251416 27606
rect 251364 27542 251416 27548
rect 251364 19304 251416 19310
rect 251364 19246 251416 19252
rect 251272 10328 251324 10334
rect 251272 10270 251324 10276
rect 251376 6186 251404 19246
rect 251364 6180 251416 6186
rect 251364 6122 251416 6128
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 250444 4140 250496 4146
rect 250444 4082 250496 4088
rect 251468 480 251496 5170
rect 251836 3398 251864 336670
rect 252664 10402 252692 340054
rect 253204 337544 253256 337550
rect 253204 337486 253256 337492
rect 252652 10396 252704 10402
rect 252652 10338 252704 10344
rect 252652 7948 252704 7954
rect 252652 7890 252704 7896
rect 251824 3392 251876 3398
rect 251824 3334 251876 3340
rect 252664 480 252692 7890
rect 253216 3330 253244 337486
rect 253492 337414 253520 340068
rect 253480 337408 253532 337414
rect 253480 337350 253532 337356
rect 253848 9240 253900 9246
rect 253848 9182 253900 9188
rect 253204 3324 253256 3330
rect 253204 3266 253256 3272
rect 253860 480 253888 9182
rect 253952 6254 253980 340068
rect 254044 340054 254518 340082
rect 254044 10470 254072 340054
rect 254964 338094 254992 340068
rect 255438 340054 255544 340082
rect 254952 338088 255004 338094
rect 254952 338030 255004 338036
rect 254584 337748 254636 337754
rect 254584 337690 254636 337696
rect 254032 10464 254084 10470
rect 254032 10406 254084 10412
rect 253940 6248 253992 6254
rect 253940 6190 253992 6196
rect 254596 3262 254624 337690
rect 255516 6322 255544 340054
rect 255608 340054 255990 340082
rect 255608 10538 255636 340054
rect 255964 337680 256016 337686
rect 255964 337622 256016 337628
rect 255596 10532 255648 10538
rect 255596 10474 255648 10480
rect 255504 6316 255556 6322
rect 255504 6258 255556 6264
rect 255044 3460 255096 3466
rect 255044 3402 255096 3408
rect 254584 3256 254636 3262
rect 254584 3198 254636 3204
rect 255056 480 255084 3402
rect 255976 3194 256004 337622
rect 256436 336734 256464 340068
rect 256804 340054 256910 340082
rect 256988 340054 257462 340082
rect 256424 336728 256476 336734
rect 256424 336670 256476 336676
rect 256240 8016 256292 8022
rect 256240 7958 256292 7964
rect 255964 3188 256016 3194
rect 255964 3130 256016 3136
rect 256252 480 256280 7958
rect 256804 6390 256832 340054
rect 256792 6384 256844 6390
rect 256792 6326 256844 6332
rect 256988 5302 257016 340054
rect 257344 337408 257396 337414
rect 257344 337350 257396 337356
rect 256976 5296 257028 5302
rect 256976 5238 257028 5244
rect 257356 3126 257384 337350
rect 257908 337210 257936 340068
rect 258276 340054 258382 340082
rect 258552 340054 258934 340082
rect 257896 337204 257948 337210
rect 257896 337146 257948 337152
rect 258172 334756 258224 334762
rect 258172 334698 258224 334704
rect 258184 13190 258212 334698
rect 258172 13184 258224 13190
rect 258172 13126 258224 13132
rect 258276 6458 258304 340054
rect 258552 334762 258580 340054
rect 258724 337952 258776 337958
rect 258724 337894 258776 337900
rect 258540 334756 258592 334762
rect 258540 334698 258592 334704
rect 258264 6452 258316 6458
rect 258264 6394 258316 6400
rect 257436 4004 257488 4010
rect 257436 3946 257488 3952
rect 257344 3120 257396 3126
rect 257344 3062 257396 3068
rect 257448 480 257476 3946
rect 258632 3528 258684 3534
rect 258632 3470 258684 3476
rect 258644 480 258672 3470
rect 258736 3058 258764 337894
rect 259380 337550 259408 340068
rect 259472 340054 259854 340082
rect 260116 340054 260406 340082
rect 259368 337544 259420 337550
rect 259368 337486 259420 337492
rect 258816 337476 258868 337482
rect 258816 337418 258868 337424
rect 258724 3052 258776 3058
rect 258724 2994 258776 3000
rect 258828 2990 258856 337418
rect 259366 17096 259422 17105
rect 259366 17031 259422 17040
rect 259380 16697 259408 17031
rect 259366 16688 259422 16697
rect 259366 16623 259422 16632
rect 259472 6526 259500 340054
rect 260116 337822 260144 340054
rect 259644 337816 259696 337822
rect 259644 337758 259696 337764
rect 260104 337816 260156 337822
rect 260104 337758 260156 337764
rect 259656 331226 259684 337758
rect 260104 337680 260156 337686
rect 260104 337622 260156 337628
rect 259644 331220 259696 331226
rect 259644 331162 259696 331168
rect 259828 331220 259880 331226
rect 259828 331162 259880 331168
rect 259840 328438 259868 331162
rect 259828 328432 259880 328438
rect 259828 328374 259880 328380
rect 259920 318844 259972 318850
rect 259920 318786 259972 318792
rect 259932 311914 259960 318786
rect 259736 311908 259788 311914
rect 259736 311850 259788 311856
rect 259920 311908 259972 311914
rect 259920 311850 259972 311856
rect 259748 309126 259776 311850
rect 259736 309120 259788 309126
rect 259736 309062 259788 309068
rect 259644 299600 259696 299606
rect 259644 299542 259696 299548
rect 259656 299470 259684 299542
rect 259644 299464 259696 299470
rect 259644 299406 259696 299412
rect 259828 299464 259880 299470
rect 259828 299406 259880 299412
rect 259840 289898 259868 299406
rect 259748 289870 259868 289898
rect 259748 289814 259776 289870
rect 259736 289808 259788 289814
rect 259736 289750 259788 289756
rect 259920 289808 259972 289814
rect 259920 289750 259972 289756
rect 259932 280265 259960 289750
rect 259550 280256 259606 280265
rect 259550 280191 259606 280200
rect 259918 280256 259974 280265
rect 259918 280191 259974 280200
rect 259564 280158 259592 280191
rect 259552 280152 259604 280158
rect 259552 280094 259604 280100
rect 259552 273080 259604 273086
rect 259552 273022 259604 273028
rect 259564 260846 259592 273022
rect 259552 260840 259604 260846
rect 259552 260782 259604 260788
rect 259552 253768 259604 253774
rect 259552 253710 259604 253716
rect 259564 251190 259592 253710
rect 259552 251184 259604 251190
rect 259552 251126 259604 251132
rect 259644 244180 259696 244186
rect 259644 244122 259696 244128
rect 259656 241398 259684 244122
rect 259644 241392 259696 241398
rect 259644 241334 259696 241340
rect 259828 241392 259880 241398
rect 259828 241334 259880 241340
rect 259840 222222 259868 241334
rect 259644 222216 259696 222222
rect 259644 222158 259696 222164
rect 259828 222216 259880 222222
rect 259828 222158 259880 222164
rect 259656 222086 259684 222158
rect 259644 222080 259696 222086
rect 259644 222022 259696 222028
rect 259828 222080 259880 222086
rect 259828 222022 259880 222028
rect 259840 215234 259868 222022
rect 259748 215206 259868 215234
rect 259748 205578 259776 215206
rect 259656 205550 259776 205578
rect 259656 202881 259684 205550
rect 259642 202872 259698 202881
rect 259642 202807 259698 202816
rect 259918 202872 259974 202881
rect 259918 202807 259974 202816
rect 259932 193254 259960 202807
rect 259736 193248 259788 193254
rect 259736 193190 259788 193196
rect 259920 193248 259972 193254
rect 259920 193190 259972 193196
rect 259748 186266 259776 193190
rect 259656 186238 259776 186266
rect 259656 179586 259684 186238
rect 259644 179580 259696 179586
rect 259644 179522 259696 179528
rect 259736 174004 259788 174010
rect 259736 173946 259788 173952
rect 259748 169114 259776 173946
rect 259736 169108 259788 169114
rect 259736 169050 259788 169056
rect 259920 169108 259972 169114
rect 259920 169050 259972 169056
rect 259932 164257 259960 169050
rect 259642 164248 259698 164257
rect 259918 164248 259974 164257
rect 259642 164183 259644 164192
rect 259696 164183 259698 164192
rect 259828 164212 259880 164218
rect 259644 164154 259696 164160
rect 259918 164183 259974 164192
rect 259828 164154 259880 164160
rect 259840 154222 259868 164154
rect 259828 154216 259880 154222
rect 259828 154158 259880 154164
rect 259644 142180 259696 142186
rect 259644 142122 259696 142128
rect 259656 142066 259684 142122
rect 259656 142050 259776 142066
rect 259656 142044 259788 142050
rect 259656 142038 259736 142044
rect 259736 141986 259788 141992
rect 259828 124228 259880 124234
rect 259828 124170 259880 124176
rect 259840 115462 259868 124170
rect 259828 115456 259880 115462
rect 259828 115398 259880 115404
rect 259828 115320 259880 115326
rect 259828 115262 259880 115268
rect 259840 106298 259868 115262
rect 259748 106282 259868 106298
rect 259736 106276 259880 106282
rect 259788 106270 259828 106276
rect 259736 106218 259788 106224
rect 259828 106218 259880 106224
rect 259840 99362 259868 106218
rect 259748 99334 259868 99362
rect 259748 91746 259776 99334
rect 259748 91718 259868 91746
rect 259840 86986 259868 91718
rect 259840 86958 259960 86986
rect 259932 77738 259960 86958
rect 259748 77710 259960 77738
rect 259748 62694 259776 77710
rect 259736 62688 259788 62694
rect 259736 62630 259788 62636
rect 259920 62620 259972 62626
rect 259920 62562 259972 62568
rect 259932 48226 259960 62562
rect 259748 48198 259960 48226
rect 259748 37262 259776 48198
rect 259736 37256 259788 37262
rect 259736 37198 259788 37204
rect 259736 27668 259788 27674
rect 259736 27610 259788 27616
rect 259748 22114 259776 27610
rect 259656 22086 259776 22114
rect 259656 14482 259684 22086
rect 259644 14476 259696 14482
rect 259644 14418 259696 14424
rect 259828 8084 259880 8090
rect 259828 8026 259880 8032
rect 259460 6520 259512 6526
rect 259460 6462 259512 6468
rect 258816 2984 258868 2990
rect 258816 2926 258868 2932
rect 259840 480 259868 8026
rect 260116 2922 260144 337622
rect 260852 337346 260880 340068
rect 261036 340054 261326 340082
rect 261496 340054 261878 340082
rect 260840 337340 260892 337346
rect 260840 337282 260892 337288
rect 260932 335640 260984 335646
rect 260932 335582 260984 335588
rect 260654 87136 260710 87145
rect 260654 87071 260656 87080
rect 260708 87071 260710 87080
rect 260656 87042 260708 87048
rect 260746 63744 260802 63753
rect 260746 63679 260802 63688
rect 260760 63617 260788 63679
rect 260746 63608 260802 63617
rect 260746 63543 260802 63552
rect 260944 14550 260972 335582
rect 260932 14544 260984 14550
rect 260932 14486 260984 14492
rect 261036 6594 261064 340054
rect 261392 337612 261444 337618
rect 261392 337554 261444 337560
rect 261404 334370 261432 337554
rect 261496 335646 261524 340054
rect 262324 337754 262352 340068
rect 262416 340054 262798 340082
rect 263060 340054 263350 340082
rect 262312 337748 262364 337754
rect 262312 337690 262364 337696
rect 261484 335640 261536 335646
rect 261484 335582 261536 335588
rect 261404 334342 261524 334370
rect 261024 6588 261076 6594
rect 261024 6530 261076 6536
rect 261024 4072 261076 4078
rect 261024 4014 261076 4020
rect 260104 2916 260156 2922
rect 260104 2858 260156 2864
rect 261036 480 261064 4014
rect 261496 2854 261524 334342
rect 262416 8158 262444 340054
rect 263060 336734 263088 340054
rect 263796 337278 263824 340068
rect 263888 340054 264270 340082
rect 264440 340054 264822 340082
rect 263784 337272 263836 337278
rect 263784 337214 263836 337220
rect 262864 336728 262916 336734
rect 262864 336670 262916 336676
rect 263048 336728 263100 336734
rect 263048 336670 263100 336676
rect 262876 327162 262904 336670
rect 263692 335640 263744 335646
rect 263692 335582 263744 335588
rect 262784 327134 262904 327162
rect 262784 322318 262812 327134
rect 262772 322312 262824 322318
rect 262772 322254 262824 322260
rect 262680 317484 262732 317490
rect 262680 317426 262732 317432
rect 262692 315994 262720 317426
rect 262680 315988 262732 315994
rect 262680 315930 262732 315936
rect 262680 306400 262732 306406
rect 262600 306348 262680 306354
rect 262600 306342 262732 306348
rect 262600 306326 262720 306342
rect 262600 299538 262628 306326
rect 262588 299532 262640 299538
rect 262588 299474 262640 299480
rect 262680 299464 262732 299470
rect 262680 299406 262732 299412
rect 262692 283642 262720 299406
rect 262600 283614 262720 283642
rect 262600 278746 262628 283614
rect 262508 278718 262628 278746
rect 262508 269142 262536 278718
rect 262496 269136 262548 269142
rect 262496 269078 262548 269084
rect 262588 269136 262640 269142
rect 262588 269078 262640 269084
rect 262600 260846 262628 269078
rect 262588 260840 262640 260846
rect 262588 260782 262640 260788
rect 262680 260772 262732 260778
rect 262680 260714 262732 260720
rect 262692 251954 262720 260714
rect 262508 251926 262720 251954
rect 262508 247081 262536 251926
rect 262494 247072 262550 247081
rect 262494 247007 262550 247016
rect 262770 246936 262826 246945
rect 262770 246871 262826 246880
rect 262784 235958 262812 246871
rect 262772 235952 262824 235958
rect 262772 235894 262824 235900
rect 262588 226364 262640 226370
rect 262588 226306 262640 226312
rect 262600 219502 262628 226306
rect 262588 219496 262640 219502
rect 262588 219438 262640 219444
rect 262680 219360 262732 219366
rect 262680 219302 262732 219308
rect 262692 202910 262720 219302
rect 262588 202904 262640 202910
rect 262588 202846 262640 202852
rect 262680 202904 262732 202910
rect 262680 202846 262732 202852
rect 262600 201482 262628 202846
rect 262588 201476 262640 201482
rect 262588 201418 262640 201424
rect 262772 201476 262824 201482
rect 262772 201418 262824 201424
rect 262784 191842 262812 201418
rect 262692 191814 262812 191842
rect 262692 186266 262720 191814
rect 262600 186238 262720 186266
rect 262600 173942 262628 186238
rect 262588 173936 262640 173942
rect 262588 173878 262640 173884
rect 262680 173936 262732 173942
rect 262680 173878 262732 173884
rect 262692 164354 262720 173878
rect 262680 164348 262732 164354
rect 262680 164290 262732 164296
rect 262588 164280 262640 164286
rect 262588 164222 262640 164228
rect 262600 157434 262628 164222
rect 262508 157406 262628 157434
rect 262508 153218 262536 157406
rect 262508 153190 262628 153218
rect 262600 144906 262628 153190
rect 262588 144900 262640 144906
rect 262588 144842 262640 144848
rect 262772 144900 262824 144906
rect 262772 144842 262824 144848
rect 262784 139992 262812 144842
rect 262692 139964 262812 139992
rect 262692 128466 262720 139964
rect 262692 128438 262812 128466
rect 262784 125633 262812 128438
rect 262586 125624 262642 125633
rect 262586 125559 262588 125568
rect 262640 125559 262642 125568
rect 262770 125624 262826 125633
rect 262770 125559 262772 125568
rect 262588 125530 262640 125536
rect 262824 125559 262826 125568
rect 262772 125530 262824 125536
rect 262784 118046 262812 125530
rect 262588 118040 262640 118046
rect 262588 117982 262640 117988
rect 262772 118040 262824 118046
rect 262772 117982 262824 117988
rect 262600 113234 262628 117982
rect 262600 113206 262720 113234
rect 262692 106298 262720 113206
rect 262692 106270 262812 106298
rect 262784 103714 262812 106270
rect 262600 103686 262812 103714
rect 262600 103494 262628 103686
rect 262588 103488 262640 103494
rect 262588 103430 262640 103436
rect 262772 103488 262824 103494
rect 262772 103430 262824 103436
rect 262784 102134 262812 103430
rect 262772 102128 262824 102134
rect 262772 102070 262824 102076
rect 262772 92540 262824 92546
rect 262772 92482 262824 92488
rect 262784 89010 262812 92482
rect 262772 89004 262824 89010
rect 262772 88946 262824 88952
rect 262680 75948 262732 75954
rect 262680 75890 262732 75896
rect 262692 67640 262720 75890
rect 262600 67612 262720 67640
rect 262600 62830 262628 67612
rect 263414 63744 263470 63753
rect 263598 63744 263654 63753
rect 263470 63702 263598 63730
rect 263414 63679 263470 63688
rect 263598 63679 263654 63688
rect 262588 62824 262640 62830
rect 262588 62766 262640 62772
rect 262772 62824 262824 62830
rect 262772 62766 262824 62772
rect 262784 47002 262812 62766
rect 262600 46974 262812 47002
rect 262600 46918 262628 46974
rect 262588 46912 262640 46918
rect 262588 46854 262640 46860
rect 262772 46912 262824 46918
rect 262772 46854 262824 46860
rect 262784 45558 262812 46854
rect 262772 45552 262824 45558
rect 262772 45494 262824 45500
rect 262772 35964 262824 35970
rect 262772 35906 262824 35912
rect 262784 32450 262812 35906
rect 262600 32422 262812 32450
rect 262600 28914 262628 32422
rect 262600 28886 262720 28914
rect 262692 27606 262720 28886
rect 262588 27600 262640 27606
rect 262588 27542 262640 27548
rect 262680 27600 262732 27606
rect 262680 27542 262732 27548
rect 262600 14618 262628 27542
rect 263704 14686 263732 335582
rect 263692 14680 263744 14686
rect 263692 14622 263744 14628
rect 262588 14612 262640 14618
rect 262588 14554 262640 14560
rect 263888 8226 263916 340054
rect 264440 335646 264468 340054
rect 265268 337074 265296 340068
rect 265452 340054 265742 340082
rect 265912 340054 266294 340082
rect 265256 337068 265308 337074
rect 265256 337010 265308 337016
rect 264428 335640 264480 335646
rect 264428 335582 264480 335588
rect 265072 335640 265124 335646
rect 265452 335594 265480 340054
rect 265912 335646 265940 340054
rect 266740 337414 266768 340068
rect 266924 340054 267214 340082
rect 267384 340054 267674 340082
rect 266728 337408 266780 337414
rect 266728 337350 266780 337356
rect 265072 335582 265124 335588
rect 264980 186992 265032 186998
rect 264980 186934 265032 186940
rect 264992 182209 265020 186934
rect 264978 182200 265034 182209
rect 264978 182135 265034 182144
rect 265084 14754 265112 335582
rect 265268 335566 265480 335594
rect 265900 335640 265952 335646
rect 265900 335582 265952 335588
rect 266452 335640 266504 335646
rect 266924 335594 266952 340054
rect 267384 335646 267412 340054
rect 268212 336938 268240 340068
rect 268396 340054 268686 340082
rect 269146 340054 269252 340082
rect 268200 336932 268252 336938
rect 268200 336874 268252 336880
rect 266452 335582 266504 335588
rect 265268 318918 265296 335566
rect 265256 318912 265308 318918
rect 265256 318854 265308 318860
rect 265256 317484 265308 317490
rect 265256 317426 265308 317432
rect 265268 309126 265296 317426
rect 265256 309120 265308 309126
rect 265256 309062 265308 309068
rect 265256 299532 265308 299538
rect 265256 299474 265308 299480
rect 265268 278934 265296 299474
rect 265256 278928 265308 278934
rect 265256 278870 265308 278876
rect 265348 278724 265400 278730
rect 265348 278666 265400 278672
rect 265360 255950 265388 278666
rect 265348 255944 265400 255950
rect 265348 255886 265400 255892
rect 265348 248260 265400 248266
rect 265348 248202 265400 248208
rect 265360 234734 265388 248202
rect 265164 234728 265216 234734
rect 265164 234670 265216 234676
rect 265348 234728 265400 234734
rect 265348 234670 265400 234676
rect 265176 229090 265204 234670
rect 265164 229084 265216 229090
rect 265164 229026 265216 229032
rect 265532 229084 265584 229090
rect 265532 229026 265584 229032
rect 265544 219473 265572 229026
rect 265346 219464 265402 219473
rect 265346 219399 265402 219408
rect 265530 219464 265586 219473
rect 265530 219399 265586 219408
rect 265360 211177 265388 219399
rect 265162 211168 265218 211177
rect 265162 211103 265218 211112
rect 265346 211168 265402 211177
rect 265346 211103 265402 211112
rect 265176 200122 265204 211103
rect 265164 200116 265216 200122
rect 265164 200058 265216 200064
rect 265164 195288 265216 195294
rect 265164 195230 265216 195236
rect 265176 186998 265204 195230
rect 265164 186992 265216 186998
rect 265164 186934 265216 186940
rect 265254 182200 265310 182209
rect 265254 182135 265310 182144
rect 265268 164354 265296 182135
rect 265256 164348 265308 164354
rect 265256 164290 265308 164296
rect 265164 164280 265216 164286
rect 265164 164222 265216 164228
rect 265176 157418 265204 164222
rect 265164 157412 265216 157418
rect 265164 157354 265216 157360
rect 265256 157276 265308 157282
rect 265256 157218 265308 157224
rect 265268 133890 265296 157218
rect 265256 133884 265308 133890
rect 265256 133826 265308 133832
rect 265256 124228 265308 124234
rect 265256 124170 265308 124176
rect 265268 113370 265296 124170
rect 265176 113342 265296 113370
rect 265176 113234 265204 113342
rect 265176 113206 265296 113234
rect 265268 113150 265296 113206
rect 265256 113144 265308 113150
rect 265256 113086 265308 113092
rect 265256 103556 265308 103562
rect 265256 103498 265308 103504
rect 265268 93906 265296 103498
rect 265164 93900 265216 93906
rect 265164 93842 265216 93848
rect 265256 93900 265308 93906
rect 265256 93842 265308 93848
rect 265176 89010 265204 93842
rect 265164 89004 265216 89010
rect 265164 88946 265216 88952
rect 265440 74588 265492 74594
rect 265440 74530 265492 74536
rect 265452 67538 265480 74530
rect 265360 67510 265480 67538
rect 265360 62694 265388 67510
rect 265348 62688 265400 62694
rect 265348 62630 265400 62636
rect 265164 57928 265216 57934
rect 265164 57870 265216 57876
rect 265176 53174 265204 57870
rect 265164 53168 265216 53174
rect 265164 53110 265216 53116
rect 265348 53168 265400 53174
rect 265348 53110 265400 53116
rect 265360 42106 265388 53110
rect 265268 42078 265388 42106
rect 265268 27606 265296 42078
rect 265256 27600 265308 27606
rect 265256 27542 265308 27548
rect 265164 18012 265216 18018
rect 265164 17954 265216 17960
rect 265072 14748 265124 14754
rect 265072 14690 265124 14696
rect 265176 8294 265204 17954
rect 266464 14822 266492 335582
rect 266740 335566 266952 335594
rect 267372 335640 267424 335646
rect 268396 335594 268424 340054
rect 269028 337408 269080 337414
rect 269028 337350 269080 337356
rect 267372 335582 267424 335588
rect 267844 335566 268424 335594
rect 266740 321638 266768 335566
rect 267844 321638 267872 335566
rect 266728 321632 266780 321638
rect 266728 321574 266780 321580
rect 267832 321632 267884 321638
rect 267832 321574 267884 321580
rect 266636 318844 266688 318850
rect 266636 318786 266688 318792
rect 267740 318844 267792 318850
rect 267740 318786 267792 318792
rect 266648 309262 266676 318786
rect 267752 310978 267780 318786
rect 267752 310950 267872 310978
rect 266636 309256 266688 309262
rect 266636 309198 266688 309204
rect 266636 309120 266688 309126
rect 266636 309062 266688 309068
rect 266648 298178 266676 309062
rect 267844 299606 267872 310950
rect 267832 299600 267884 299606
rect 267832 299542 267884 299548
rect 267740 299464 267792 299470
rect 267740 299406 267792 299412
rect 266636 298172 266688 298178
rect 266636 298114 266688 298120
rect 266636 296744 266688 296750
rect 266636 296686 266688 296692
rect 266648 287094 266676 296686
rect 267752 288454 267780 299406
rect 267740 288448 267792 288454
rect 267740 288390 267792 288396
rect 267832 288448 267884 288454
rect 267832 288390 267884 288396
rect 266636 287088 266688 287094
rect 266636 287030 266688 287036
rect 266728 287088 266780 287094
rect 266728 287030 266780 287036
rect 266740 285666 266768 287030
rect 266728 285660 266780 285666
rect 266728 285602 266780 285608
rect 267844 283642 267872 288390
rect 267752 283614 267872 283642
rect 267752 278769 267780 283614
rect 267738 278760 267794 278769
rect 267738 278695 267794 278704
rect 267830 278624 267886 278633
rect 267830 278559 267886 278568
rect 266728 276072 266780 276078
rect 266648 276020 266728 276026
rect 266648 276014 266780 276020
rect 266648 275998 266768 276014
rect 266648 274650 266676 275998
rect 266636 274644 266688 274650
rect 266636 274586 266688 274592
rect 267844 265690 267872 278559
rect 267752 265662 267872 265690
rect 267752 260846 267780 265662
rect 266636 260840 266688 260846
rect 266636 260782 266688 260788
rect 267740 260840 267792 260846
rect 267740 260782 267792 260788
rect 266648 256714 266676 260782
rect 267832 260772 267884 260778
rect 267832 260714 267884 260720
rect 267844 258058 267872 260714
rect 267832 258052 267884 258058
rect 267832 257994 267884 258000
rect 268016 257984 268068 257990
rect 268016 257926 268068 257932
rect 266648 256686 266768 256714
rect 266740 251190 266768 256686
rect 266728 251184 266780 251190
rect 266728 251126 266780 251132
rect 266820 251184 266872 251190
rect 266820 251126 266872 251132
rect 266832 241534 266860 251126
rect 268028 248441 268056 257926
rect 267738 248432 267794 248441
rect 267738 248367 267794 248376
rect 268014 248432 268070 248441
rect 268014 248367 268070 248376
rect 266728 241528 266780 241534
rect 266728 241470 266780 241476
rect 266820 241528 266872 241534
rect 266820 241470 266872 241476
rect 266740 234818 266768 241470
rect 267752 240106 267780 248367
rect 267740 240100 267792 240106
rect 267740 240042 267792 240048
rect 267924 240100 267976 240106
rect 267924 240042 267976 240048
rect 266740 234790 266860 234818
rect 266832 231826 266860 234790
rect 266740 231798 266860 231826
rect 266740 220674 266768 231798
rect 266740 220646 266860 220674
rect 266832 211177 266860 220646
rect 266634 211168 266690 211177
rect 266634 211103 266690 211112
rect 266818 211168 266874 211177
rect 266818 211103 266874 211112
rect 266648 202910 266676 211103
rect 267936 209817 267964 240042
rect 267738 209808 267794 209817
rect 267738 209743 267794 209752
rect 267922 209808 267978 209817
rect 267922 209743 267978 209752
rect 266636 202904 266688 202910
rect 266636 202846 266688 202852
rect 266728 202904 266780 202910
rect 266728 202846 266780 202852
rect 266740 194834 266768 202846
rect 267752 201414 267780 209743
rect 267740 201408 267792 201414
rect 267740 201350 267792 201356
rect 267924 201408 267976 201414
rect 267924 201350 267976 201356
rect 266648 194806 266768 194834
rect 266648 191826 266676 194806
rect 266636 191820 266688 191826
rect 266636 191762 266688 191768
rect 266636 186312 266688 186318
rect 266636 186254 266688 186260
rect 266648 182186 266676 186254
rect 267936 182209 267964 201350
rect 267738 182200 267794 182209
rect 266648 182158 266768 182186
rect 266740 178786 266768 182158
rect 267738 182135 267794 182144
rect 267922 182200 267978 182209
rect 267922 182135 267978 182144
rect 266740 178758 266860 178786
rect 266832 173942 266860 178758
rect 267752 173942 267780 182135
rect 266636 173936 266688 173942
rect 266634 173904 266636 173913
rect 266820 173936 266872 173942
rect 266688 173904 266690 173913
rect 266634 173839 266690 173848
rect 266818 173904 266820 173913
rect 267740 173936 267792 173942
rect 266872 173904 266874 173913
rect 267740 173878 267792 173884
rect 267832 173936 267884 173942
rect 267832 173878 267884 173884
rect 266818 173839 266874 173848
rect 266832 166818 266860 173839
rect 266740 166790 266860 166818
rect 266740 144974 266768 166790
rect 267844 164354 267872 173878
rect 267832 164348 267884 164354
rect 267832 164290 267884 164296
rect 267740 164280 267792 164286
rect 267740 164222 267792 164228
rect 267752 157486 267780 164222
rect 267740 157480 267792 157486
rect 267740 157422 267792 157428
rect 267740 157344 267792 157350
rect 267740 157286 267792 157292
rect 266728 144968 266780 144974
rect 266728 144910 266780 144916
rect 267752 144906 267780 157286
rect 267740 144900 267792 144906
rect 267740 144842 267792 144848
rect 267924 144900 267976 144906
rect 267924 144842 267976 144848
rect 266728 144832 266780 144838
rect 266728 144774 266780 144780
rect 266740 135425 266768 144774
rect 267936 139992 267964 144842
rect 267844 139964 267964 139992
rect 266726 135416 266782 135425
rect 266726 135351 266782 135360
rect 266634 135280 266690 135289
rect 266634 135215 266636 135224
rect 266688 135215 266690 135224
rect 266728 135244 266780 135250
rect 266636 135186 266688 135192
rect 266728 135186 266780 135192
rect 266740 116113 266768 135186
rect 267844 128466 267872 139964
rect 267844 128438 267964 128466
rect 267936 125633 267964 128438
rect 267738 125624 267794 125633
rect 267738 125559 267740 125568
rect 267792 125559 267794 125568
rect 267922 125624 267978 125633
rect 267922 125559 267924 125568
rect 267740 125530 267792 125536
rect 267976 125559 267978 125568
rect 267924 125530 267976 125536
rect 267936 120680 267964 125530
rect 267844 120652 267964 120680
rect 266726 116104 266782 116113
rect 266726 116039 266782 116048
rect 266634 115968 266690 115977
rect 266634 115903 266690 115912
rect 266648 106298 266676 115903
rect 267844 111092 267872 120652
rect 267752 111064 267872 111092
rect 266648 106282 266768 106298
rect 266648 106276 266780 106282
rect 266648 106270 266728 106276
rect 266728 106218 266780 106224
rect 266820 106276 266872 106282
rect 267752 106264 267780 111064
rect 267832 106276 267884 106282
rect 267752 106236 267832 106264
rect 266820 106218 266872 106224
rect 267832 106218 267884 106224
rect 267924 106276 267976 106282
rect 267924 106218 267976 106224
rect 266832 103494 266860 106218
rect 267936 103494 267964 106218
rect 266820 103488 266872 103494
rect 266820 103430 266872 103436
rect 267924 103488 267976 103494
rect 267924 103430 267976 103436
rect 266820 96484 266872 96490
rect 266820 96426 266872 96432
rect 266832 58002 266860 96426
rect 267740 93900 267792 93906
rect 267740 93842 267792 93848
rect 267752 85542 267780 93842
rect 267740 85536 267792 85542
rect 267740 85478 267792 85484
rect 267832 85536 267884 85542
rect 267832 85478 267884 85484
rect 267844 66298 267872 85478
rect 267740 66292 267792 66298
rect 267740 66234 267792 66240
rect 267832 66292 267884 66298
rect 267832 66234 267884 66240
rect 267752 58002 267780 66234
rect 266728 57996 266780 58002
rect 266728 57938 266780 57944
rect 266820 57996 266872 58002
rect 266820 57938 266872 57944
rect 267740 57996 267792 58002
rect 267740 57938 267792 57944
rect 267832 57996 267884 58002
rect 267832 57938 267884 57944
rect 266740 46986 266768 57938
rect 267844 48346 267872 57938
rect 267832 48340 267884 48346
rect 267832 48282 267884 48288
rect 267924 48204 267976 48210
rect 267924 48146 267976 48152
rect 266544 46980 266596 46986
rect 266544 46922 266596 46928
rect 266728 46980 266780 46986
rect 266728 46922 266780 46928
rect 266556 37330 266584 46922
rect 266544 37324 266596 37330
rect 266544 37266 266596 37272
rect 266636 37324 266688 37330
rect 266636 37266 266688 37272
rect 266648 17898 266676 37266
rect 267936 37262 267964 48146
rect 267924 37256 267976 37262
rect 267924 37198 267976 37204
rect 267832 28620 267884 28626
rect 267832 28562 267884 28568
rect 267844 22114 267872 28562
rect 267844 22086 267964 22114
rect 267936 21978 267964 22086
rect 266556 17870 266676 17898
rect 267752 21950 267964 21978
rect 266452 14816 266504 14822
rect 266452 14758 266504 14764
rect 266556 10606 266584 17870
rect 267752 10674 267780 21950
rect 267740 10668 267792 10674
rect 267740 10610 267792 10616
rect 266544 10600 266596 10606
rect 266544 10542 266596 10548
rect 265164 8288 265216 8294
rect 265164 8230 265216 8236
rect 263876 8220 263928 8226
rect 263876 8162 263928 8168
rect 267004 8220 267056 8226
rect 267004 8162 267056 8168
rect 262404 8152 262456 8158
rect 262404 8094 262456 8100
rect 263416 8152 263468 8158
rect 263416 8094 263468 8100
rect 262220 3664 262272 3670
rect 262220 3606 262272 3612
rect 261484 2848 261536 2854
rect 261484 2790 261536 2796
rect 262232 480 262260 3606
rect 263428 480 263456 8094
rect 264612 3936 264664 3942
rect 264612 3878 264664 3884
rect 264624 480 264652 3878
rect 265808 3596 265860 3602
rect 265808 3538 265860 3544
rect 265820 480 265848 3538
rect 267016 480 267044 8162
rect 269040 4146 269068 337350
rect 269224 14890 269252 340054
rect 269684 337482 269712 340068
rect 269868 340054 270158 340082
rect 269672 337476 269724 337482
rect 269672 337418 269724 337424
rect 269868 335594 269896 340054
rect 269316 335566 269896 335594
rect 269212 14884 269264 14890
rect 269212 14826 269264 14832
rect 269316 10742 269344 335566
rect 270498 325680 270554 325689
rect 270498 325615 270554 325624
rect 270512 316062 270540 325615
rect 270500 316056 270552 316062
rect 270500 315998 270552 316004
rect 270500 202156 270552 202162
rect 270500 202098 270552 202104
rect 270512 195838 270540 202098
rect 270500 195832 270552 195838
rect 270500 195774 270552 195780
rect 270500 130416 270552 130422
rect 270500 130358 270552 130364
rect 270512 125633 270540 130358
rect 270498 125624 270554 125633
rect 270498 125559 270554 125568
rect 270604 18018 270632 340068
rect 271156 337142 271184 340068
rect 271248 340054 271630 340082
rect 271984 340054 272090 340082
rect 271144 337136 271196 337142
rect 271144 337078 271196 337084
rect 271248 334354 271276 340054
rect 271788 337476 271840 337482
rect 271788 337418 271840 337424
rect 271328 337272 271380 337278
rect 271328 337214 271380 337220
rect 270776 334348 270828 334354
rect 270776 334290 270828 334296
rect 271236 334348 271288 334354
rect 271236 334290 271288 334296
rect 270788 325689 270816 334290
rect 271340 334234 271368 337214
rect 271156 334206 271368 334234
rect 270774 325680 270830 325689
rect 270774 325615 270830 325624
rect 270684 316056 270736 316062
rect 270684 315998 270736 316004
rect 270696 314673 270724 315998
rect 270682 314664 270738 314673
rect 270682 314599 270738 314608
rect 270866 314664 270922 314673
rect 270866 314599 270922 314608
rect 270880 304994 270908 314599
rect 270880 304966 271000 304994
rect 270972 296750 271000 304966
rect 270776 296744 270828 296750
rect 270776 296686 270828 296692
rect 270960 296744 271012 296750
rect 270960 296686 271012 296692
rect 270788 295322 270816 296686
rect 270776 295316 270828 295322
rect 270776 295258 270828 295264
rect 270960 295316 271012 295322
rect 270960 295258 271012 295264
rect 270972 282266 271000 295258
rect 270776 282260 270828 282266
rect 270776 282202 270828 282208
rect 270960 282260 271012 282266
rect 270960 282202 271012 282208
rect 270788 273306 270816 282202
rect 270696 273278 270816 273306
rect 270696 263634 270724 273278
rect 270684 263628 270736 263634
rect 270684 263570 270736 263576
rect 270684 263492 270736 263498
rect 270684 263434 270736 263440
rect 270696 260846 270724 263434
rect 270684 260840 270736 260846
rect 270684 260782 270736 260788
rect 270684 240236 270736 240242
rect 270684 240178 270736 240184
rect 270696 238746 270724 240178
rect 270684 238740 270736 238746
rect 270684 238682 270736 238688
rect 270684 233844 270736 233850
rect 270684 233786 270736 233792
rect 270696 220833 270724 233786
rect 270682 220824 270738 220833
rect 270682 220759 270738 220768
rect 270958 220824 271014 220833
rect 270958 220759 271014 220768
rect 270972 219434 271000 220759
rect 270776 219428 270828 219434
rect 270776 219370 270828 219376
rect 270960 219428 271012 219434
rect 270960 219370 271012 219376
rect 270788 209817 270816 219370
rect 270774 209808 270830 209817
rect 270774 209743 270830 209752
rect 270958 209808 271014 209817
rect 270958 209743 271014 209752
rect 270972 202162 271000 209743
rect 270960 202156 271012 202162
rect 270960 202098 271012 202104
rect 270684 195832 270736 195838
rect 270684 195774 270736 195780
rect 270696 191826 270724 195774
rect 270684 191820 270736 191826
rect 270684 191762 270736 191768
rect 270868 191820 270920 191826
rect 270868 191762 270920 191768
rect 270880 190466 270908 191762
rect 270868 190460 270920 190466
rect 270868 190402 270920 190408
rect 271052 190460 271104 190466
rect 271052 190402 271104 190408
rect 271064 180849 271092 190402
rect 270774 180840 270830 180849
rect 270774 180775 270830 180784
rect 271050 180840 271106 180849
rect 271050 180775 271106 180784
rect 270788 172582 270816 180775
rect 270776 172576 270828 172582
rect 270776 172518 270828 172524
rect 270868 172440 270920 172446
rect 270868 172382 270920 172388
rect 270880 167142 270908 172382
rect 270868 167136 270920 167142
rect 270868 167078 270920 167084
rect 270684 167000 270736 167006
rect 270684 166942 270736 166948
rect 270696 144906 270724 166942
rect 270684 144900 270736 144906
rect 270684 144842 270736 144848
rect 270684 140004 270736 140010
rect 270684 139946 270736 139952
rect 270696 130422 270724 139946
rect 270684 130416 270736 130422
rect 270684 130358 270736 130364
rect 270682 125624 270738 125633
rect 270682 125559 270684 125568
rect 270736 125559 270738 125568
rect 270684 125530 270736 125536
rect 270684 120692 270736 120698
rect 270684 120634 270736 120640
rect 270696 111110 270724 120634
rect 270684 111104 270736 111110
rect 270684 111046 270736 111052
rect 270868 111104 270920 111110
rect 270868 111046 270920 111052
rect 270880 106321 270908 111046
rect 270682 106312 270738 106321
rect 270682 106247 270684 106256
rect 270736 106247 270738 106256
rect 270866 106312 270922 106321
rect 270866 106247 270922 106256
rect 270684 106218 270736 106224
rect 270684 101380 270736 101386
rect 270684 101322 270736 101328
rect 270696 96626 270724 101322
rect 270684 96620 270736 96626
rect 270684 96562 270736 96568
rect 270868 96620 270920 96626
rect 270868 96562 270920 96568
rect 270880 86986 270908 96562
rect 270788 86958 270908 86986
rect 270788 80782 270816 86958
rect 270776 80776 270828 80782
rect 270776 80718 270828 80724
rect 270776 67652 270828 67658
rect 270776 67594 270828 67600
rect 270788 66230 270816 67594
rect 270776 66224 270828 66230
rect 270776 66166 270828 66172
rect 270776 56636 270828 56642
rect 270776 56578 270828 56584
rect 270788 53122 270816 56578
rect 270788 53094 270908 53122
rect 270880 38690 270908 53094
rect 270776 38684 270828 38690
rect 270776 38626 270828 38632
rect 270868 38684 270920 38690
rect 270868 38626 270920 38632
rect 270788 22166 270816 38626
rect 270776 22160 270828 22166
rect 270776 22102 270828 22108
rect 270592 18012 270644 18018
rect 270592 17954 270644 17960
rect 270500 17944 270552 17950
rect 270500 17886 270552 17892
rect 270512 10810 270540 17886
rect 270592 17876 270644 17882
rect 270592 17818 270644 17824
rect 270604 14958 270632 17818
rect 270592 14952 270644 14958
rect 270592 14894 270644 14900
rect 270500 10804 270552 10810
rect 270500 10746 270552 10752
rect 269304 10736 269356 10742
rect 269304 10678 269356 10684
rect 270500 8288 270552 8294
rect 270500 8230 270552 8236
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 269028 4140 269080 4146
rect 269028 4082 269080 4088
rect 268120 480 268148 4082
rect 269304 3256 269356 3262
rect 269304 3198 269356 3204
rect 269316 480 269344 3198
rect 270512 480 270540 8230
rect 271156 4418 271184 334206
rect 271144 4412 271196 4418
rect 271144 4354 271196 4360
rect 271800 626 271828 337418
rect 271880 243092 271932 243098
rect 271880 243034 271932 243040
rect 271892 229129 271920 243034
rect 271878 229120 271934 229129
rect 271878 229055 271934 229064
rect 271880 26172 271932 26178
rect 271880 26114 271932 26120
rect 271892 10878 271920 26114
rect 271984 18018 272012 340054
rect 272628 337958 272656 340068
rect 272720 340054 273102 340082
rect 273364 340054 273562 340082
rect 272616 337952 272668 337958
rect 272616 337894 272668 337900
rect 272720 334354 272748 340054
rect 272800 337340 272852 337346
rect 272800 337282 272852 337288
rect 272248 334348 272300 334354
rect 272248 334290 272300 334296
rect 272708 334348 272760 334354
rect 272708 334290 272760 334296
rect 272260 324358 272288 334290
rect 272812 334234 272840 337282
rect 272536 334206 272840 334234
rect 272156 324352 272208 324358
rect 272156 324294 272208 324300
rect 272248 324352 272300 324358
rect 272248 324294 272300 324300
rect 272168 314634 272196 324294
rect 272156 314628 272208 314634
rect 272156 314570 272208 314576
rect 272248 296744 272300 296750
rect 272248 296686 272300 296692
rect 272260 295322 272288 296686
rect 272248 295316 272300 295322
rect 272248 295258 272300 295264
rect 272156 285728 272208 285734
rect 272156 285670 272208 285676
rect 272168 282282 272196 285670
rect 272168 282254 272288 282282
rect 272260 269113 272288 282254
rect 272062 269104 272118 269113
rect 272062 269039 272118 269048
rect 272246 269104 272302 269113
rect 272246 269039 272302 269048
rect 272076 259486 272104 269039
rect 272064 259480 272116 259486
rect 272156 259480 272208 259486
rect 272064 259422 272116 259428
rect 272154 259448 272156 259457
rect 272208 259448 272210 259457
rect 272154 259383 272210 259392
rect 272430 259448 272486 259457
rect 272430 259383 272486 259392
rect 272444 258058 272472 259383
rect 272432 258052 272484 258058
rect 272432 257994 272484 258000
rect 272432 249756 272484 249762
rect 272432 249698 272484 249704
rect 272444 243098 272472 249698
rect 272432 243092 272484 243098
rect 272432 243034 272484 243040
rect 272062 229120 272118 229129
rect 272062 229055 272064 229064
rect 272116 229055 272118 229064
rect 272064 229026 272116 229032
rect 272156 220788 272208 220794
rect 272156 220730 272208 220736
rect 272168 214690 272196 220730
rect 272168 214662 272288 214690
rect 272260 214418 272288 214662
rect 272168 214390 272288 214418
rect 272168 202881 272196 214390
rect 272154 202872 272210 202881
rect 272154 202807 272210 202816
rect 272338 202736 272394 202745
rect 272338 202671 272394 202680
rect 272352 201482 272380 202671
rect 272340 201476 272392 201482
rect 272340 201418 272392 201424
rect 272340 193180 272392 193186
rect 272340 193122 272392 193128
rect 272352 191842 272380 193122
rect 272352 191814 272472 191842
rect 272444 186318 272472 191814
rect 272156 186312 272208 186318
rect 272156 186254 272208 186260
rect 272432 186312 272484 186318
rect 272432 186254 272484 186260
rect 272168 183569 272196 186254
rect 272154 183560 272210 183569
rect 272154 183495 272210 183504
rect 272338 183424 272394 183433
rect 272338 183359 272394 183368
rect 272352 172582 272380 183359
rect 272248 172576 272300 172582
rect 272248 172518 272300 172524
rect 272340 172576 272392 172582
rect 272340 172518 272392 172524
rect 272260 167686 272288 172518
rect 272064 167680 272116 167686
rect 272064 167622 272116 167628
rect 272248 167680 272300 167686
rect 272248 167622 272300 167628
rect 272076 162874 272104 167622
rect 272076 162846 272196 162874
rect 272168 158030 272196 162846
rect 272156 158024 272208 158030
rect 272156 157966 272208 157972
rect 272156 148980 272208 148986
rect 272156 148922 272208 148928
rect 272168 144906 272196 148922
rect 272156 144900 272208 144906
rect 272156 144842 272208 144848
rect 272432 144900 272484 144906
rect 272432 144842 272484 144848
rect 272444 143546 272472 144842
rect 272432 143540 272484 143546
rect 272432 143482 272484 143488
rect 272432 135244 272484 135250
rect 272432 135186 272484 135192
rect 272444 125866 272472 135186
rect 272156 125860 272208 125866
rect 272156 125802 272208 125808
rect 272432 125860 272484 125866
rect 272432 125802 272484 125808
rect 272168 125594 272196 125802
rect 272156 125588 272208 125594
rect 272156 125530 272208 125536
rect 272432 125588 272484 125594
rect 272432 125530 272484 125536
rect 272444 124166 272472 125530
rect 272432 124160 272484 124166
rect 272432 124102 272484 124108
rect 272432 114572 272484 114578
rect 272432 114514 272484 114520
rect 272444 106554 272472 114514
rect 272156 106548 272208 106554
rect 272156 106490 272208 106496
rect 272432 106548 272484 106554
rect 272432 106490 272484 106496
rect 272168 106282 272196 106490
rect 272156 106276 272208 106282
rect 272156 106218 272208 106224
rect 272432 106276 272484 106282
rect 272432 106218 272484 106224
rect 272444 90386 272472 106218
rect 272352 90358 272472 90386
rect 272352 84182 272380 90358
rect 272340 84176 272392 84182
rect 272340 84118 272392 84124
rect 272248 74588 272300 74594
rect 272248 74530 272300 74536
rect 272260 67726 272288 74530
rect 272248 67720 272300 67726
rect 272248 67662 272300 67668
rect 272248 67108 272300 67114
rect 272248 67050 272300 67056
rect 272260 57916 272288 67050
rect 272168 57888 272288 57916
rect 272168 38690 272196 57888
rect 272156 38684 272208 38690
rect 272156 38626 272208 38632
rect 272248 38684 272300 38690
rect 272248 38626 272300 38632
rect 272260 37262 272288 38626
rect 272248 37256 272300 37262
rect 272248 37198 272300 37204
rect 272340 37256 272392 37262
rect 272340 37198 272392 37204
rect 272352 35902 272380 37198
rect 272340 35896 272392 35902
rect 272340 35838 272392 35844
rect 272248 26308 272300 26314
rect 272248 26250 272300 26256
rect 272260 26178 272288 26250
rect 272248 26172 272300 26178
rect 272248 26114 272300 26120
rect 271972 18012 272024 18018
rect 271972 17954 272024 17960
rect 271972 17876 272024 17882
rect 271972 17818 272024 17824
rect 271984 15026 272012 17818
rect 271972 15020 272024 15026
rect 271972 14962 272024 14968
rect 271880 10872 271932 10878
rect 271880 10814 271932 10820
rect 272536 4350 272564 334206
rect 273074 63744 273130 63753
rect 273258 63744 273314 63753
rect 273130 63702 273258 63730
rect 273074 63679 273130 63688
rect 273258 63679 273314 63688
rect 273074 40216 273130 40225
rect 273258 40216 273314 40225
rect 273130 40174 273258 40202
rect 273074 40151 273130 40160
rect 273258 40151 273314 40160
rect 273364 15094 273392 340054
rect 274100 337006 274128 340068
rect 274284 340054 274574 340082
rect 274744 340054 275034 340082
rect 274088 337000 274140 337006
rect 274088 336942 274140 336948
rect 274284 331242 274312 340054
rect 273640 331214 274312 331242
rect 273548 316062 273576 316093
rect 273640 316062 273668 331214
rect 273536 316056 273588 316062
rect 273456 316004 273536 316010
rect 273456 315998 273588 316004
rect 273628 316056 273680 316062
rect 273628 315998 273680 316004
rect 273456 315982 273576 315998
rect 273456 309330 273484 315982
rect 273444 309324 273496 309330
rect 273444 309266 273496 309272
rect 273536 301572 273588 301578
rect 273536 301514 273588 301520
rect 273548 293162 273576 301514
rect 273548 293134 273668 293162
rect 273640 282826 273668 293134
rect 273548 282798 273668 282826
rect 273548 280158 273576 282798
rect 273536 280152 273588 280158
rect 273536 280094 273588 280100
rect 273628 280152 273680 280158
rect 273628 280094 273680 280100
rect 273640 263514 273668 280094
rect 273548 263486 273668 263514
rect 273548 260846 273576 263486
rect 273536 260840 273588 260846
rect 273536 260782 273588 260788
rect 273628 260840 273680 260846
rect 273628 260782 273680 260788
rect 273640 244202 273668 260782
rect 273548 244174 273668 244202
rect 273548 234682 273576 244174
rect 273456 234654 273576 234682
rect 273456 234598 273484 234654
rect 273444 234592 273496 234598
rect 273444 234534 273496 234540
rect 273628 234592 273680 234598
rect 273628 234534 273680 234540
rect 273640 220862 273668 234534
rect 273536 220856 273588 220862
rect 273536 220798 273588 220804
rect 273628 220856 273680 220862
rect 273628 220798 273680 220804
rect 273548 215370 273576 220798
rect 273456 215342 273576 215370
rect 273456 215286 273484 215342
rect 273444 215280 273496 215286
rect 273444 215222 273496 215228
rect 273628 215280 273680 215286
rect 273628 215222 273680 215228
rect 273640 207754 273668 215222
rect 273548 207726 273668 207754
rect 273548 202842 273576 207726
rect 273536 202836 273588 202842
rect 273536 202778 273588 202784
rect 273628 202836 273680 202842
rect 273628 202778 273680 202784
rect 273640 186266 273668 202778
rect 273548 186238 273668 186266
rect 273548 183530 273576 186238
rect 273536 183524 273588 183530
rect 273536 183466 273588 183472
rect 273628 183524 273680 183530
rect 273628 183466 273680 183472
rect 273640 157434 273668 183466
rect 273456 157406 273668 157434
rect 273456 157298 273484 157406
rect 273456 157270 273576 157298
rect 273548 137850 273576 157270
rect 273548 137822 273668 137850
rect 273640 128330 273668 137822
rect 273548 128302 273668 128330
rect 273548 118726 273576 128302
rect 273536 118720 273588 118726
rect 273536 118662 273588 118668
rect 273628 118652 273680 118658
rect 273628 118594 273680 118600
rect 273640 109018 273668 118594
rect 273548 108990 273668 109018
rect 273548 95334 273576 108990
rect 273536 95328 273588 95334
rect 273536 95270 273588 95276
rect 273628 95328 273680 95334
rect 273628 95270 273680 95276
rect 273640 85542 273668 95270
rect 273536 85536 273588 85542
rect 273536 85478 273588 85484
rect 273628 85536 273680 85542
rect 273628 85478 273680 85484
rect 273548 67538 273576 85478
rect 273456 67510 273576 67538
rect 273456 66230 273484 67510
rect 273444 66224 273496 66230
rect 273444 66166 273496 66172
rect 273536 50992 273588 50998
rect 273536 50934 273588 50940
rect 273548 48278 273576 50934
rect 273536 48272 273588 48278
rect 273536 48214 273588 48220
rect 273536 38684 273588 38690
rect 273536 38626 273588 38632
rect 273548 22114 273576 38626
rect 273456 22086 273576 22114
rect 273456 17950 273484 22086
rect 273444 17944 273496 17950
rect 273444 17886 273496 17892
rect 274744 15162 274772 340054
rect 275572 337550 275600 340068
rect 275560 337544 275612 337550
rect 275560 337486 275612 337492
rect 275928 337544 275980 337550
rect 275928 337486 275980 337492
rect 274732 15156 274784 15162
rect 274732 15098 274784 15104
rect 273352 15088 273404 15094
rect 273352 15030 273404 15036
rect 274088 6180 274140 6186
rect 274088 6122 274140 6128
rect 272524 4344 272576 4350
rect 272524 4286 272576 4292
rect 272892 3188 272944 3194
rect 272892 3130 272944 3136
rect 271708 598 271828 626
rect 271708 480 271736 598
rect 272904 480 272932 3130
rect 274100 480 274128 6122
rect 275940 3942 275968 337486
rect 276032 11014 276060 340068
rect 276124 340054 276506 340082
rect 276124 14414 276152 340054
rect 277044 337686 277072 340068
rect 277518 340054 277624 340082
rect 277032 337680 277084 337686
rect 277032 337622 277084 337628
rect 276112 14408 276164 14414
rect 276112 14350 276164 14356
rect 276020 11008 276072 11014
rect 276020 10950 276072 10956
rect 277596 10266 277624 340054
rect 277688 340054 277978 340082
rect 277688 14346 277716 340054
rect 278516 336870 278544 340068
rect 278792 340054 278990 340082
rect 279068 340054 279450 340082
rect 278504 336864 278556 336870
rect 278504 336806 278556 336812
rect 278792 333334 278820 340054
rect 278780 333328 278832 333334
rect 278780 333270 278832 333276
rect 278964 333328 279016 333334
rect 278964 333270 279016 333276
rect 278872 328500 278924 328506
rect 278872 328442 278924 328448
rect 278884 157434 278912 328442
rect 278792 157406 278912 157434
rect 278792 157298 278820 157406
rect 278792 157270 278912 157298
rect 278884 80186 278912 157270
rect 278792 80158 278912 80186
rect 278792 41290 278820 80158
rect 278792 41262 278912 41290
rect 278778 29336 278834 29345
rect 278778 29271 278780 29280
rect 278832 29271 278834 29280
rect 278780 29242 278832 29248
rect 278780 16584 278832 16590
rect 278778 16552 278780 16561
rect 278832 16552 278834 16561
rect 278778 16487 278834 16496
rect 277676 14340 277728 14346
rect 277676 14282 277728 14288
rect 278884 14278 278912 41262
rect 278872 14272 278924 14278
rect 278872 14214 278924 14220
rect 277584 10260 277636 10266
rect 277584 10202 277636 10208
rect 278976 10198 279004 333270
rect 279068 328506 279096 340054
rect 279988 337618 280016 340068
rect 280356 340054 280462 340082
rect 280632 340054 280922 340082
rect 281184 340054 281474 340082
rect 281644 340054 281934 340082
rect 282104 340054 282394 340082
rect 282946 340054 283144 340082
rect 279976 337612 280028 337618
rect 279976 337554 280028 337560
rect 280252 335640 280304 335646
rect 280252 335582 280304 335588
rect 279056 328500 279108 328506
rect 279056 328442 279108 328448
rect 280264 14210 280292 335582
rect 280252 14204 280304 14210
rect 280252 14146 280304 14152
rect 278964 10192 279016 10198
rect 278964 10134 279016 10140
rect 280356 10130 280384 340054
rect 280632 335646 280660 340054
rect 281184 336802 281212 340054
rect 281448 337612 281500 337618
rect 281448 337554 281500 337560
rect 281172 336796 281224 336802
rect 281172 336738 281224 336744
rect 280620 335640 280672 335646
rect 280620 335582 280672 335588
rect 281264 29300 281316 29306
rect 281264 29242 281316 29248
rect 281276 29209 281304 29242
rect 281262 29200 281318 29209
rect 281262 29135 281318 29144
rect 280344 10124 280396 10130
rect 280344 10066 280396 10072
rect 280068 6248 280120 6254
rect 280068 6190 280120 6196
rect 275284 3936 275336 3942
rect 275284 3878 275336 3884
rect 275928 3936 275980 3942
rect 275928 3878 275980 3884
rect 275296 480 275324 3878
rect 278872 3800 278924 3806
rect 278872 3742 278924 3748
rect 276480 3256 276532 3262
rect 276480 3198 276532 3204
rect 276492 480 276520 3198
rect 277676 3188 277728 3194
rect 277676 3130 277728 3136
rect 277688 480 277716 3130
rect 278884 480 278912 3742
rect 280080 480 280108 6190
rect 281460 610 281488 337554
rect 281540 335640 281592 335646
rect 281540 335582 281592 335588
rect 281552 11898 281580 335582
rect 281540 11892 281592 11898
rect 281540 11834 281592 11840
rect 281644 11830 281672 340054
rect 282104 335646 282132 340054
rect 282092 335640 282144 335646
rect 282092 335582 282144 335588
rect 283012 335640 283064 335646
rect 283012 335582 283064 335588
rect 282734 40216 282790 40225
rect 282918 40216 282974 40225
rect 282790 40174 282918 40202
rect 282734 40151 282790 40160
rect 282918 40151 282974 40160
rect 281632 11824 281684 11830
rect 281632 11766 281684 11772
rect 283024 6662 283052 335582
rect 283116 7585 283144 340054
rect 283208 340054 283406 340082
rect 283576 340054 283866 340082
rect 283102 7576 283158 7585
rect 283102 7511 283158 7520
rect 283012 6656 283064 6662
rect 283012 6598 283064 6604
rect 283208 5370 283236 340054
rect 283576 335646 283604 340054
rect 284404 336734 284432 340068
rect 284588 340054 284878 340082
rect 285140 340054 285338 340082
rect 285798 340054 285904 340082
rect 284392 336728 284444 336734
rect 284392 336670 284444 336676
rect 283564 335640 283616 335646
rect 283564 335582 283616 335588
rect 284484 335232 284536 335238
rect 284484 335174 284536 335180
rect 284300 329588 284352 329594
rect 284300 329530 284352 329536
rect 284312 5438 284340 329530
rect 284496 8945 284524 335174
rect 284588 329594 284616 340054
rect 285140 332586 285168 340054
rect 285588 337680 285640 337686
rect 285588 337622 285640 337628
rect 284668 332580 284720 332586
rect 284668 332522 284720 332528
rect 285128 332580 285180 332586
rect 285128 332522 285180 332528
rect 284576 329588 284628 329594
rect 284576 329530 284628 329536
rect 284680 318850 284708 332522
rect 284668 318844 284720 318850
rect 284668 318786 284720 318792
rect 284760 318844 284812 318850
rect 284760 318786 284812 318792
rect 284772 316010 284800 318786
rect 284680 315982 284800 316010
rect 284680 311914 284708 315982
rect 284668 311908 284720 311914
rect 284668 311850 284720 311856
rect 284576 306400 284628 306406
rect 284576 306342 284628 306348
rect 284588 289814 284616 306342
rect 284576 289808 284628 289814
rect 284576 289750 284628 289756
rect 284760 289740 284812 289746
rect 284760 289682 284812 289688
rect 284772 280158 284800 289682
rect 284576 280152 284628 280158
rect 284576 280094 284628 280100
rect 284760 280152 284812 280158
rect 284760 280094 284812 280100
rect 284588 278769 284616 280094
rect 284574 278760 284630 278769
rect 284574 278695 284630 278704
rect 284758 278760 284814 278769
rect 284758 278695 284814 278704
rect 284772 269142 284800 278695
rect 284576 269136 284628 269142
rect 284576 269078 284628 269084
rect 284760 269136 284812 269142
rect 284760 269078 284812 269084
rect 284588 260914 284616 269078
rect 284576 260908 284628 260914
rect 284576 260850 284628 260856
rect 284760 260908 284812 260914
rect 284760 260850 284812 260856
rect 284772 249898 284800 260850
rect 284668 249892 284720 249898
rect 284668 249834 284720 249840
rect 284760 249892 284812 249898
rect 284760 249834 284812 249840
rect 284680 249762 284708 249834
rect 284668 249756 284720 249762
rect 284668 249698 284720 249704
rect 284852 240168 284904 240174
rect 284852 240110 284904 240116
rect 284864 225078 284892 240110
rect 284852 225072 284904 225078
rect 284852 225014 284904 225020
rect 284852 224936 284904 224942
rect 284852 224878 284904 224884
rect 284864 220833 284892 224878
rect 284666 220824 284722 220833
rect 284666 220759 284722 220768
rect 284850 220824 284906 220833
rect 284850 220759 284906 220768
rect 284680 212498 284708 220759
rect 284668 212492 284720 212498
rect 284668 212434 284720 212440
rect 284852 212492 284904 212498
rect 284852 212434 284904 212440
rect 284864 211154 284892 212434
rect 284864 211138 284984 211154
rect 284668 211132 284720 211138
rect 284864 211132 284996 211138
rect 284864 211126 284944 211132
rect 284668 211074 284720 211080
rect 284944 211074 284996 211080
rect 284680 201521 284708 211074
rect 284956 211043 284984 211074
rect 284666 201512 284722 201521
rect 284666 201447 284722 201456
rect 284850 201512 284906 201521
rect 284850 201447 284906 201456
rect 284864 193225 284892 201447
rect 284666 193216 284722 193225
rect 284666 193151 284722 193160
rect 284850 193216 284906 193225
rect 284850 193151 284906 193160
rect 284680 183666 284708 193151
rect 284668 183660 284720 183666
rect 284668 183602 284720 183608
rect 284668 183524 284720 183530
rect 284668 183466 284720 183472
rect 284680 180810 284708 183466
rect 284668 180804 284720 180810
rect 284668 180746 284720 180752
rect 284760 171148 284812 171154
rect 284760 171090 284812 171096
rect 284772 132546 284800 171090
rect 285494 157992 285550 158001
rect 285494 157927 285550 157936
rect 285508 157457 285536 157927
rect 285494 157448 285550 157457
rect 285494 157383 285550 157392
rect 284680 132518 284800 132546
rect 284680 128382 284708 132518
rect 284668 128376 284720 128382
rect 284668 128318 284720 128324
rect 284760 128308 284812 128314
rect 284760 128250 284812 128256
rect 284772 122806 284800 128250
rect 284760 122800 284812 122806
rect 284760 122742 284812 122748
rect 284760 122664 284812 122670
rect 284760 122606 284812 122612
rect 284772 117994 284800 122606
rect 284680 117966 284800 117994
rect 284680 113150 284708 117966
rect 284668 113144 284720 113150
rect 284668 113086 284720 113092
rect 284668 103556 284720 103562
rect 284668 103498 284720 103504
rect 284680 95198 284708 103498
rect 284668 95192 284720 95198
rect 284668 95134 284720 95140
rect 284760 95124 284812 95130
rect 284760 95066 284812 95072
rect 284772 84182 284800 95066
rect 284760 84176 284812 84182
rect 284760 84118 284812 84124
rect 284668 66292 284720 66298
rect 284668 66234 284720 66240
rect 284680 58002 284708 66234
rect 284668 57996 284720 58002
rect 284668 57938 284720 57944
rect 284760 57996 284812 58002
rect 284760 57938 284812 57944
rect 284772 48346 284800 57938
rect 284668 48340 284720 48346
rect 284668 48282 284720 48288
rect 284760 48340 284812 48346
rect 284760 48282 284812 48288
rect 284680 44742 284708 48282
rect 284668 44736 284720 44742
rect 284668 44678 284720 44684
rect 284760 29028 284812 29034
rect 284760 28970 284812 28976
rect 284772 27606 284800 28970
rect 284760 27600 284812 27606
rect 284760 27542 284812 27548
rect 284760 18012 284812 18018
rect 284760 17954 284812 17960
rect 284772 11898 284800 17954
rect 284576 11892 284628 11898
rect 284576 11834 284628 11840
rect 284760 11892 284812 11898
rect 284760 11834 284812 11840
rect 284482 8936 284538 8945
rect 284482 8871 284538 8880
rect 284588 7546 284616 11834
rect 284576 7540 284628 7546
rect 284576 7482 284628 7488
rect 284300 5432 284352 5438
rect 284300 5374 284352 5380
rect 283196 5364 283248 5370
rect 283196 5306 283248 5312
rect 283656 5296 283708 5302
rect 283656 5238 283708 5244
rect 282460 3936 282512 3942
rect 282460 3878 282512 3884
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281448 604 281500 610
rect 281448 546 281500 552
rect 281276 480 281304 546
rect 282472 480 282500 3878
rect 283668 480 283696 5238
rect 285600 3330 285628 337622
rect 285680 335640 285732 335646
rect 285680 335582 285732 335588
rect 285692 5506 285720 335582
rect 285772 306468 285824 306474
rect 285772 306410 285824 306416
rect 285784 296750 285812 306410
rect 285772 296744 285824 296750
rect 285772 296686 285824 296692
rect 285772 291916 285824 291922
rect 285772 291858 285824 291864
rect 285784 278798 285812 291858
rect 285772 278792 285824 278798
rect 285772 278734 285824 278740
rect 285770 202872 285826 202881
rect 285770 202807 285826 202816
rect 285784 198082 285812 202807
rect 285772 198076 285824 198082
rect 285772 198018 285824 198024
rect 285876 9314 285904 340054
rect 285968 340054 286350 340082
rect 286612 340054 286810 340082
rect 287164 340054 287270 340082
rect 287348 340054 287822 340082
rect 287992 340054 288282 340082
rect 288544 340054 288742 340082
rect 289004 340054 289294 340082
rect 289464 340054 289754 340082
rect 289832 340054 290214 340082
rect 285968 335646 285996 340054
rect 286612 335646 286640 340054
rect 285956 335640 286008 335646
rect 285956 335582 286008 335588
rect 286048 335640 286100 335646
rect 286048 335582 286100 335588
rect 286600 335640 286652 335646
rect 286600 335582 286652 335588
rect 287060 335640 287112 335646
rect 287060 335582 287112 335588
rect 286060 318866 286088 335582
rect 285968 318838 286088 318866
rect 285968 311914 285996 318838
rect 285956 311908 286008 311914
rect 285956 311850 286008 311856
rect 286048 296744 286100 296750
rect 286048 296686 286100 296692
rect 286060 291922 286088 296686
rect 286048 291916 286100 291922
rect 286048 291858 286100 291864
rect 286048 278792 286100 278798
rect 286048 278734 286100 278740
rect 286060 261089 286088 278734
rect 286046 261080 286102 261089
rect 286046 261015 286102 261024
rect 285954 260944 286010 260953
rect 285954 260879 286010 260888
rect 285968 249830 285996 260879
rect 285956 249824 286008 249830
rect 286048 249824 286100 249830
rect 285956 249766 286008 249772
rect 286046 249792 286048 249801
rect 286100 249792 286102 249801
rect 286046 249727 286102 249736
rect 285954 249656 286010 249665
rect 285954 249591 286010 249600
rect 285968 245002 285996 249591
rect 285956 244996 286008 245002
rect 285956 244938 286008 244944
rect 285956 234524 286008 234530
rect 285956 234466 286008 234472
rect 285968 222193 285996 234466
rect 285954 222184 286010 222193
rect 285954 222119 286010 222128
rect 286138 222184 286194 222193
rect 286138 222119 286194 222128
rect 286152 220833 286180 222119
rect 285954 220824 286010 220833
rect 285954 220759 286010 220768
rect 286138 220824 286194 220833
rect 286138 220759 286194 220768
rect 285968 211834 285996 220759
rect 285968 211806 286180 211834
rect 286152 202910 286180 211806
rect 285956 202904 286008 202910
rect 285954 202872 285956 202881
rect 286140 202904 286192 202910
rect 286008 202872 286010 202881
rect 286140 202846 286192 202852
rect 285954 202807 286010 202816
rect 285956 198076 286008 198082
rect 285956 198018 286008 198024
rect 285968 183734 285996 198018
rect 285956 183728 286008 183734
rect 285956 183670 286008 183676
rect 285956 183592 286008 183598
rect 285956 183534 286008 183540
rect 285968 172689 285996 183534
rect 285954 172680 286010 172689
rect 285954 172615 286010 172624
rect 286046 172544 286102 172553
rect 286046 172479 286102 172488
rect 286060 171086 286088 172479
rect 286048 171080 286100 171086
rect 286048 171022 286100 171028
rect 285956 161492 286008 161498
rect 285956 161434 286008 161440
rect 285968 158710 285996 161434
rect 285956 158704 286008 158710
rect 285956 158646 286008 158652
rect 286048 140820 286100 140826
rect 286048 140762 286100 140768
rect 286060 140706 286088 140762
rect 285968 140678 286088 140706
rect 285968 122777 285996 140678
rect 285954 122768 286010 122777
rect 285954 122703 286010 122712
rect 286230 122768 286286 122777
rect 286230 122703 286286 122712
rect 286244 113218 286272 122703
rect 286048 113212 286100 113218
rect 286048 113154 286100 113160
rect 286232 113212 286284 113218
rect 286232 113154 286284 113160
rect 286060 113082 286088 113154
rect 286048 113076 286100 113082
rect 286048 113018 286100 113024
rect 286232 113076 286284 113082
rect 286232 113018 286284 113024
rect 286244 85678 286272 113018
rect 286232 85672 286284 85678
rect 286232 85614 286284 85620
rect 285956 85604 286008 85610
rect 285956 85546 286008 85552
rect 285968 84182 285996 85546
rect 285956 84176 286008 84182
rect 285956 84118 286008 84124
rect 285956 66292 286008 66298
rect 285956 66234 286008 66240
rect 285968 58002 285996 66234
rect 285956 57996 286008 58002
rect 285956 57938 286008 57944
rect 286048 57996 286100 58002
rect 286048 57938 286100 57944
rect 286060 48414 286088 57938
rect 286048 48408 286100 48414
rect 286048 48350 286100 48356
rect 285956 48340 286008 48346
rect 285956 48282 286008 48288
rect 285968 38865 285996 48282
rect 285954 38856 286010 38865
rect 285954 38791 286010 38800
rect 285954 38584 286010 38593
rect 285954 38519 286010 38528
rect 285968 29034 285996 38519
rect 285956 29028 286008 29034
rect 285956 28970 286008 28976
rect 286048 29028 286100 29034
rect 286048 28970 286100 28976
rect 286060 27606 286088 28970
rect 286048 27600 286100 27606
rect 286048 27542 286100 27548
rect 285956 18012 286008 18018
rect 285956 17954 286008 17960
rect 285864 9308 285916 9314
rect 285864 9250 285916 9256
rect 285968 7478 285996 17954
rect 285956 7472 286008 7478
rect 285956 7414 286008 7420
rect 287072 7410 287100 335582
rect 287164 9382 287192 340054
rect 287348 11966 287376 340054
rect 287992 335646 288020 340054
rect 288256 337816 288308 337822
rect 288256 337758 288308 337764
rect 287980 335640 288032 335646
rect 287980 335582 288032 335588
rect 287336 11960 287388 11966
rect 287336 11902 287388 11908
rect 287152 9376 287204 9382
rect 287152 9318 287204 9324
rect 287060 7404 287112 7410
rect 287060 7346 287112 7352
rect 285680 5500 285732 5506
rect 285680 5442 285732 5448
rect 287152 5364 287204 5370
rect 287152 5306 287204 5312
rect 285956 3800 286008 3806
rect 285956 3742 286008 3748
rect 284760 3324 284812 3330
rect 284760 3266 284812 3272
rect 285588 3324 285640 3330
rect 285588 3266 285640 3272
rect 284772 480 284800 3266
rect 285968 480 285996 3742
rect 287164 480 287192 5306
rect 288268 626 288296 337758
rect 288440 335640 288492 335646
rect 288440 335582 288492 335588
rect 288452 7342 288480 335582
rect 288544 10062 288572 340054
rect 289004 336734 289032 340054
rect 288992 336728 289044 336734
rect 288992 336670 289044 336676
rect 289464 335646 289492 340054
rect 289452 335640 289504 335646
rect 289452 335582 289504 335588
rect 288808 319116 288860 319122
rect 288808 319058 288860 319064
rect 288820 311982 288848 319058
rect 288808 311976 288860 311982
rect 288808 311918 288860 311924
rect 288716 290012 288768 290018
rect 288716 289954 288768 289960
rect 288728 289814 288756 289954
rect 288716 289808 288768 289814
rect 288716 289750 288768 289756
rect 288808 289808 288860 289814
rect 288808 289750 288860 289756
rect 288820 278798 288848 289750
rect 288716 278792 288768 278798
rect 288716 278734 288768 278740
rect 288808 278792 288860 278798
rect 288808 278734 288860 278740
rect 288728 267782 288756 278734
rect 288716 267776 288768 267782
rect 288716 267718 288768 267724
rect 288808 267776 288860 267782
rect 288808 267718 288860 267724
rect 288820 258233 288848 267718
rect 288806 258224 288862 258233
rect 288806 258159 288862 258168
rect 288806 258088 288862 258097
rect 288806 258023 288862 258032
rect 288820 253994 288848 258023
rect 288820 253966 288940 253994
rect 288912 245614 288940 253966
rect 288900 245608 288952 245614
rect 288900 245550 288952 245556
rect 288992 236020 289044 236026
rect 288992 235962 289044 235968
rect 289004 224210 289032 235962
rect 288820 224182 289032 224210
rect 288820 218906 288848 224182
rect 288820 218878 289032 218906
rect 289004 201521 289032 218878
rect 288806 201512 288862 201521
rect 288806 201447 288862 201456
rect 288990 201512 289046 201521
rect 288990 201447 289046 201456
rect 288820 191826 288848 201447
rect 288808 191820 288860 191826
rect 288808 191762 288860 191768
rect 288808 179444 288860 179450
rect 288808 179386 288860 179392
rect 288820 176662 288848 179386
rect 288808 176656 288860 176662
rect 288808 176598 288860 176604
rect 288808 167068 288860 167074
rect 288808 167010 288860 167016
rect 288820 158658 288848 167010
rect 288820 158630 288940 158658
rect 288912 153898 288940 158630
rect 288820 153870 288940 153898
rect 288820 140758 288848 153870
rect 288808 140752 288860 140758
rect 288808 140694 288860 140700
rect 288624 131164 288676 131170
rect 288624 131106 288676 131112
rect 288636 121514 288664 131106
rect 288624 121508 288676 121514
rect 288624 121450 288676 121456
rect 288900 121508 288952 121514
rect 288900 121450 288952 121456
rect 288912 103562 288940 121450
rect 288808 103556 288860 103562
rect 288808 103498 288860 103504
rect 288900 103556 288952 103562
rect 288900 103498 288952 103504
rect 288820 100042 288848 103498
rect 288820 100014 288940 100042
rect 288912 89026 288940 100014
rect 288728 88998 288940 89026
rect 288728 82822 288756 88998
rect 288716 82816 288768 82822
rect 288716 82758 288768 82764
rect 288900 64932 288952 64938
rect 288900 64874 288952 64880
rect 288912 64841 288940 64874
rect 288714 64832 288770 64841
rect 288714 64767 288770 64776
rect 288898 64832 288954 64841
rect 288898 64767 288954 64776
rect 288728 55350 288756 64767
rect 288716 55344 288768 55350
rect 288716 55286 288768 55292
rect 288900 55276 288952 55282
rect 288900 55218 288952 55224
rect 288912 46986 288940 55218
rect 288716 46980 288768 46986
rect 288716 46922 288768 46928
rect 288900 46980 288952 46986
rect 288900 46922 288952 46928
rect 288728 37262 288756 46922
rect 288716 37256 288768 37262
rect 288716 37198 288768 37204
rect 288808 37188 288860 37194
rect 288808 37130 288860 37136
rect 288820 22250 288848 37130
rect 288636 22222 288848 22250
rect 288636 19258 288664 22222
rect 288636 19230 288848 19258
rect 288820 12034 288848 19230
rect 288808 12028 288860 12034
rect 288808 11970 288860 11976
rect 288532 10056 288584 10062
rect 288532 9998 288584 10004
rect 289832 9994 289860 340054
rect 290292 331242 290320 340190
rect 290464 337884 290516 337890
rect 290464 337826 290516 337832
rect 290108 331214 290320 331242
rect 290108 309194 290136 331214
rect 290004 309188 290056 309194
rect 290004 309130 290056 309136
rect 290096 309188 290148 309194
rect 290096 309130 290148 309136
rect 290016 302954 290044 309130
rect 290016 302926 290228 302954
rect 290200 294642 290228 302926
rect 290004 294636 290056 294642
rect 290004 294578 290056 294584
rect 290188 294636 290240 294642
rect 290188 294578 290240 294584
rect 290016 289814 290044 294578
rect 290004 289808 290056 289814
rect 290004 289750 290056 289756
rect 290188 289808 290240 289814
rect 290188 289750 290240 289756
rect 290200 269142 290228 289750
rect 290096 269136 290148 269142
rect 290096 269078 290148 269084
rect 290188 269136 290240 269142
rect 290188 269078 290240 269084
rect 290108 251258 290136 269078
rect 290004 251252 290056 251258
rect 290004 251194 290056 251200
rect 290096 251252 290148 251258
rect 290096 251194 290148 251200
rect 290016 247042 290044 251194
rect 290004 247036 290056 247042
rect 290004 246978 290056 246984
rect 290372 247036 290424 247042
rect 290372 246978 290424 246984
rect 290384 219609 290412 246978
rect 290370 219600 290426 219609
rect 290370 219535 290426 219544
rect 290094 219464 290150 219473
rect 290094 219399 290150 219408
rect 290108 218006 290136 219399
rect 290096 218000 290148 218006
rect 290096 217942 290148 217948
rect 290096 208412 290148 208418
rect 290096 208354 290148 208360
rect 290108 201550 290136 208354
rect 290096 201544 290148 201550
rect 290096 201486 290148 201492
rect 290188 201408 290240 201414
rect 290188 201350 290240 201356
rect 290200 193322 290228 201350
rect 290188 193316 290240 193322
rect 290188 193258 290240 193264
rect 290096 193180 290148 193186
rect 290096 193122 290148 193128
rect 290108 188698 290136 193122
rect 290096 188692 290148 188698
rect 290096 188634 290148 188640
rect 290004 179444 290056 179450
rect 290004 179386 290056 179392
rect 290016 153202 290044 179386
rect 290004 153196 290056 153202
rect 290004 153138 290056 153144
rect 290096 153196 290148 153202
rect 290096 153138 290148 153144
rect 290108 138106 290136 153138
rect 290096 138100 290148 138106
rect 290096 138042 290148 138048
rect 289912 132456 289964 132462
rect 289912 132398 289964 132404
rect 289924 104922 289952 132398
rect 289912 104916 289964 104922
rect 289912 104858 289964 104864
rect 290004 104916 290056 104922
rect 290004 104858 290056 104864
rect 290016 103494 290044 104858
rect 290004 103488 290056 103494
rect 290004 103430 290056 103436
rect 290096 103420 290148 103426
rect 290096 103362 290148 103368
rect 290108 75954 290136 103362
rect 289912 75948 289964 75954
rect 289912 75890 289964 75896
rect 290096 75948 290148 75954
rect 290096 75890 290148 75896
rect 289924 75834 289952 75890
rect 289924 75806 290044 75834
rect 290016 12102 290044 75806
rect 290004 12096 290056 12102
rect 290004 12038 290056 12044
rect 289820 9988 289872 9994
rect 289820 9930 289872 9936
rect 288440 7336 288492 7342
rect 288440 7278 288492 7284
rect 289820 6520 289872 6526
rect 289820 6462 289872 6468
rect 288440 6452 288492 6458
rect 288440 6394 288492 6400
rect 288452 3262 288480 6394
rect 288532 6384 288584 6390
rect 288532 6326 288584 6332
rect 288440 3256 288492 3262
rect 288440 3198 288492 3204
rect 288544 3194 288572 6326
rect 289544 3868 289596 3874
rect 289544 3810 289596 3816
rect 288532 3188 288584 3194
rect 288532 3130 288584 3136
rect 288268 598 288388 626
rect 288360 480 288388 598
rect 289556 480 289584 3810
rect 289832 3398 289860 6462
rect 289820 3392 289872 3398
rect 289820 3334 289872 3340
rect 290476 3126 290504 337826
rect 290554 16688 290610 16697
rect 290554 16623 290610 16632
rect 290568 16590 290596 16623
rect 290556 16584 290608 16590
rect 290556 16526 290608 16532
rect 291212 7274 291240 340068
rect 291304 340054 291686 340082
rect 291304 9926 291332 340054
rect 291764 335594 291792 340190
rect 291580 335566 291792 335594
rect 292592 340054 292698 340082
rect 292868 340054 293158 340082
rect 293328 340054 293710 340082
rect 293972 340054 294170 340082
rect 294248 340054 294630 340082
rect 291580 319410 291608 335566
rect 291488 319382 291608 319410
rect 291488 319138 291516 319382
rect 291488 319110 291608 319138
rect 291580 311250 291608 319110
rect 291488 311222 291608 311250
rect 291488 306377 291516 311222
rect 291474 306368 291530 306377
rect 291474 306303 291530 306312
rect 291750 306368 291806 306377
rect 291750 306303 291806 306312
rect 291764 287094 291792 306303
rect 291568 287088 291620 287094
rect 291568 287030 291620 287036
rect 291752 287088 291804 287094
rect 291752 287030 291804 287036
rect 291580 277506 291608 287030
rect 291568 277500 291620 277506
rect 291568 277442 291620 277448
rect 291568 277364 291620 277370
rect 291568 277306 291620 277312
rect 291580 276026 291608 277306
rect 291580 275998 291700 276026
rect 291672 267782 291700 275998
rect 291568 267776 291620 267782
rect 291568 267718 291620 267724
rect 291660 267776 291712 267782
rect 291660 267718 291712 267724
rect 291580 240106 291608 267718
rect 291568 240100 291620 240106
rect 291568 240042 291620 240048
rect 291844 240100 291896 240106
rect 291844 240042 291896 240048
rect 291856 236314 291884 240042
rect 291856 236286 292068 236314
rect 292040 219473 292068 236286
rect 291658 219464 291714 219473
rect 291658 219399 291714 219408
rect 292026 219464 292082 219473
rect 292026 219399 292082 219408
rect 291672 214606 291700 219399
rect 291660 214600 291712 214606
rect 291660 214542 291712 214548
rect 291660 204060 291712 204066
rect 291660 204002 291712 204008
rect 291672 193202 291700 204002
rect 291580 193174 291700 193202
rect 291580 191826 291608 193174
rect 291568 191820 291620 191826
rect 291568 191762 291620 191768
rect 291660 191820 291712 191826
rect 291660 191762 291712 191768
rect 291672 164257 291700 191762
rect 291474 164248 291530 164257
rect 291474 164183 291530 164192
rect 291658 164248 291714 164257
rect 291658 164183 291714 164192
rect 291488 153202 291516 164183
rect 291476 153196 291528 153202
rect 291476 153138 291528 153144
rect 291568 153196 291620 153202
rect 291568 153138 291620 153144
rect 291580 133906 291608 153138
rect 291488 133878 291608 133906
rect 291488 131102 291516 133878
rect 291476 131096 291528 131102
rect 291476 131038 291528 131044
rect 291568 122732 291620 122738
rect 291568 122674 291620 122680
rect 291580 113150 291608 122674
rect 291568 113144 291620 113150
rect 291568 113086 291620 113092
rect 291660 103624 291712 103630
rect 291660 103566 291712 103572
rect 291672 102134 291700 103566
rect 291660 102128 291712 102134
rect 291660 102070 291712 102076
rect 291660 92540 291712 92546
rect 291660 92482 291712 92488
rect 291672 85610 291700 92482
rect 291660 85604 291712 85610
rect 291660 85546 291712 85552
rect 291568 84244 291620 84250
rect 291568 84186 291620 84192
rect 291580 75954 291608 84186
rect 291384 75948 291436 75954
rect 291384 75890 291436 75896
rect 291568 75948 291620 75954
rect 291568 75890 291620 75896
rect 291396 75834 291424 75890
rect 291396 75806 291516 75834
rect 291488 58070 291516 75806
rect 291476 58064 291528 58070
rect 291476 58006 291528 58012
rect 291384 57928 291436 57934
rect 291384 57870 291436 57876
rect 291396 47054 291424 57870
rect 291384 47048 291436 47054
rect 291384 46990 291436 46996
rect 291476 46980 291528 46986
rect 291476 46922 291528 46928
rect 291488 28966 291516 46922
rect 291476 28960 291528 28966
rect 291476 28902 291528 28908
rect 291660 28960 291712 28966
rect 291660 28902 291712 28908
rect 291672 27554 291700 28902
rect 291580 27526 291700 27554
rect 291580 19990 291608 27526
rect 291568 19984 291620 19990
rect 291568 19926 291620 19932
rect 291568 19848 291620 19854
rect 291568 19790 291620 19796
rect 291580 12170 291608 19790
rect 291568 12164 291620 12170
rect 291568 12106 291620 12112
rect 291292 9920 291344 9926
rect 291292 9862 291344 9868
rect 291200 7268 291252 7274
rect 291200 7210 291252 7216
rect 292592 7206 292620 340054
rect 292764 335640 292816 335646
rect 292764 335582 292816 335588
rect 292776 13258 292804 335582
rect 292764 13252 292816 13258
rect 292764 13194 292816 13200
rect 292868 9858 292896 340054
rect 293328 335646 293356 340054
rect 293316 335640 293368 335646
rect 293316 335582 293368 335588
rect 292856 9852 292908 9858
rect 292856 9794 292908 9800
rect 292580 7200 292632 7206
rect 292580 7142 292632 7148
rect 293972 7138 294000 340054
rect 294248 335696 294276 340054
rect 294064 335668 294276 335696
rect 294064 9790 294092 335668
rect 294708 331242 294736 340190
rect 294248 331214 294736 331242
rect 295352 340054 295642 340082
rect 295720 340054 296102 340082
rect 296272 340054 296654 340082
rect 296732 340054 297114 340082
rect 297284 340054 297574 340082
rect 298126 340054 298232 340082
rect 294248 316062 294276 331214
rect 294144 316056 294196 316062
rect 294144 315998 294196 316004
rect 294236 316056 294288 316062
rect 294236 315998 294288 316004
rect 294156 296750 294184 315998
rect 294144 296744 294196 296750
rect 294144 296686 294196 296692
rect 294328 296744 294380 296750
rect 294328 296686 294380 296692
rect 294340 287094 294368 296686
rect 294236 287088 294288 287094
rect 294236 287030 294288 287036
rect 294328 287088 294380 287094
rect 294328 287030 294380 287036
rect 294248 278798 294276 287030
rect 294236 278792 294288 278798
rect 294236 278734 294288 278740
rect 294328 278792 294380 278798
rect 294328 278734 294380 278740
rect 294340 264994 294368 278734
rect 294236 264988 294288 264994
rect 294236 264930 294288 264936
rect 294328 264988 294380 264994
rect 294328 264930 294380 264936
rect 294248 247042 294276 264930
rect 294236 247036 294288 247042
rect 294236 246978 294288 246984
rect 294420 246900 294472 246906
rect 294420 246842 294472 246848
rect 294432 222222 294460 246842
rect 294328 222216 294380 222222
rect 294328 222158 294380 222164
rect 294420 222216 294472 222222
rect 294420 222158 294472 222164
rect 294340 202910 294368 222158
rect 294236 202904 294288 202910
rect 294236 202846 294288 202852
rect 294328 202904 294380 202910
rect 294328 202846 294380 202852
rect 294248 198082 294276 202846
rect 294236 198076 294288 198082
rect 294236 198018 294288 198024
rect 294420 198076 294472 198082
rect 294420 198018 294472 198024
rect 294432 184278 294460 198018
rect 294420 184272 294472 184278
rect 294420 184214 294472 184220
rect 294328 179444 294380 179450
rect 294328 179386 294380 179392
rect 294340 178022 294368 179386
rect 294328 178016 294380 178022
rect 294328 177958 294380 177964
rect 294328 168428 294380 168434
rect 294328 168370 294380 168376
rect 294340 158710 294368 168370
rect 294328 158704 294380 158710
rect 294328 158646 294380 158652
rect 294328 149116 294380 149122
rect 294328 149058 294380 149064
rect 294340 140842 294368 149058
rect 294248 140814 294368 140842
rect 294248 140758 294276 140814
rect 294236 140752 294288 140758
rect 294236 140694 294288 140700
rect 294420 140752 294472 140758
rect 294420 140694 294472 140700
rect 294432 139398 294460 140694
rect 294420 139392 294472 139398
rect 294420 139334 294472 139340
rect 294420 129804 294472 129810
rect 294420 129746 294472 129752
rect 294432 121514 294460 129746
rect 294328 121508 294380 121514
rect 294328 121450 294380 121456
rect 294420 121508 294472 121514
rect 294420 121450 294472 121456
rect 294340 109750 294368 121450
rect 294328 109744 294380 109750
rect 294328 109686 294380 109692
rect 294328 102196 294380 102202
rect 294328 102138 294380 102144
rect 294340 85610 294368 102138
rect 295246 87544 295302 87553
rect 295246 87479 295302 87488
rect 295260 87009 295288 87479
rect 295246 87000 295302 87009
rect 295246 86935 295302 86944
rect 294236 85604 294288 85610
rect 294236 85546 294288 85552
rect 294328 85604 294380 85610
rect 294328 85546 294380 85552
rect 294248 64870 294276 85546
rect 295246 75984 295302 75993
rect 295246 75919 295302 75928
rect 295260 75585 295288 75919
rect 295246 75576 295302 75585
rect 295246 75511 295302 75520
rect 294236 64864 294288 64870
rect 294236 64806 294288 64812
rect 294236 46980 294288 46986
rect 294236 46922 294288 46928
rect 294248 45558 294276 46922
rect 294236 45552 294288 45558
rect 294236 45494 294288 45500
rect 294420 26308 294472 26314
rect 294420 26250 294472 26256
rect 294432 17898 294460 26250
rect 294340 17870 294460 17898
rect 294340 13326 294368 17870
rect 294328 13320 294380 13326
rect 294328 13262 294380 13268
rect 294052 9784 294104 9790
rect 294052 9726 294104 9732
rect 293960 7132 294012 7138
rect 293960 7074 294012 7080
rect 295352 7070 295380 340054
rect 295720 335696 295748 340054
rect 295444 335668 295748 335696
rect 295444 9722 295472 335668
rect 296272 335594 296300 340054
rect 295536 335566 296300 335594
rect 295536 328438 295564 335566
rect 295524 328432 295576 328438
rect 295524 328374 295576 328380
rect 295708 328432 295760 328438
rect 295708 328374 295760 328380
rect 295720 323490 295748 328374
rect 295628 323462 295748 323490
rect 295628 302190 295656 323462
rect 295616 302184 295668 302190
rect 295616 302126 295668 302132
rect 295708 302116 295760 302122
rect 295708 302058 295760 302064
rect 295720 288522 295748 302058
rect 295708 288516 295760 288522
rect 295708 288458 295760 288464
rect 295524 287088 295576 287094
rect 295524 287030 295576 287036
rect 295536 280838 295564 287030
rect 295524 280832 295576 280838
rect 295524 280774 295576 280780
rect 295800 280832 295852 280838
rect 295800 280774 295852 280780
rect 295812 276049 295840 280774
rect 295614 276040 295670 276049
rect 295614 275975 295670 275984
rect 295798 276040 295854 276049
rect 295798 275975 295854 275984
rect 295628 267782 295656 275975
rect 295616 267776 295668 267782
rect 295616 267718 295668 267724
rect 295800 267776 295852 267782
rect 295800 267718 295852 267724
rect 295812 262970 295840 267718
rect 295720 262942 295840 262970
rect 295720 256698 295748 262942
rect 295708 256692 295760 256698
rect 295708 256634 295760 256640
rect 295892 256692 295944 256698
rect 295892 256634 295944 256640
rect 295904 247081 295932 256634
rect 295522 247072 295578 247081
rect 295522 247007 295578 247016
rect 295890 247072 295946 247081
rect 295890 247007 295946 247016
rect 295536 241482 295564 247007
rect 295536 241454 295656 241482
rect 295536 222222 295564 222253
rect 295628 222222 295656 241454
rect 295524 222216 295576 222222
rect 295616 222216 295668 222222
rect 295576 222164 295616 222170
rect 295524 222158 295668 222164
rect 295536 222142 295656 222158
rect 295536 202910 295564 202941
rect 295628 202910 295656 222142
rect 295524 202904 295576 202910
rect 295616 202904 295668 202910
rect 295576 202852 295616 202858
rect 295524 202846 295668 202852
rect 295536 202830 295656 202846
rect 295628 186454 295656 202830
rect 295616 186448 295668 186454
rect 295616 186390 295668 186396
rect 295524 186312 295576 186318
rect 295524 186254 295576 186260
rect 295536 178770 295564 186254
rect 295524 178764 295576 178770
rect 295524 178706 295576 178712
rect 295708 178764 295760 178770
rect 295708 178706 295760 178712
rect 295720 160138 295748 178706
rect 295616 160132 295668 160138
rect 295616 160074 295668 160080
rect 295708 160132 295760 160138
rect 295708 160074 295760 160080
rect 295628 153202 295656 160074
rect 295524 153196 295576 153202
rect 295524 153138 295576 153144
rect 295616 153196 295668 153202
rect 295616 153138 295668 153144
rect 295536 140758 295564 153138
rect 295524 140752 295576 140758
rect 295524 140694 295576 140700
rect 295616 131164 295668 131170
rect 295616 131106 295668 131112
rect 295628 103494 295656 131106
rect 295616 103488 295668 103494
rect 295616 103430 295668 103436
rect 295616 93900 295668 93906
rect 295616 93842 295668 93848
rect 295628 90386 295656 93842
rect 295628 90358 295748 90386
rect 295720 75954 295748 90358
rect 296626 87136 296682 87145
rect 296626 87071 296682 87080
rect 296640 87009 296668 87071
rect 296626 87000 296682 87009
rect 296626 86935 296682 86944
rect 295524 75948 295576 75954
rect 295524 75890 295576 75896
rect 295708 75948 295760 75954
rect 295708 75890 295760 75896
rect 295536 28966 295564 75890
rect 296626 29608 296682 29617
rect 296626 29543 296682 29552
rect 296640 29345 296668 29543
rect 296626 29336 296682 29345
rect 296626 29271 296682 29280
rect 295524 28960 295576 28966
rect 295524 28902 295576 28908
rect 295616 28960 295668 28966
rect 295616 28902 295668 28908
rect 295628 12510 295656 28902
rect 295616 12504 295668 12510
rect 295616 12446 295668 12452
rect 295432 9716 295484 9722
rect 295432 9658 295484 9664
rect 295340 7064 295392 7070
rect 295340 7006 295392 7012
rect 296732 6730 296760 340054
rect 297284 335696 297312 340054
rect 297916 337204 297968 337210
rect 297916 337146 297968 337152
rect 296824 335668 297312 335696
rect 296824 328438 296852 335668
rect 296812 328432 296864 328438
rect 296812 328374 296864 328380
rect 296996 328432 297048 328438
rect 296996 328374 297048 328380
rect 297008 323490 297036 328374
rect 296916 323462 297036 323490
rect 296916 298194 296944 323462
rect 296824 298166 296944 298194
rect 296824 292602 296852 298166
rect 296812 292596 296864 292602
rect 296812 292538 296864 292544
rect 296904 292528 296956 292534
rect 296904 292470 296956 292476
rect 296916 287026 296944 292470
rect 296904 287020 296956 287026
rect 296904 286962 296956 286968
rect 297088 276072 297140 276078
rect 297088 276014 297140 276020
rect 297100 267730 297128 276014
rect 297008 267702 297128 267730
rect 297008 251326 297036 267702
rect 296996 251320 297048 251326
rect 296996 251262 297048 251268
rect 296812 251116 296864 251122
rect 296812 251058 296864 251064
rect 296824 241482 296852 251058
rect 296824 241454 296944 241482
rect 296824 222222 296852 222253
rect 296916 222222 296944 241454
rect 296812 222216 296864 222222
rect 296904 222216 296956 222222
rect 296864 222164 296904 222170
rect 296812 222158 296956 222164
rect 296824 222142 296944 222158
rect 296824 202910 296852 202941
rect 296916 202910 296944 222142
rect 296812 202904 296864 202910
rect 296904 202904 296956 202910
rect 296864 202852 296904 202858
rect 296812 202846 296956 202852
rect 296824 202830 296944 202846
rect 296916 186454 296944 202830
rect 296904 186448 296956 186454
rect 296904 186390 296956 186396
rect 296812 186312 296864 186318
rect 296812 186254 296864 186260
rect 296824 178770 296852 186254
rect 296812 178764 296864 178770
rect 296812 178706 296864 178712
rect 296996 178764 297048 178770
rect 296996 178706 297048 178712
rect 297008 160138 297036 178706
rect 296904 160132 296956 160138
rect 296904 160074 296956 160080
rect 296996 160132 297048 160138
rect 296996 160074 297048 160080
rect 296916 151722 296944 160074
rect 296824 151694 296944 151722
rect 296824 138038 296852 151694
rect 296812 138032 296864 138038
rect 296812 137974 296864 137980
rect 297272 138032 297324 138038
rect 297272 137974 297324 137980
rect 297284 131186 297312 137974
rect 297192 131158 297312 131186
rect 297192 131102 297220 131158
rect 297180 131096 297232 131102
rect 297180 131038 297232 131044
rect 296904 121508 296956 121514
rect 296904 121450 296956 121456
rect 296916 114646 296944 121450
rect 296904 114640 296956 114646
rect 296904 114582 296956 114588
rect 296812 114504 296864 114510
rect 296812 114446 296864 114452
rect 296824 113150 296852 114446
rect 296812 113144 296864 113150
rect 296812 113086 296864 113092
rect 296812 103556 296864 103562
rect 296812 103498 296864 103504
rect 296824 103442 296852 103498
rect 296824 103426 296944 103442
rect 296824 103420 296956 103426
rect 296824 103414 296904 103420
rect 296904 103362 296956 103368
rect 297088 103420 297140 103426
rect 297088 103362 297140 103368
rect 297100 95146 297128 103362
rect 297008 95118 297128 95146
rect 297008 84318 297036 95118
rect 296996 84312 297048 84318
rect 296996 84254 297048 84260
rect 297088 84244 297140 84250
rect 297088 84186 297140 84192
rect 297100 74662 297128 84186
rect 296812 74656 296864 74662
rect 296812 74598 296864 74604
rect 297088 74656 297140 74662
rect 297088 74598 297140 74604
rect 296824 66298 296852 74598
rect 296812 66292 296864 66298
rect 296812 66234 296864 66240
rect 296904 66156 296956 66162
rect 296904 66098 296956 66104
rect 296916 55162 296944 66098
rect 296824 55134 296944 55162
rect 296824 38690 296852 55134
rect 296812 38684 296864 38690
rect 296812 38626 296864 38632
rect 296904 38548 296956 38554
rect 296904 38490 296956 38496
rect 296916 13394 296944 38490
rect 296904 13388 296956 13394
rect 296904 13330 296956 13336
rect 296720 6724 296772 6730
rect 296720 6666 296772 6672
rect 297364 6656 297416 6662
rect 297364 6598 297416 6604
rect 295892 6588 295944 6594
rect 295892 6530 295944 6536
rect 294328 6316 294380 6322
rect 294328 6258 294380 6264
rect 290740 5432 290792 5438
rect 290740 5374 290792 5380
rect 290464 3120 290516 3126
rect 290464 3062 290516 3068
rect 290752 480 290780 5374
rect 291936 3256 291988 3262
rect 291936 3198 291988 3204
rect 291948 480 291976 3198
rect 293132 3052 293184 3058
rect 293132 2994 293184 3000
rect 293144 480 293172 2994
rect 294340 480 294368 6258
rect 295904 4146 295932 6530
rect 295892 4140 295944 4146
rect 295892 4082 295944 4088
rect 296720 4140 296772 4146
rect 296720 4082 296772 4088
rect 295524 3120 295576 3126
rect 295524 3062 295576 3068
rect 295536 480 295564 3062
rect 296732 480 296760 4082
rect 297376 4078 297404 6598
rect 297824 5500 297876 5506
rect 297824 5442 297876 5448
rect 297364 4072 297416 4078
rect 297364 4014 297416 4020
rect 297836 4026 297864 5442
rect 297928 4146 297956 337146
rect 298098 29336 298154 29345
rect 298098 29271 298154 29280
rect 298112 28937 298140 29271
rect 298098 28928 298154 28937
rect 298098 28863 298154 28872
rect 298006 16824 298062 16833
rect 298062 16782 298140 16810
rect 298006 16759 298062 16768
rect 298112 16697 298140 16782
rect 298098 16688 298154 16697
rect 298098 16623 298154 16632
rect 298204 12306 298232 340054
rect 298388 340054 298586 340082
rect 298664 340054 299046 340082
rect 298284 335640 298336 335646
rect 298284 335582 298336 335588
rect 298296 13462 298324 335582
rect 298284 13456 298336 13462
rect 298284 13398 298336 13404
rect 298192 12300 298244 12306
rect 298192 12242 298244 12248
rect 298388 6798 298416 340054
rect 298664 335646 298692 340054
rect 298652 335640 298704 335646
rect 298652 335582 298704 335588
rect 299584 331294 299612 340068
rect 299768 340054 300058 340082
rect 300228 340054 300518 340082
rect 300964 340054 301070 340082
rect 301240 340054 301530 340082
rect 301700 340054 301990 340082
rect 302344 340054 302542 340082
rect 302712 340054 303002 340082
rect 303080 340054 303462 340082
rect 303724 340054 303922 340082
rect 304184 340054 304474 340082
rect 304644 340054 304934 340082
rect 305104 340054 305394 340082
rect 305656 340054 305946 340082
rect 299572 331288 299624 331294
rect 299768 331242 299796 340054
rect 299572 331230 299624 331236
rect 299676 331214 299796 331242
rect 299572 331152 299624 331158
rect 299572 331094 299624 331100
rect 299480 331084 299532 331090
rect 299480 331026 299532 331032
rect 299492 241466 299520 331026
rect 299480 241460 299532 241466
rect 299480 241402 299532 241408
rect 299480 231872 299532 231878
rect 299480 231814 299532 231820
rect 299492 222154 299520 231814
rect 299480 222148 299532 222154
rect 299480 222090 299532 222096
rect 299480 212560 299532 212566
rect 299480 212502 299532 212508
rect 299492 202842 299520 212502
rect 299480 202836 299532 202842
rect 299480 202778 299532 202784
rect 299480 193248 299532 193254
rect 299480 193190 299532 193196
rect 299492 6866 299520 193190
rect 299584 12374 299612 331094
rect 299676 331090 299704 331214
rect 300228 331158 300256 340054
rect 300860 335640 300912 335646
rect 300860 335582 300912 335588
rect 299756 331152 299808 331158
rect 299756 331094 299808 331100
rect 300216 331152 300268 331158
rect 300216 331094 300268 331100
rect 299664 331084 299716 331090
rect 299664 331026 299716 331032
rect 299768 327162 299796 331094
rect 299768 327134 299888 327162
rect 299860 327078 299888 327134
rect 299848 327072 299900 327078
rect 299848 327014 299900 327020
rect 299848 317484 299900 317490
rect 299848 317426 299900 317432
rect 299860 312066 299888 317426
rect 299676 312038 299888 312066
rect 299676 308122 299704 312038
rect 299676 308094 299888 308122
rect 299860 289882 299888 308094
rect 299756 289876 299808 289882
rect 299756 289818 299808 289824
rect 299848 289876 299900 289882
rect 299848 289818 299900 289824
rect 299768 285138 299796 289818
rect 299768 285110 299980 285138
rect 299952 282826 299980 285110
rect 299768 282798 299980 282826
rect 299768 280242 299796 282798
rect 299768 280214 299888 280242
rect 299860 259418 299888 280214
rect 299848 259412 299900 259418
rect 299848 259354 299900 259360
rect 300032 259412 300084 259418
rect 300032 259354 300084 259360
rect 300044 240174 300072 259354
rect 299940 240168 299992 240174
rect 299940 240110 299992 240116
rect 300032 240168 300084 240174
rect 300032 240110 300084 240116
rect 299952 231878 299980 240110
rect 299940 231872 299992 231878
rect 299940 231814 299992 231820
rect 299756 231804 299808 231810
rect 299756 231746 299808 231752
rect 299768 222222 299796 231746
rect 299756 222216 299808 222222
rect 299756 222158 299808 222164
rect 299940 222216 299992 222222
rect 299940 222158 299992 222164
rect 299952 212634 299980 222158
rect 299940 212628 299992 212634
rect 299940 212570 299992 212576
rect 299756 212492 299808 212498
rect 299756 212434 299808 212440
rect 299768 202910 299796 212434
rect 299756 202904 299808 202910
rect 299756 202846 299808 202852
rect 299940 202904 299992 202910
rect 299940 202846 299992 202852
rect 299952 193338 299980 202846
rect 299952 193310 300072 193338
rect 300044 191842 300072 193310
rect 299860 191814 300072 191842
rect 299860 188494 299888 191814
rect 299848 188488 299900 188494
rect 299848 188430 299900 188436
rect 299848 183592 299900 183598
rect 299848 183534 299900 183540
rect 299860 180810 299888 183534
rect 299848 180804 299900 180810
rect 299848 180746 299900 180752
rect 299848 171148 299900 171154
rect 299848 171090 299900 171096
rect 299860 154562 299888 171090
rect 299756 154556 299808 154562
rect 299756 154498 299808 154504
rect 299848 154556 299900 154562
rect 299848 154498 299900 154504
rect 299768 149546 299796 154498
rect 299768 149518 299888 149546
rect 299860 128602 299888 149518
rect 299860 128574 299980 128602
rect 299952 128194 299980 128574
rect 299860 128166 299980 128194
rect 299860 124166 299888 128166
rect 299848 124160 299900 124166
rect 299848 124102 299900 124108
rect 299848 114572 299900 114578
rect 299848 114514 299900 114520
rect 299860 96642 299888 114514
rect 299768 96614 299888 96642
rect 299768 90386 299796 96614
rect 299768 90358 299888 90386
rect 299860 85542 299888 90358
rect 299848 85536 299900 85542
rect 299848 85478 299900 85484
rect 299848 75948 299900 75954
rect 299848 75890 299900 75896
rect 299860 67658 299888 75890
rect 299756 67652 299808 67658
rect 299756 67594 299808 67600
rect 299848 67652 299900 67658
rect 299848 67594 299900 67600
rect 299768 57984 299796 67594
rect 299676 57956 299796 57984
rect 299676 56574 299704 57956
rect 299664 56568 299716 56574
rect 299664 56510 299716 56516
rect 299756 45620 299808 45626
rect 299756 45562 299808 45568
rect 299768 45490 299796 45562
rect 299756 45484 299808 45490
rect 299756 45426 299808 45432
rect 299848 45484 299900 45490
rect 299848 45426 299900 45432
rect 299860 32314 299888 45426
rect 299768 32286 299888 32314
rect 299768 13530 299796 32286
rect 299756 13524 299808 13530
rect 299756 13466 299808 13472
rect 299572 12368 299624 12374
rect 299572 12310 299624 12316
rect 299480 6860 299532 6866
rect 299480 6802 299532 6808
rect 298376 6792 298428 6798
rect 298376 6734 298428 6740
rect 298100 6724 298152 6730
rect 298100 6666 298152 6672
rect 297916 4140 297968 4146
rect 297916 4082 297968 4088
rect 297836 3998 297956 4026
rect 298112 4010 298140 6666
rect 300872 6118 300900 335582
rect 300964 12442 300992 340054
rect 301240 335646 301268 340054
rect 301228 335640 301280 335646
rect 301228 335582 301280 335588
rect 301700 331906 301728 340054
rect 302240 335708 302292 335714
rect 302240 335650 302292 335656
rect 301044 331900 301096 331906
rect 301044 331842 301096 331848
rect 301688 331900 301740 331906
rect 301688 331842 301740 331848
rect 301056 327162 301084 331842
rect 301056 327134 301176 327162
rect 301148 327078 301176 327134
rect 301136 327072 301188 327078
rect 301136 327014 301188 327020
rect 301320 327072 301372 327078
rect 301320 327014 301372 327020
rect 301332 317529 301360 327014
rect 301318 317520 301374 317529
rect 301318 317455 301374 317464
rect 301226 317384 301282 317393
rect 301226 317319 301282 317328
rect 301240 307834 301268 317319
rect 301044 307828 301096 307834
rect 301044 307770 301096 307776
rect 301228 307828 301280 307834
rect 301228 307770 301280 307776
rect 301056 292602 301084 307770
rect 301044 292596 301096 292602
rect 301044 292538 301096 292544
rect 301136 292528 301188 292534
rect 301136 292470 301188 292476
rect 301148 283014 301176 292470
rect 301136 283008 301188 283014
rect 301136 282950 301188 282956
rect 301044 282872 301096 282878
rect 301044 282814 301096 282820
rect 301056 269142 301084 282814
rect 301044 269136 301096 269142
rect 301044 269078 301096 269084
rect 301228 269136 301280 269142
rect 301228 269078 301280 269084
rect 301240 246242 301268 269078
rect 301056 246214 301268 246242
rect 301056 241505 301084 246214
rect 301042 241496 301098 241505
rect 301042 241431 301098 241440
rect 301134 241360 301190 241369
rect 301134 241295 301190 241304
rect 301148 231946 301176 241295
rect 301136 231940 301188 231946
rect 301136 231882 301188 231888
rect 301044 231804 301096 231810
rect 301044 231746 301096 231752
rect 301056 222193 301084 231746
rect 301042 222184 301098 222193
rect 301042 222119 301098 222128
rect 301134 222048 301190 222057
rect 301134 221983 301190 221992
rect 301148 212634 301176 221983
rect 301136 212628 301188 212634
rect 301136 212570 301188 212576
rect 301044 212492 301096 212498
rect 301044 212434 301096 212440
rect 301056 202881 301084 212434
rect 301042 202872 301098 202881
rect 301042 202807 301098 202816
rect 301134 202736 301190 202745
rect 301134 202671 301190 202680
rect 301148 196602 301176 202671
rect 301148 196574 301268 196602
rect 301240 183598 301268 196574
rect 301044 183592 301096 183598
rect 301044 183534 301096 183540
rect 301228 183592 301280 183598
rect 301228 183534 301280 183540
rect 301056 180810 301084 183534
rect 301044 180804 301096 180810
rect 301044 180746 301096 180752
rect 301044 171148 301096 171154
rect 301044 171090 301096 171096
rect 301056 154494 301084 171090
rect 301044 154488 301096 154494
rect 301044 154430 301096 154436
rect 301228 154488 301280 154494
rect 301228 154430 301280 154436
rect 301240 144945 301268 154430
rect 301042 144936 301098 144945
rect 301042 144871 301098 144880
rect 301226 144936 301282 144945
rect 301226 144871 301282 144880
rect 301056 143546 301084 144871
rect 301044 143540 301096 143546
rect 301044 143482 301096 143488
rect 301228 143540 301280 143546
rect 301228 143482 301280 143488
rect 301240 138530 301268 143482
rect 301148 138502 301268 138530
rect 301148 111058 301176 138502
rect 301148 111030 301268 111058
rect 301240 103494 301268 111030
rect 301228 103488 301280 103494
rect 301228 103430 301280 103436
rect 301136 93900 301188 93906
rect 301136 93842 301188 93848
rect 301148 90658 301176 93842
rect 301148 90630 301268 90658
rect 301240 85542 301268 90630
rect 301044 85536 301096 85542
rect 301044 85478 301096 85484
rect 301228 85536 301280 85542
rect 301228 85478 301280 85484
rect 301056 84130 301084 85478
rect 301056 84102 301268 84130
rect 301240 66337 301268 84102
rect 301226 66328 301282 66337
rect 301226 66263 301282 66272
rect 301226 66056 301282 66065
rect 301226 65991 301282 66000
rect 301240 56710 301268 65991
rect 301044 56704 301096 56710
rect 301044 56646 301096 56652
rect 301228 56704 301280 56710
rect 301228 56646 301280 56652
rect 301056 56574 301084 56646
rect 301044 56568 301096 56574
rect 301044 56510 301096 56516
rect 301044 46980 301096 46986
rect 301044 46922 301096 46928
rect 301056 38690 301084 46922
rect 301044 38684 301096 38690
rect 301044 38626 301096 38632
rect 301320 38616 301372 38622
rect 301320 38558 301372 38564
rect 301332 35902 301360 38558
rect 301320 35896 301372 35902
rect 301320 35838 301372 35844
rect 301136 26308 301188 26314
rect 301136 26250 301188 26256
rect 301148 13598 301176 26250
rect 301136 13592 301188 13598
rect 301136 13534 301188 13540
rect 300952 12436 301004 12442
rect 300952 12378 301004 12384
rect 300860 6112 300912 6118
rect 300860 6054 300912 6060
rect 302252 6050 302280 335650
rect 302344 11694 302372 340054
rect 302712 335714 302740 340054
rect 302700 335708 302752 335714
rect 302700 335650 302752 335656
rect 303080 334762 303108 340054
rect 303160 337952 303212 337958
rect 303160 337894 303212 337900
rect 303068 334756 303120 334762
rect 303068 334698 303120 334704
rect 303172 334642 303200 337894
rect 303620 335640 303672 335646
rect 303620 335582 303672 335588
rect 302896 334614 303200 334642
rect 302516 328500 302568 328506
rect 302516 328442 302568 328448
rect 302528 318850 302556 328442
rect 302516 318844 302568 318850
rect 302516 318786 302568 318792
rect 302608 318844 302660 318850
rect 302608 318786 302660 318792
rect 302620 292618 302648 318786
rect 302528 292590 302648 292618
rect 302528 289814 302556 292590
rect 302516 289808 302568 289814
rect 302516 289750 302568 289756
rect 302700 289808 302752 289814
rect 302700 289750 302752 289756
rect 302712 269210 302740 289750
rect 302700 269204 302752 269210
rect 302700 269146 302752 269152
rect 302608 269136 302660 269142
rect 302608 269078 302660 269084
rect 302620 259418 302648 269078
rect 302608 259412 302660 259418
rect 302608 259354 302660 259360
rect 302792 259412 302844 259418
rect 302792 259354 302844 259360
rect 302804 240174 302832 259354
rect 302700 240168 302752 240174
rect 302700 240110 302752 240116
rect 302792 240168 302844 240174
rect 302792 240110 302844 240116
rect 302712 231860 302740 240110
rect 302620 231832 302740 231860
rect 302620 222306 302648 231832
rect 302620 222278 302740 222306
rect 302712 212650 302740 222278
rect 302712 212622 302832 212650
rect 302804 212378 302832 212622
rect 302620 212350 302832 212378
rect 302620 202994 302648 212350
rect 302620 202966 302740 202994
rect 302712 193322 302740 202966
rect 302700 193316 302752 193322
rect 302700 193258 302752 193264
rect 302516 193180 302568 193186
rect 302516 193122 302568 193128
rect 302528 183666 302556 193122
rect 302516 183660 302568 183666
rect 302516 183602 302568 183608
rect 302608 183592 302660 183598
rect 302608 183534 302660 183540
rect 302620 180810 302648 183534
rect 302608 180804 302660 180810
rect 302608 180746 302660 180752
rect 302608 171148 302660 171154
rect 302608 171090 302660 171096
rect 302620 161430 302648 171090
rect 302516 161424 302568 161430
rect 302516 161366 302568 161372
rect 302608 161424 302660 161430
rect 302608 161366 302660 161372
rect 302528 144922 302556 161366
rect 302528 144894 302648 144922
rect 302620 128382 302648 144894
rect 302608 128376 302660 128382
rect 302608 128318 302660 128324
rect 302608 128240 302660 128246
rect 302608 128182 302660 128188
rect 302620 75954 302648 128182
rect 302516 75948 302568 75954
rect 302516 75890 302568 75896
rect 302608 75948 302660 75954
rect 302608 75890 302660 75896
rect 302528 53122 302556 75890
rect 302528 53094 302648 53122
rect 302620 38690 302648 53094
rect 302516 38684 302568 38690
rect 302516 38626 302568 38632
rect 302608 38684 302660 38690
rect 302608 38626 302660 38632
rect 302528 29102 302556 38626
rect 302516 29096 302568 29102
rect 302516 29038 302568 29044
rect 302516 28960 302568 28966
rect 302516 28902 302568 28908
rect 302528 17898 302556 28902
rect 302528 17870 302648 17898
rect 302620 13666 302648 17870
rect 302608 13660 302660 13666
rect 302608 13602 302660 13608
rect 302332 11688 302384 11694
rect 302332 11630 302384 11636
rect 302240 6044 302292 6050
rect 302240 5986 302292 5992
rect 301412 4412 301464 4418
rect 301412 4354 301464 4360
rect 300308 4140 300360 4146
rect 300308 4082 300360 4088
rect 297928 480 297956 3998
rect 298100 4004 298152 4010
rect 298100 3946 298152 3952
rect 299112 3392 299164 3398
rect 299112 3334 299164 3340
rect 299124 480 299152 3334
rect 300320 480 300348 4082
rect 301424 480 301452 4354
rect 302608 4072 302660 4078
rect 302608 4014 302660 4020
rect 302620 480 302648 4014
rect 302896 3398 302924 334614
rect 303632 5982 303660 335582
rect 303724 11626 303752 340054
rect 304184 335646 304212 340054
rect 304172 335640 304224 335646
rect 304172 335582 304224 335588
rect 304644 328506 304672 340054
rect 305000 335640 305052 335646
rect 305000 335582 305052 335588
rect 303896 328500 303948 328506
rect 303896 328442 303948 328448
rect 304632 328500 304684 328506
rect 304632 328442 304684 328448
rect 303908 311930 303936 328442
rect 303816 311902 303936 311930
rect 303816 311794 303844 311902
rect 303816 311766 303936 311794
rect 303908 292482 303936 311766
rect 303816 292454 303936 292482
rect 303816 292210 303844 292454
rect 303816 292182 303936 292210
rect 303908 176746 303936 292182
rect 303816 176718 303936 176746
rect 303816 176610 303844 176718
rect 303816 176582 303936 176610
rect 303908 80102 303936 176582
rect 303896 80096 303948 80102
rect 303896 80038 303948 80044
rect 303896 79960 303948 79966
rect 303896 79902 303948 79908
rect 303908 77246 303936 79902
rect 303896 77240 303948 77246
rect 303896 77182 303948 77188
rect 303988 77240 304040 77246
rect 303988 77182 304040 77188
rect 304000 58002 304028 77182
rect 303896 57996 303948 58002
rect 303896 57938 303948 57944
rect 303988 57996 304040 58002
rect 303988 57938 304040 57944
rect 303908 46986 303936 57938
rect 303804 46980 303856 46986
rect 303804 46922 303856 46928
rect 303896 46980 303948 46986
rect 303896 46922 303948 46928
rect 303816 38622 303844 46922
rect 303804 38616 303856 38622
rect 303804 38558 303856 38564
rect 303896 32428 303948 32434
rect 303896 32370 303948 32376
rect 303908 13734 303936 32370
rect 303896 13728 303948 13734
rect 303896 13670 303948 13676
rect 303712 11620 303764 11626
rect 303712 11562 303764 11568
rect 303620 5976 303672 5982
rect 303620 5918 303672 5924
rect 305012 5914 305040 335582
rect 305104 11558 305132 340054
rect 305656 335646 305684 340054
rect 306196 338020 306248 338026
rect 306196 337962 306248 337968
rect 305644 335640 305696 335646
rect 305644 335582 305696 335588
rect 305092 11552 305144 11558
rect 305092 11494 305144 11500
rect 305000 5908 305052 5914
rect 305000 5850 305052 5856
rect 305000 4344 305052 4350
rect 305000 4286 305052 4292
rect 302884 3392 302936 3398
rect 302884 3334 302936 3340
rect 303804 3324 303856 3330
rect 303804 3266 303856 3272
rect 303816 480 303844 3266
rect 305012 480 305040 4286
rect 306208 480 306236 337962
rect 306392 333418 306420 340068
rect 306668 340054 306866 340082
rect 307036 340054 307418 340082
rect 307878 340054 307984 340082
rect 306392 333390 306604 333418
rect 306472 331084 306524 331090
rect 306472 331026 306524 331032
rect 306380 160064 306432 160070
rect 306380 160006 306432 160012
rect 306392 142186 306420 160006
rect 306380 142180 306432 142186
rect 306380 142122 306432 142128
rect 306286 76120 306342 76129
rect 306286 76055 306342 76064
rect 306300 75857 306328 76055
rect 306286 75848 306342 75857
rect 306286 75783 306342 75792
rect 306378 40216 306434 40225
rect 306378 40151 306380 40160
rect 306432 40151 306434 40160
rect 306380 40122 306432 40128
rect 306378 28928 306434 28937
rect 306378 28863 306380 28872
rect 306432 28863 306434 28872
rect 306380 28834 306432 28840
rect 306484 11490 306512 331026
rect 306576 13802 306604 333390
rect 306668 331090 306696 340054
rect 307036 331242 307064 340054
rect 307760 337748 307812 337754
rect 307760 337690 307812 337696
rect 307772 337657 307800 337690
rect 307758 337648 307814 337657
rect 307758 337583 307814 337592
rect 307760 335640 307812 335646
rect 307760 335582 307812 335588
rect 306760 331214 307064 331242
rect 306656 331084 306708 331090
rect 306656 331026 306708 331032
rect 306760 318850 306788 331214
rect 306748 318844 306800 318850
rect 306748 318786 306800 318792
rect 306840 318844 306892 318850
rect 306840 318786 306892 318792
rect 306852 312610 306880 318786
rect 306852 312582 306972 312610
rect 306944 294642 306972 312582
rect 306748 294636 306800 294642
rect 306748 294578 306800 294584
rect 306932 294636 306984 294642
rect 306932 294578 306984 294584
rect 306760 289814 306788 294578
rect 306748 289808 306800 289814
rect 306748 289750 306800 289756
rect 306932 289808 306984 289814
rect 306932 289750 306984 289756
rect 306944 269210 306972 289750
rect 306932 269204 306984 269210
rect 306932 269146 306984 269152
rect 306840 269136 306892 269142
rect 306840 269078 306892 269084
rect 306852 241602 306880 269078
rect 306840 241596 306892 241602
rect 306840 241538 306892 241544
rect 306840 241460 306892 241466
rect 306840 241402 306892 241408
rect 306852 222358 306880 241402
rect 306840 222352 306892 222358
rect 306840 222294 306892 222300
rect 306932 222352 306984 222358
rect 306932 222294 306984 222300
rect 306944 212548 306972 222294
rect 306852 212520 306972 212548
rect 306852 202994 306880 212520
rect 306852 202966 306972 202994
rect 306944 193338 306972 202966
rect 306944 193310 307064 193338
rect 307036 191842 307064 193310
rect 306852 191814 307064 191842
rect 306852 188494 306880 191814
rect 306840 188488 306892 188494
rect 306840 188430 306892 188436
rect 306840 183592 306892 183598
rect 306840 183534 306892 183540
rect 306852 176746 306880 183534
rect 306852 176718 306972 176746
rect 306944 171154 306972 176718
rect 306656 171148 306708 171154
rect 306656 171090 306708 171096
rect 306932 171148 306984 171154
rect 306932 171090 306984 171096
rect 306668 171034 306696 171090
rect 306668 171006 306788 171034
rect 306760 161514 306788 171006
rect 306760 161486 306880 161514
rect 306852 160070 306880 161486
rect 306840 160064 306892 160070
rect 306840 160006 306892 160012
rect 307024 142180 307076 142186
rect 307024 142122 307076 142128
rect 307036 133958 307064 142122
rect 307024 133952 307076 133958
rect 307024 133894 307076 133900
rect 307024 133816 307076 133822
rect 307024 133758 307076 133764
rect 307036 124273 307064 133758
rect 306838 124264 306894 124273
rect 306838 124199 306894 124208
rect 307022 124264 307078 124273
rect 307022 124199 307078 124208
rect 306852 124166 306880 124199
rect 306840 124160 306892 124166
rect 306840 124102 306892 124108
rect 306748 113280 306800 113286
rect 306800 113228 306880 113234
rect 306748 113222 306880 113228
rect 306760 113206 306880 113222
rect 306852 113150 306880 113206
rect 306840 113144 306892 113150
rect 306840 113086 306892 113092
rect 307024 113144 307076 113150
rect 307024 113086 307076 113092
rect 307036 103601 307064 113086
rect 306838 103592 306894 103601
rect 306838 103527 306894 103536
rect 307022 103592 307078 103601
rect 307022 103527 307078 103536
rect 306852 103494 306880 103527
rect 306840 103488 306892 103494
rect 306840 103430 306892 103436
rect 306840 93900 306892 93906
rect 306840 93842 306892 93848
rect 306852 85542 306880 93842
rect 306656 85536 306708 85542
rect 306656 85478 306708 85484
rect 306840 85536 306892 85542
rect 306840 85478 306892 85484
rect 306668 65822 306696 85478
rect 306656 65816 306708 65822
rect 306656 65758 306708 65764
rect 306840 65816 306892 65822
rect 306840 65758 306892 65764
rect 306852 46986 306880 65758
rect 306748 46980 306800 46986
rect 306748 46922 306800 46928
rect 306840 46980 306892 46986
rect 306840 46922 306892 46928
rect 306760 38622 306788 46922
rect 306748 38616 306800 38622
rect 306748 38558 306800 38564
rect 306840 38616 306892 38622
rect 306840 38558 306892 38564
rect 306852 19378 306880 38558
rect 306748 19372 306800 19378
rect 306748 19314 306800 19320
rect 306840 19372 306892 19378
rect 306840 19314 306892 19320
rect 306564 13796 306616 13802
rect 306564 13738 306616 13744
rect 306472 11484 306524 11490
rect 306472 11426 306524 11432
rect 306760 9790 306788 19314
rect 306748 9784 306800 9790
rect 306748 9726 306800 9732
rect 306656 9716 306708 9722
rect 306656 9658 306708 9664
rect 306668 5846 306696 9658
rect 306656 5840 306708 5846
rect 306656 5782 306708 5788
rect 307772 5778 307800 335582
rect 307956 13054 307984 340054
rect 308048 340054 308338 340082
rect 308600 340054 308890 340082
rect 309244 340054 309350 340082
rect 309428 340054 309810 340082
rect 310072 340054 310362 340082
rect 310624 340054 310822 340082
rect 311084 340054 311282 340082
rect 311544 340054 311834 340082
rect 312004 340054 312294 340082
rect 307944 13048 307996 13054
rect 307944 12990 307996 12996
rect 308048 11422 308076 340054
rect 308600 335646 308628 340054
rect 308588 335640 308640 335646
rect 308588 335582 308640 335588
rect 309140 335640 309192 335646
rect 309140 335582 309192 335588
rect 308036 11416 308088 11422
rect 308036 11358 308088 11364
rect 307760 5772 307812 5778
rect 307760 5714 307812 5720
rect 309152 5710 309180 335582
rect 309244 9450 309272 340054
rect 309428 11354 309456 340054
rect 309784 337340 309836 337346
rect 309784 337282 309836 337288
rect 309416 11348 309468 11354
rect 309416 11290 309468 11296
rect 309232 9444 309284 9450
rect 309232 9386 309284 9392
rect 309140 5704 309192 5710
rect 309140 5646 309192 5652
rect 308588 4276 308640 4282
rect 308588 4218 308640 4224
rect 307390 3360 307446 3369
rect 307390 3295 307446 3304
rect 307404 480 307432 3295
rect 308600 480 308628 4218
rect 309796 4078 309824 337282
rect 310072 335646 310100 340054
rect 310060 335640 310112 335646
rect 310060 335582 310112 335588
rect 310520 332104 310572 332110
rect 310520 332046 310572 332052
rect 310532 5642 310560 332046
rect 310624 9518 310652 340054
rect 311084 331242 311112 340054
rect 311544 332110 311572 340054
rect 311532 332104 311584 332110
rect 311532 332046 311584 332052
rect 310808 331214 311112 331242
rect 310808 321638 310836 331214
rect 310796 321632 310848 321638
rect 310796 321574 310848 321580
rect 310888 321496 310940 321502
rect 310888 321438 310940 321444
rect 310900 311982 310928 321438
rect 310888 311976 310940 311982
rect 310888 311918 310940 311924
rect 310704 307896 310756 307902
rect 310704 307838 310756 307844
rect 310716 307766 310744 307838
rect 310704 307760 310756 307766
rect 310704 307702 310756 307708
rect 310888 298172 310940 298178
rect 310888 298114 310940 298120
rect 310900 293078 310928 298114
rect 310888 293072 310940 293078
rect 310888 293014 310940 293020
rect 310888 282804 310940 282810
rect 310888 282746 310940 282752
rect 310900 278730 310928 282746
rect 310888 278724 310940 278730
rect 310888 278666 310940 278672
rect 310888 263492 310940 263498
rect 310888 263434 310940 263440
rect 310900 256086 310928 263434
rect 310888 256080 310940 256086
rect 310888 256022 310940 256028
rect 310704 251320 310756 251326
rect 310704 251262 310756 251268
rect 310716 251190 310744 251262
rect 310704 251184 310756 251190
rect 310704 251126 310756 251132
rect 310888 241528 310940 241534
rect 310888 241470 310940 241476
rect 310900 234734 310928 241470
rect 310888 234728 310940 234734
rect 310888 234670 310940 234676
rect 310796 234592 310848 234598
rect 310796 234534 310848 234540
rect 310808 231810 310836 234534
rect 310796 231804 310848 231810
rect 310796 231746 310848 231752
rect 310888 222216 310940 222222
rect 310888 222158 310940 222164
rect 310900 215422 310928 222158
rect 310888 215416 310940 215422
rect 310888 215358 310940 215364
rect 310796 215280 310848 215286
rect 310796 215222 310848 215228
rect 310808 212498 310836 215222
rect 310796 212492 310848 212498
rect 310796 212434 310848 212440
rect 310888 202904 310940 202910
rect 310888 202846 310940 202852
rect 310900 196110 310928 202846
rect 310888 196104 310940 196110
rect 310888 196046 310940 196052
rect 310796 195968 310848 195974
rect 310796 195910 310848 195916
rect 310808 193225 310836 195910
rect 310794 193216 310850 193225
rect 310794 193151 310850 193160
rect 311070 193216 311126 193225
rect 311070 193151 311126 193160
rect 311084 183598 311112 193151
rect 310888 183592 310940 183598
rect 310888 183534 310940 183540
rect 311072 183592 311124 183598
rect 311072 183534 311124 183540
rect 310900 176798 310928 183534
rect 310888 176792 310940 176798
rect 310888 176734 310940 176740
rect 310796 176656 310848 176662
rect 310796 176598 310848 176604
rect 310808 167074 310836 176598
rect 310796 167068 310848 167074
rect 310796 167010 310848 167016
rect 310888 166932 310940 166938
rect 310888 166874 310940 166880
rect 310900 153377 310928 166874
rect 310886 153368 310942 153377
rect 310886 153303 310942 153312
rect 310794 153232 310850 153241
rect 310794 153167 310796 153176
rect 310848 153167 310850 153176
rect 310796 153138 310848 153144
rect 310796 147620 310848 147626
rect 310796 147562 310848 147568
rect 310808 143562 310836 147562
rect 310808 143534 310928 143562
rect 310900 133906 310928 143534
rect 310900 133878 311020 133906
rect 310992 116113 311020 133878
rect 310978 116104 311034 116113
rect 310978 116039 311034 116048
rect 310794 115968 310850 115977
rect 310794 115903 310850 115912
rect 310808 109070 310836 115903
rect 310796 109064 310848 109070
rect 310796 109006 310848 109012
rect 310888 108996 310940 109002
rect 310888 108938 310940 108944
rect 310900 96830 310928 108938
rect 310888 96824 310940 96830
rect 310888 96766 310940 96772
rect 310796 96688 310848 96694
rect 310796 96630 310848 96636
rect 310808 95198 310836 96630
rect 310796 95192 310848 95198
rect 310796 95134 310848 95140
rect 310796 85604 310848 85610
rect 310796 85546 310848 85552
rect 310808 76158 310836 85546
rect 310796 76152 310848 76158
rect 310796 76094 310848 76100
rect 310796 76016 310848 76022
rect 310796 75958 310848 75964
rect 310808 75886 310836 75958
rect 310796 75880 310848 75886
rect 310796 75822 310848 75828
rect 310796 66360 310848 66366
rect 310796 66302 310848 66308
rect 310808 66230 310836 66302
rect 310796 66224 310848 66230
rect 310796 66166 310848 66172
rect 310888 60036 310940 60042
rect 310888 59978 310940 59984
rect 310900 55214 310928 59978
rect 310888 55208 310940 55214
rect 310888 55150 310940 55156
rect 311072 55208 311124 55214
rect 311072 55150 311124 55156
rect 311084 45665 311112 55150
rect 310886 45656 310942 45665
rect 310886 45591 310942 45600
rect 311070 45656 311126 45665
rect 311070 45591 311126 45600
rect 310900 45558 310928 45591
rect 310888 45552 310940 45558
rect 310888 45494 310940 45500
rect 311072 45552 311124 45558
rect 311072 45494 311124 45500
rect 311084 35902 311112 45494
rect 311072 35896 311124 35902
rect 311072 35838 311124 35844
rect 310888 26308 310940 26314
rect 310888 26250 310940 26256
rect 310900 24834 310928 26250
rect 310808 24806 310928 24834
rect 310808 22166 310836 24806
rect 310796 22160 310848 22166
rect 310796 22102 310848 22108
rect 310888 15224 310940 15230
rect 310888 15166 310940 15172
rect 310900 11286 310928 15166
rect 310888 11280 310940 11286
rect 310888 11222 310940 11228
rect 312004 9586 312032 340054
rect 312544 337272 312596 337278
rect 312544 337214 312596 337220
rect 311992 9580 312044 9586
rect 311992 9522 312044 9528
rect 310612 9512 310664 9518
rect 310612 9454 310664 9460
rect 310520 5636 310572 5642
rect 310520 5578 310572 5584
rect 312082 4992 312138 5001
rect 312082 4927 312138 4936
rect 312096 4214 312124 4927
rect 312084 4208 312136 4214
rect 312084 4150 312136 4156
rect 312176 4208 312228 4214
rect 312176 4150 312228 4156
rect 309784 4072 309836 4078
rect 309784 4014 309836 4020
rect 310980 3392 311032 3398
rect 310980 3334 311032 3340
rect 309784 3188 309836 3194
rect 309784 3130 309836 3136
rect 309796 480 309824 3130
rect 310992 480 311020 3334
rect 312188 480 312216 4150
rect 312556 3058 312584 337214
rect 312740 337142 312768 340068
rect 312728 337136 312780 337142
rect 312728 337078 312780 337084
rect 313292 5574 313320 340068
rect 313384 340054 313766 340082
rect 313384 9654 313412 340054
rect 314212 337210 314240 340068
rect 314778 340054 314884 340082
rect 314660 338088 314712 338094
rect 314660 338030 314712 338036
rect 314200 337204 314252 337210
rect 314200 337146 314252 337152
rect 313372 9648 313424 9654
rect 313372 9590 313424 9596
rect 313280 5568 313332 5574
rect 313280 5510 313332 5516
rect 314672 4865 314700 338030
rect 314856 12986 314884 340054
rect 314948 340054 315238 340082
rect 315408 340054 315698 340082
rect 314844 12980 314896 12986
rect 314844 12922 314896 12928
rect 314948 8906 314976 340054
rect 315408 338094 315436 340054
rect 316132 338156 316184 338162
rect 316132 338098 316184 338104
rect 315396 338088 315448 338094
rect 315396 338030 315448 338036
rect 316040 337340 316092 337346
rect 316040 337282 316092 337288
rect 315946 87408 316002 87417
rect 315946 87343 316002 87352
rect 315960 87145 315988 87343
rect 315946 87136 316002 87145
rect 315946 87071 316002 87080
rect 315948 40180 316000 40186
rect 315948 40122 316000 40128
rect 315960 40089 315988 40122
rect 315946 40080 316002 40089
rect 315946 40015 316002 40024
rect 315946 28928 316002 28937
rect 315946 28863 315948 28872
rect 316000 28863 316002 28872
rect 315948 28834 316000 28840
rect 314936 8900 314988 8906
rect 314936 8842 314988 8848
rect 315948 5024 316000 5030
rect 315946 4992 315948 5001
rect 316000 4992 316002 5001
rect 315946 4927 316002 4936
rect 314658 4856 314714 4865
rect 314658 4791 314714 4800
rect 316052 4758 316080 337282
rect 316144 8838 316172 338098
rect 316236 12918 316264 340068
rect 316328 340054 316710 340082
rect 316880 340054 317170 340082
rect 317616 340054 317722 340082
rect 317892 340054 318182 340082
rect 318352 340054 318642 340082
rect 318996 340054 319194 340082
rect 319272 340054 319654 340082
rect 319824 340054 320114 340082
rect 320284 340054 320666 340082
rect 320744 340054 321126 340082
rect 316328 338162 316356 340054
rect 316316 338156 316368 338162
rect 316316 338098 316368 338104
rect 316880 337346 316908 340054
rect 317328 337748 317380 337754
rect 317328 337690 317380 337696
rect 317340 337657 317368 337690
rect 317326 337648 317382 337657
rect 317326 337583 317382 337592
rect 316868 337340 316920 337346
rect 316868 337282 316920 337288
rect 317420 337340 317472 337346
rect 317420 337282 317472 337288
rect 316684 337136 316736 337142
rect 316684 337078 316736 337084
rect 316224 12912 316276 12918
rect 316224 12854 316276 12860
rect 316132 8832 316184 8838
rect 316132 8774 316184 8780
rect 316040 4752 316092 4758
rect 316040 4694 316092 4700
rect 314568 4072 314620 4078
rect 314568 4014 314620 4020
rect 313372 4004 313424 4010
rect 313372 3946 313424 3952
rect 312544 3052 312596 3058
rect 312544 2994 312596 3000
rect 313384 480 313412 3946
rect 314580 480 314608 4014
rect 316696 3262 316724 337078
rect 317326 29336 317382 29345
rect 317326 29271 317382 29280
rect 317340 28937 317368 29271
rect 317326 28928 317382 28937
rect 317326 28863 317382 28872
rect 317432 4690 317460 337282
rect 317512 306400 317564 306406
rect 317512 306342 317564 306348
rect 317524 219434 317552 306342
rect 317512 219428 317564 219434
rect 317512 219370 317564 219376
rect 317512 209840 317564 209846
rect 317512 209782 317564 209788
rect 317524 200122 317552 209782
rect 317512 200116 317564 200122
rect 317512 200058 317564 200064
rect 317512 190528 317564 190534
rect 317512 190470 317564 190476
rect 317524 180810 317552 190470
rect 317512 180804 317564 180810
rect 317512 180746 317564 180752
rect 317512 142180 317564 142186
rect 317512 142122 317564 142128
rect 317524 137970 317552 142122
rect 317512 137964 317564 137970
rect 317512 137906 317564 137912
rect 317512 55276 317564 55282
rect 317512 55218 317564 55224
rect 317524 45558 317552 55218
rect 317512 45552 317564 45558
rect 317512 45494 317564 45500
rect 317512 31816 317564 31822
rect 317512 31758 317564 31764
rect 317524 8770 317552 31758
rect 317616 12850 317644 340054
rect 317892 337770 317920 340054
rect 317708 337742 317920 337770
rect 317708 306406 317736 337742
rect 318352 337346 318380 340054
rect 318800 338156 318852 338162
rect 318800 338098 318852 338104
rect 318340 337340 318392 337346
rect 318340 337282 318392 337288
rect 317696 306400 317748 306406
rect 317696 306342 317748 306348
rect 317696 219428 317748 219434
rect 317696 219370 317748 219376
rect 317708 209846 317736 219370
rect 317696 209840 317748 209846
rect 317696 209782 317748 209788
rect 317696 200116 317748 200122
rect 317696 200058 317748 200064
rect 317708 190534 317736 200058
rect 317696 190528 317748 190534
rect 317696 190470 317748 190476
rect 317696 180804 317748 180810
rect 317696 180746 317748 180752
rect 317708 142186 317736 180746
rect 317696 142180 317748 142186
rect 317696 142122 317748 142128
rect 317788 137964 317840 137970
rect 317788 137906 317840 137912
rect 317800 128330 317828 137906
rect 317708 128302 317828 128330
rect 317708 125594 317736 128302
rect 317696 125588 317748 125594
rect 317696 125530 317748 125536
rect 317972 125588 318024 125594
rect 317972 125530 318024 125536
rect 317984 115977 318012 125530
rect 317786 115968 317842 115977
rect 317786 115903 317842 115912
rect 317970 115968 318026 115977
rect 317970 115903 318026 115912
rect 317800 104922 317828 115903
rect 317788 104916 317840 104922
rect 317788 104858 317840 104864
rect 317972 104916 318024 104922
rect 317972 104858 318024 104864
rect 317984 93974 318012 104858
rect 317972 93968 318024 93974
rect 317972 93910 318024 93916
rect 317696 93900 317748 93906
rect 317696 93842 317748 93848
rect 317708 88398 317736 93842
rect 317696 88392 317748 88398
rect 317696 88334 317748 88340
rect 317696 75948 317748 75954
rect 317696 75890 317748 75896
rect 317708 55282 317736 75890
rect 317696 55276 317748 55282
rect 317696 55218 317748 55224
rect 317696 45552 317748 45558
rect 317696 45494 317748 45500
rect 317708 31822 317736 45494
rect 317696 31816 317748 31822
rect 317696 31758 317748 31764
rect 317604 12844 317656 12850
rect 317604 12786 317656 12792
rect 317512 8764 317564 8770
rect 317512 8706 317564 8712
rect 318708 4956 318760 4962
rect 318708 4898 318760 4904
rect 317420 4684 317472 4690
rect 317420 4626 317472 4632
rect 318720 3466 318748 4898
rect 318812 4622 318840 338098
rect 318892 337340 318944 337346
rect 318892 337282 318944 337288
rect 318904 8702 318932 337282
rect 318996 12782 319024 340054
rect 319272 337346 319300 340054
rect 319824 338162 319852 340054
rect 319812 338156 319864 338162
rect 319812 338098 319864 338104
rect 319260 337340 319312 337346
rect 319260 337282 319312 337288
rect 320180 337340 320232 337346
rect 320180 337282 320232 337288
rect 319444 337000 319496 337006
rect 319444 336942 319496 336948
rect 318984 12776 319036 12782
rect 318984 12718 319036 12724
rect 318892 8696 318944 8702
rect 318892 8638 318944 8644
rect 318800 4616 318852 4622
rect 318800 4558 318852 4564
rect 318708 3460 318760 3466
rect 318708 3402 318760 3408
rect 316684 3256 316736 3262
rect 316684 3198 316736 3204
rect 318064 3256 318116 3262
rect 318064 3198 318116 3204
rect 315764 3052 315816 3058
rect 315764 2994 315816 3000
rect 315776 480 315804 2994
rect 316960 2984 317012 2990
rect 316960 2926 317012 2932
rect 316972 480 317000 2926
rect 318076 480 318104 3198
rect 319456 3126 319484 336942
rect 320192 8634 320220 337282
rect 320284 12714 320312 340054
rect 320744 337346 320772 340054
rect 320732 337340 320784 337346
rect 320732 337282 320784 337288
rect 321468 337204 321520 337210
rect 321468 337146 321520 337152
rect 320824 16720 320876 16726
rect 320822 16688 320824 16697
rect 320876 16688 320878 16697
rect 320822 16623 320878 16632
rect 320272 12708 320324 12714
rect 320272 12650 320324 12656
rect 320180 8628 320232 8634
rect 320180 8570 320232 8576
rect 320364 4548 320416 4554
rect 320364 4490 320416 4496
rect 320376 3534 320404 4490
rect 321480 3534 321508 337146
rect 321572 4622 321600 340068
rect 321756 340054 322138 340082
rect 322216 340054 322598 340082
rect 322952 340054 323058 340082
rect 323136 340054 323518 340082
rect 323688 340054 324070 340082
rect 324332 340054 324530 340082
rect 324700 340054 324990 340082
rect 325160 340054 325542 340082
rect 325712 340054 326002 340082
rect 326080 340054 326462 340082
rect 321652 335640 321704 335646
rect 321652 335582 321704 335588
rect 321664 8566 321692 335582
rect 321756 12646 321784 340054
rect 322216 335646 322244 340054
rect 322204 335640 322256 335646
rect 322204 335582 322256 335588
rect 322202 29336 322258 29345
rect 322202 29271 322258 29280
rect 322216 29073 322244 29271
rect 322202 29064 322258 29073
rect 322202 28999 322258 29008
rect 321744 12640 321796 12646
rect 321744 12582 321796 12588
rect 321652 8560 321704 8566
rect 321652 8502 321704 8508
rect 322952 4690 322980 340054
rect 323136 12578 323164 340054
rect 323688 328506 323716 340054
rect 323308 328500 323360 328506
rect 323308 328442 323360 328448
rect 323676 328500 323728 328506
rect 323676 328442 323728 328448
rect 323320 311982 323348 328442
rect 323308 311976 323360 311982
rect 323308 311918 323360 311924
rect 323216 311908 323268 311914
rect 323216 311850 323268 311856
rect 323228 304314 323256 311850
rect 323228 304286 323440 304314
rect 323412 302138 323440 304286
rect 323320 302110 323440 302138
rect 323320 299470 323348 302110
rect 323308 299464 323360 299470
rect 323308 299406 323360 299412
rect 323492 288516 323544 288522
rect 323492 288458 323544 288464
rect 323504 288425 323532 288458
rect 323214 288416 323270 288425
rect 323214 288351 323270 288360
rect 323490 288416 323546 288425
rect 323490 288351 323546 288360
rect 323228 278798 323256 288351
rect 323216 278792 323268 278798
rect 323216 278734 323268 278740
rect 323308 278792 323360 278798
rect 323308 278734 323360 278740
rect 323320 269113 323348 278734
rect 323306 269104 323362 269113
rect 323306 269039 323362 269048
rect 323398 268968 323454 268977
rect 323398 268903 323454 268912
rect 323412 254046 323440 268903
rect 323400 254040 323452 254046
rect 323400 253982 323452 253988
rect 323308 253904 323360 253910
rect 323308 253846 323360 253852
rect 323320 241534 323348 253846
rect 323308 241528 323360 241534
rect 323308 241470 323360 241476
rect 323400 241528 323452 241534
rect 323400 241470 323452 241476
rect 323412 234734 323440 241470
rect 323400 234728 323452 234734
rect 323400 234670 323452 234676
rect 323400 231804 323452 231810
rect 323400 231746 323452 231752
rect 323412 217546 323440 231746
rect 323412 217518 323532 217546
rect 323504 211177 323532 217518
rect 323306 211168 323362 211177
rect 323306 211103 323362 211112
rect 323490 211168 323546 211177
rect 323490 211103 323546 211112
rect 323320 205698 323348 211103
rect 323308 205692 323360 205698
rect 323308 205634 323360 205640
rect 323400 205556 323452 205562
rect 323400 205498 323452 205504
rect 323412 198098 323440 205498
rect 323412 198070 323532 198098
rect 323504 193254 323532 198070
rect 323308 193248 323360 193254
rect 323306 193216 323308 193225
rect 323492 193248 323544 193254
rect 323360 193216 323362 193225
rect 323306 193151 323362 193160
rect 323490 193216 323492 193225
rect 323544 193216 323546 193225
rect 323490 193151 323546 193160
rect 323504 186266 323532 193151
rect 323412 186238 323532 186266
rect 323412 178786 323440 186238
rect 323412 178758 323532 178786
rect 323504 173942 323532 178758
rect 323308 173936 323360 173942
rect 323308 173878 323360 173884
rect 323492 173936 323544 173942
rect 323492 173878 323544 173884
rect 323320 169402 323348 173878
rect 323320 169374 323440 169402
rect 323412 157434 323440 169374
rect 324226 157448 324282 157457
rect 323412 157406 323532 157434
rect 323504 155666 323532 157406
rect 324226 157383 324282 157392
rect 324240 157185 324268 157383
rect 324226 157176 324282 157185
rect 324226 157111 324282 157120
rect 323412 155638 323532 155666
rect 323412 144906 323440 155638
rect 323308 144900 323360 144906
rect 323308 144842 323360 144848
rect 323400 144900 323452 144906
rect 323400 144842 323452 144848
rect 323320 143546 323348 144842
rect 323308 143540 323360 143546
rect 323308 143482 323360 143488
rect 323308 133952 323360 133958
rect 323308 133894 323360 133900
rect 323320 128058 323348 133894
rect 323320 128030 323440 128058
rect 323412 116113 323440 128030
rect 323398 116104 323454 116113
rect 323398 116039 323454 116048
rect 323306 115968 323362 115977
rect 323306 115903 323362 115912
rect 323320 106298 323348 115903
rect 323320 106270 323440 106298
rect 323412 99634 323440 106270
rect 323228 99606 323440 99634
rect 323228 96608 323256 99606
rect 323228 96580 323440 96608
rect 323412 86970 323440 96580
rect 323308 86964 323360 86970
rect 323308 86906 323360 86912
rect 323400 86964 323452 86970
rect 323400 86906 323452 86912
rect 323320 67726 323348 86906
rect 323308 67720 323360 67726
rect 323308 67662 323360 67668
rect 323400 67652 323452 67658
rect 323400 67594 323452 67600
rect 323412 66230 323440 67594
rect 323400 66224 323452 66230
rect 323400 66166 323452 66172
rect 323308 48340 323360 48346
rect 323308 48282 323360 48288
rect 323320 46918 323348 48282
rect 323308 46912 323360 46918
rect 323308 46854 323360 46860
rect 323400 37324 323452 37330
rect 323400 37266 323452 37272
rect 323412 28966 323440 37266
rect 323308 28960 323360 28966
rect 323308 28902 323360 28908
rect 323400 28960 323452 28966
rect 323400 28902 323452 28908
rect 323124 12572 323176 12578
rect 323124 12514 323176 12520
rect 323320 8498 323348 28902
rect 323308 8492 323360 8498
rect 323308 8434 323360 8440
rect 324332 4826 324360 340054
rect 324700 335730 324728 340054
rect 324424 335702 324728 335730
rect 324424 7614 324452 335702
rect 325160 328506 325188 340054
rect 324688 328500 324740 328506
rect 324688 328442 324740 328448
rect 325148 328500 325200 328506
rect 325148 328442 325200 328448
rect 324700 311930 324728 328442
rect 324608 311902 324728 311930
rect 324608 304314 324636 311902
rect 325608 307760 325660 307766
rect 325608 307702 325660 307708
rect 324516 304286 324636 304314
rect 324516 302138 324544 304286
rect 324516 302110 324728 302138
rect 324700 299470 324728 302110
rect 324688 299464 324740 299470
rect 324688 299406 324740 299412
rect 325620 298217 325648 307702
rect 325606 298208 325662 298217
rect 325606 298143 325662 298152
rect 324688 289876 324740 289882
rect 324688 289818 324740 289824
rect 324700 285002 324728 289818
rect 324700 284974 324820 285002
rect 324792 270570 324820 284974
rect 324688 270564 324740 270570
rect 324688 270506 324740 270512
rect 324780 270564 324832 270570
rect 324780 270506 324832 270512
rect 324700 269113 324728 270506
rect 324686 269104 324742 269113
rect 324686 269039 324742 269048
rect 324870 269104 324926 269113
rect 324870 269039 324926 269048
rect 324884 260658 324912 269039
rect 324700 260630 324912 260658
rect 324700 241602 324728 260630
rect 324688 241596 324740 241602
rect 324688 241538 324740 241544
rect 324596 241528 324648 241534
rect 324596 241470 324648 241476
rect 324608 240106 324636 241470
rect 324596 240100 324648 240106
rect 324596 240042 324648 240048
rect 324780 231804 324832 231810
rect 324780 231746 324832 231752
rect 324792 212566 324820 231746
rect 324688 212560 324740 212566
rect 324688 212502 324740 212508
rect 324780 212560 324832 212566
rect 324780 212502 324832 212508
rect 324700 202910 324728 212502
rect 324596 202904 324648 202910
rect 324596 202846 324648 202852
rect 324688 202904 324740 202910
rect 324688 202846 324740 202852
rect 324608 193254 324636 202846
rect 324596 193248 324648 193254
rect 324688 193248 324740 193254
rect 324648 193196 324688 193202
rect 324596 193190 324740 193196
rect 324608 193174 324728 193190
rect 324608 183569 324636 193174
rect 324594 183560 324650 183569
rect 324594 183495 324650 183504
rect 324778 183560 324834 183569
rect 324778 183495 324834 183504
rect 324792 173942 324820 183495
rect 324688 173936 324740 173942
rect 324688 173878 324740 173884
rect 324780 173936 324832 173942
rect 324780 173878 324832 173884
rect 324700 164234 324728 173878
rect 324608 164206 324728 164234
rect 324608 157400 324636 164206
rect 324608 157372 324820 157400
rect 324792 154544 324820 157372
rect 324608 154516 324820 154544
rect 324608 144945 324636 154516
rect 324594 144936 324650 144945
rect 324594 144871 324650 144880
rect 324594 144800 324650 144809
rect 324594 144735 324650 144744
rect 324608 143546 324636 144735
rect 324596 143540 324648 143546
rect 324596 143482 324648 143488
rect 324688 132524 324740 132530
rect 324688 132466 324740 132472
rect 324700 122806 324728 132466
rect 324688 122800 324740 122806
rect 324688 122742 324740 122748
rect 324688 113212 324740 113218
rect 324688 113154 324740 113160
rect 324700 106264 324728 113154
rect 324608 106236 324728 106264
rect 324608 104854 324636 106236
rect 324596 104848 324648 104854
rect 324596 104790 324648 104796
rect 324688 104848 324740 104854
rect 324688 104790 324740 104796
rect 324700 103494 324728 104790
rect 324688 103488 324740 103494
rect 324688 103430 324740 103436
rect 324596 93900 324648 93906
rect 324596 93842 324648 93848
rect 324608 86970 324636 93842
rect 324596 86964 324648 86970
rect 324596 86906 324648 86912
rect 324688 86896 324740 86902
rect 324688 86838 324740 86844
rect 324700 85542 324728 86838
rect 324688 85536 324740 85542
rect 324688 85478 324740 85484
rect 324688 76016 324740 76022
rect 324688 75958 324740 75964
rect 324700 75886 324728 75958
rect 324688 75880 324740 75886
rect 324688 75822 324740 75828
rect 324596 66360 324648 66366
rect 324596 66302 324648 66308
rect 324608 66230 324636 66302
rect 324596 66224 324648 66230
rect 324596 66166 324648 66172
rect 324688 61396 324740 61402
rect 324688 61338 324740 61344
rect 324700 56658 324728 61338
rect 324700 56630 324820 56658
rect 324792 56574 324820 56630
rect 324780 56568 324832 56574
rect 324780 56510 324832 56516
rect 324596 46980 324648 46986
rect 324596 46922 324648 46928
rect 324608 46866 324636 46922
rect 324608 46838 324728 46866
rect 324700 28966 324728 46838
rect 324596 28960 324648 28966
rect 324596 28902 324648 28908
rect 324688 28960 324740 28966
rect 324688 28902 324740 28908
rect 324608 8430 324636 28902
rect 325606 16824 325662 16833
rect 325606 16759 325662 16768
rect 325620 16726 325648 16759
rect 325608 16720 325660 16726
rect 325608 16662 325660 16668
rect 324596 8424 324648 8430
rect 324596 8366 324648 8372
rect 324412 7608 324464 7614
rect 324412 7550 324464 7556
rect 325608 5024 325660 5030
rect 325608 4966 325660 4972
rect 324320 4820 324372 4826
rect 324320 4762 324372 4768
rect 324228 4752 324280 4758
rect 324228 4694 324280 4700
rect 322940 4684 322992 4690
rect 322940 4626 322992 4632
rect 321560 4616 321612 4622
rect 321560 4558 321612 4564
rect 322572 4480 322624 4486
rect 322572 4422 322624 4428
rect 322584 3670 322612 4422
rect 322572 3664 322624 3670
rect 322572 3606 322624 3612
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 320364 3528 320416 3534
rect 320364 3470 320416 3476
rect 320456 3528 320508 3534
rect 320456 3470 320508 3476
rect 321468 3528 321520 3534
rect 321468 3470 321520 3476
rect 319444 3120 319496 3126
rect 319444 3062 319496 3068
rect 319260 2916 319312 2922
rect 319260 2858 319312 2864
rect 319272 480 319300 2858
rect 320468 480 320496 3470
rect 321652 3460 321704 3466
rect 321652 3402 321704 3408
rect 321664 480 321692 3402
rect 322860 480 322888 3538
rect 324044 3528 324096 3534
rect 324044 3470 324096 3476
rect 324056 480 324084 3470
rect 324240 3058 324268 4694
rect 325620 3942 325648 4966
rect 325712 4894 325740 340054
rect 326080 335594 326108 340054
rect 325804 335566 326108 335594
rect 325804 7682 325832 335566
rect 326540 333334 326568 340190
rect 327092 340054 327474 340082
rect 327644 340054 327934 340082
rect 328486 340054 328684 340082
rect 325976 333328 326028 333334
rect 325976 333270 326028 333276
rect 326528 333328 326580 333334
rect 326528 333270 326580 333276
rect 325988 307766 326016 333270
rect 325976 307760 326028 307766
rect 325976 307702 326028 307708
rect 325882 298174 325938 298183
rect 325882 298109 325938 298118
rect 325896 296721 325924 298109
rect 325882 296712 325938 296721
rect 325882 296647 325938 296656
rect 326066 296712 326122 296721
rect 326066 296647 326122 296656
rect 326080 288386 326108 296647
rect 325884 288380 325936 288386
rect 325884 288322 325936 288328
rect 326068 288380 326120 288386
rect 326068 288322 326120 288328
rect 325896 280226 325924 288322
rect 325884 280220 325936 280226
rect 325884 280162 325936 280168
rect 325884 278792 325936 278798
rect 325884 278734 325936 278740
rect 325896 270570 325924 278734
rect 325884 270564 325936 270570
rect 325884 270506 325936 270512
rect 325976 270564 326028 270570
rect 325976 270506 326028 270512
rect 325988 260982 326016 270506
rect 325976 260976 326028 260982
rect 325976 260918 326028 260924
rect 325976 260772 326028 260778
rect 325976 260714 326028 260720
rect 325988 241602 326016 260714
rect 325976 241596 326028 241602
rect 325976 241538 326028 241544
rect 325884 241528 325936 241534
rect 325884 241470 325936 241476
rect 325896 240145 325924 241470
rect 325882 240136 325938 240145
rect 325882 240071 325938 240080
rect 326158 240136 326214 240145
rect 326158 240071 326214 240080
rect 326172 230518 326200 240071
rect 325976 230512 326028 230518
rect 325976 230454 326028 230460
rect 326160 230512 326212 230518
rect 326160 230454 326212 230460
rect 325988 227202 326016 230454
rect 325988 227174 326108 227202
rect 326080 222222 326108 227174
rect 325884 222216 325936 222222
rect 325884 222158 325936 222164
rect 326068 222216 326120 222222
rect 326068 222158 326120 222164
rect 325896 212566 325924 222158
rect 325884 212560 325936 212566
rect 325884 212502 325936 212508
rect 325976 212560 326028 212566
rect 325976 212502 326028 212508
rect 325988 202910 326016 212502
rect 325884 202904 325936 202910
rect 325884 202846 325936 202852
rect 325976 202904 326028 202910
rect 325976 202846 326028 202852
rect 325896 193254 325924 202846
rect 325884 193248 325936 193254
rect 325884 193190 325936 193196
rect 325976 193248 326028 193254
rect 325976 193190 326028 193196
rect 325988 188442 326016 193190
rect 325896 188414 326016 188442
rect 325896 173942 325924 188414
rect 325884 173936 325936 173942
rect 325884 173878 325936 173884
rect 325976 173936 326028 173942
rect 325976 173878 326028 173884
rect 325988 164234 326016 173878
rect 325896 164206 326016 164234
rect 325896 157418 325924 164206
rect 325884 157412 325936 157418
rect 325884 157354 325936 157360
rect 325976 157208 326028 157214
rect 325976 157150 326028 157156
rect 325988 149818 326016 157150
rect 325988 149790 326108 149818
rect 326080 144945 326108 149790
rect 325882 144936 325938 144945
rect 325882 144871 325884 144880
rect 325936 144871 325938 144880
rect 326066 144936 326122 144945
rect 326066 144871 326068 144880
rect 325884 144842 325936 144848
rect 326120 144871 326122 144880
rect 326068 144842 326120 144848
rect 326080 137714 326108 144842
rect 325988 137686 326108 137714
rect 325988 128450 326016 137686
rect 325976 128444 326028 128450
rect 325976 128386 326028 128392
rect 325884 128308 325936 128314
rect 325884 128250 325936 128256
rect 325896 125594 325924 128250
rect 325884 125588 325936 125594
rect 325884 125530 325936 125536
rect 326068 125588 326120 125594
rect 326068 125530 326120 125536
rect 326080 118402 326108 125530
rect 325988 118374 326108 118402
rect 325988 106350 326016 118374
rect 325976 106344 326028 106350
rect 325976 106286 326028 106292
rect 325976 104916 326028 104922
rect 325976 104858 326028 104864
rect 325988 100042 326016 104858
rect 325896 100014 326016 100042
rect 325896 86970 325924 100014
rect 325884 86964 325936 86970
rect 325884 86906 325936 86912
rect 325976 86896 326028 86902
rect 325976 86838 326028 86844
rect 325988 67674 326016 86838
rect 325896 67646 326016 67674
rect 325896 61418 325924 67646
rect 325896 61390 326108 61418
rect 326080 29034 326108 61390
rect 325976 29028 326028 29034
rect 325976 28970 326028 28976
rect 326068 29028 326120 29034
rect 326068 28970 326120 28976
rect 325988 19310 326016 28970
rect 325976 19304 326028 19310
rect 325976 19246 326028 19252
rect 325976 19168 326028 19174
rect 325976 19110 326028 19116
rect 325988 8974 326016 19110
rect 325976 8968 326028 8974
rect 325976 8910 326028 8916
rect 325792 7676 325844 7682
rect 325792 7618 325844 7624
rect 327092 5098 327120 340054
rect 327644 336734 327672 340054
rect 327724 336864 327776 336870
rect 327724 336806 327776 336812
rect 327632 336728 327684 336734
rect 327632 336670 327684 336676
rect 327264 327140 327316 327146
rect 327264 327082 327316 327088
rect 327276 309058 327304 327082
rect 327264 309052 327316 309058
rect 327264 308994 327316 309000
rect 327356 309052 327408 309058
rect 327356 308994 327408 309000
rect 327368 302190 327396 308994
rect 327356 302184 327408 302190
rect 327356 302126 327408 302132
rect 327264 298172 327316 298178
rect 327264 298114 327316 298120
rect 327276 289814 327304 298114
rect 327264 289808 327316 289814
rect 327264 289750 327316 289756
rect 327356 289740 327408 289746
rect 327356 289682 327408 289688
rect 327368 273850 327396 289682
rect 327276 273822 327396 273850
rect 327276 259622 327304 273822
rect 327264 259616 327316 259622
rect 327264 259558 327316 259564
rect 327264 259412 327316 259418
rect 327264 259354 327316 259360
rect 327276 253978 327304 259354
rect 327264 253972 327316 253978
rect 327264 253914 327316 253920
rect 327172 240236 327224 240242
rect 327172 240178 327224 240184
rect 327184 240106 327212 240178
rect 327172 240100 327224 240106
rect 327172 240042 327224 240048
rect 327172 230580 327224 230586
rect 327172 230522 327224 230528
rect 327184 230489 327212 230522
rect 327170 230480 327226 230489
rect 327170 230415 327226 230424
rect 327538 230480 327594 230489
rect 327538 230415 327594 230424
rect 327552 220862 327580 230415
rect 327356 220856 327408 220862
rect 327356 220798 327408 220804
rect 327540 220856 327592 220862
rect 327540 220798 327592 220804
rect 327368 217274 327396 220798
rect 327276 217246 327396 217274
rect 327276 212537 327304 217246
rect 327262 212528 327318 212537
rect 327262 212463 327318 212472
rect 327354 212392 327410 212401
rect 327354 212327 327410 212336
rect 327368 197962 327396 212327
rect 327276 197934 327396 197962
rect 327276 186454 327304 197934
rect 327264 186448 327316 186454
rect 327264 186390 327316 186396
rect 327172 186312 327224 186318
rect 327172 186254 327224 186260
rect 327184 173942 327212 186254
rect 327172 173936 327224 173942
rect 327172 173878 327224 173884
rect 327264 173936 327316 173942
rect 327264 173878 327316 173884
rect 327276 164234 327304 173878
rect 327184 164206 327304 164234
rect 327184 157418 327212 164206
rect 327172 157412 327224 157418
rect 327172 157354 327224 157360
rect 327264 157276 327316 157282
rect 327264 157218 327316 157224
rect 327276 145081 327304 157218
rect 327262 145072 327318 145081
rect 327262 145007 327318 145016
rect 327170 144936 327226 144945
rect 327170 144871 327172 144880
rect 327224 144871 327226 144880
rect 327356 144900 327408 144906
rect 327172 144842 327224 144848
rect 327356 144842 327408 144848
rect 327368 137850 327396 144842
rect 327276 137822 327396 137850
rect 327276 128450 327304 137822
rect 327264 128444 327316 128450
rect 327264 128386 327316 128392
rect 327172 128308 327224 128314
rect 327172 128250 327224 128256
rect 327184 125594 327212 128250
rect 327172 125588 327224 125594
rect 327172 125530 327224 125536
rect 327356 125588 327408 125594
rect 327356 125530 327408 125536
rect 327368 118522 327396 125530
rect 327264 118516 327316 118522
rect 327264 118458 327316 118464
rect 327356 118516 327408 118522
rect 327356 118458 327408 118464
rect 327276 114510 327304 118458
rect 327264 114504 327316 114510
rect 327264 114446 327316 114452
rect 327172 104916 327224 104922
rect 327172 104858 327224 104864
rect 327184 86970 327212 104858
rect 327172 86964 327224 86970
rect 327172 86906 327224 86912
rect 327264 86964 327316 86970
rect 327264 86906 327316 86912
rect 327276 77466 327304 86906
rect 327276 77438 327396 77466
rect 327368 74610 327396 77438
rect 327276 74582 327396 74610
rect 327276 66298 327304 74582
rect 327264 66292 327316 66298
rect 327264 66234 327316 66240
rect 327356 66156 327408 66162
rect 327356 66098 327408 66104
rect 327368 60602 327396 66098
rect 327276 60574 327396 60602
rect 327276 46918 327304 60574
rect 327264 46912 327316 46918
rect 327264 46854 327316 46860
rect 327264 37324 327316 37330
rect 327264 37266 327316 37272
rect 327276 31822 327304 37266
rect 327264 31816 327316 31822
rect 327264 31758 327316 31764
rect 327264 31612 327316 31618
rect 327264 31554 327316 31560
rect 327276 19310 327304 31554
rect 327264 19304 327316 19310
rect 327264 19246 327316 19252
rect 327264 19168 327316 19174
rect 327264 19110 327316 19116
rect 327276 7002 327304 19110
rect 327264 6996 327316 7002
rect 327264 6938 327316 6944
rect 327080 5092 327132 5098
rect 327080 5034 327132 5040
rect 325700 4888 325752 4894
rect 325700 4830 325752 4836
rect 327080 4888 327132 4894
rect 327080 4830 327132 4836
rect 326528 4684 326580 4690
rect 326528 4626 326580 4632
rect 325608 3936 325660 3942
rect 325608 3878 325660 3884
rect 326436 3732 326488 3738
rect 326436 3674 326488 3680
rect 325240 3664 325292 3670
rect 325240 3606 325292 3612
rect 324228 3052 324280 3058
rect 324228 2994 324280 3000
rect 325252 480 325280 3606
rect 326448 480 326476 3674
rect 326540 2922 326568 4626
rect 327092 3602 327120 4830
rect 327080 3596 327132 3602
rect 327080 3538 327132 3544
rect 327736 3126 327764 336806
rect 328552 331356 328604 331362
rect 328552 331298 328604 331304
rect 328458 87272 328514 87281
rect 328458 87207 328514 87216
rect 328366 87136 328422 87145
rect 328472 87122 328500 87207
rect 328422 87094 328500 87122
rect 328366 87071 328422 87080
rect 328564 7750 328592 331298
rect 328656 9042 328684 340054
rect 328748 340054 328946 340082
rect 329024 340054 329406 340082
rect 329958 340054 330064 340082
rect 328644 9036 328696 9042
rect 328644 8978 328696 8984
rect 328552 7744 328604 7750
rect 328552 7686 328604 7692
rect 328748 4962 328776 340054
rect 329024 331362 329052 340054
rect 329840 335640 329892 335646
rect 329840 335582 329892 335588
rect 329012 331356 329064 331362
rect 329012 331298 329064 331304
rect 328920 76152 328972 76158
rect 328920 76094 328972 76100
rect 328932 75993 328960 76094
rect 328918 75984 328974 75993
rect 328918 75919 328974 75928
rect 329852 5098 329880 335582
rect 329932 297764 329984 297770
rect 329932 297706 329984 297712
rect 329944 288386 329972 297706
rect 329932 288380 329984 288386
rect 329932 288322 329984 288328
rect 329932 113144 329984 113150
rect 329932 113086 329984 113092
rect 329944 103601 329972 113086
rect 329930 103592 329986 103601
rect 329930 103527 329986 103536
rect 330036 9110 330064 340054
rect 330128 340054 330418 340082
rect 330588 340054 330878 340082
rect 331324 340054 331430 340082
rect 331508 340054 331890 340082
rect 331968 340054 332350 340082
rect 332796 340054 332902 340082
rect 333072 340054 333362 340082
rect 333440 340054 333822 340082
rect 334176 340054 334374 340082
rect 334544 340054 334834 340082
rect 334912 340054 335294 340082
rect 335464 340054 335846 340082
rect 336016 340054 336306 340082
rect 330128 335646 330156 340054
rect 330588 338042 330616 340054
rect 330496 338014 330616 338042
rect 330116 335640 330168 335646
rect 330116 335582 330168 335588
rect 330496 327214 330524 338014
rect 331324 333282 331352 340054
rect 331324 333254 331444 333282
rect 331220 332172 331272 332178
rect 331220 332114 331272 332120
rect 330484 327208 330536 327214
rect 330484 327150 330536 327156
rect 330116 327140 330168 327146
rect 330116 327082 330168 327088
rect 330128 318850 330156 327082
rect 330116 318844 330168 318850
rect 330116 318786 330168 318792
rect 330208 318708 330260 318714
rect 330208 318650 330260 318656
rect 330220 316033 330248 318650
rect 330206 316024 330262 316033
rect 330206 315959 330262 315968
rect 330390 316024 330446 316033
rect 330390 315959 330446 315968
rect 330404 297770 330432 315959
rect 330392 297764 330444 297770
rect 330392 297706 330444 297712
rect 330300 288380 330352 288386
rect 330300 288322 330352 288328
rect 330312 282826 330340 288322
rect 330128 282798 330340 282826
rect 330128 273970 330156 282798
rect 330116 273964 330168 273970
rect 330116 273906 330168 273912
rect 330116 260908 330168 260914
rect 330116 260850 330168 260856
rect 330128 258890 330156 260850
rect 330128 258862 330248 258890
rect 330220 249801 330248 258862
rect 330206 249792 330262 249801
rect 330206 249727 330262 249736
rect 330390 249792 330446 249801
rect 330390 249727 330446 249736
rect 330404 241346 330432 249727
rect 330220 241318 330432 241346
rect 330220 240122 330248 241318
rect 330220 240094 330432 240122
rect 330404 220862 330432 240094
rect 330208 220856 330260 220862
rect 330208 220798 330260 220804
rect 330392 220856 330444 220862
rect 330392 220798 330444 220804
rect 330220 212498 330248 220798
rect 330208 212492 330260 212498
rect 330208 212434 330260 212440
rect 330300 212492 330352 212498
rect 330300 212434 330352 212440
rect 330312 195922 330340 212434
rect 330220 195894 330340 195922
rect 330220 186454 330248 195894
rect 330208 186448 330260 186454
rect 330208 186390 330260 186396
rect 330208 186244 330260 186250
rect 330208 186186 330260 186192
rect 330220 183410 330248 186186
rect 330128 183382 330248 183410
rect 330128 172514 330156 183382
rect 330116 172508 330168 172514
rect 330116 172450 330168 172456
rect 330116 162988 330168 162994
rect 330116 162930 330168 162936
rect 330128 161430 330156 162930
rect 330116 161424 330168 161430
rect 330116 161366 330168 161372
rect 330116 151836 330168 151842
rect 330116 151778 330168 151784
rect 330128 147694 330156 151778
rect 330116 147688 330168 147694
rect 330116 147630 330168 147636
rect 330208 147620 330260 147626
rect 330208 147562 330260 147568
rect 330220 143546 330248 147562
rect 330208 143540 330260 143546
rect 330208 143482 330260 143488
rect 330116 137964 330168 137970
rect 330116 137906 330168 137912
rect 330128 121530 330156 137906
rect 330128 121502 330248 121530
rect 330220 113150 330248 121502
rect 330208 113144 330260 113150
rect 330208 113086 330260 113092
rect 330114 103592 330170 103601
rect 330114 103527 330170 103536
rect 330128 103494 330156 103527
rect 330116 103488 330168 103494
rect 330116 103430 330168 103436
rect 330208 103488 330260 103494
rect 330208 103430 330260 103436
rect 330220 102134 330248 103430
rect 330208 102128 330260 102134
rect 330208 102070 330260 102076
rect 330208 77308 330260 77314
rect 330208 77250 330260 77256
rect 330220 67674 330248 77250
rect 330128 67646 330248 67674
rect 330128 66230 330156 67646
rect 330116 66224 330168 66230
rect 330116 66166 330168 66172
rect 330208 56636 330260 56642
rect 330208 56578 330260 56584
rect 330220 48362 330248 56578
rect 330128 48334 330248 48362
rect 330128 46918 330156 48334
rect 330116 46912 330168 46918
rect 330116 46854 330168 46860
rect 330116 37324 330168 37330
rect 330116 37266 330168 37272
rect 330128 28937 330156 37266
rect 330114 28928 330170 28937
rect 330114 28863 330170 28872
rect 330206 28792 330262 28801
rect 330206 28727 330262 28736
rect 330024 9104 330076 9110
rect 330024 9046 330076 9052
rect 330220 7818 330248 28727
rect 330208 7812 330260 7818
rect 330208 7754 330260 7760
rect 331232 5166 331260 332114
rect 331312 331764 331364 331770
rect 331312 331706 331364 331712
rect 331324 7886 331352 331706
rect 331416 8362 331444 333254
rect 331508 332178 331536 340054
rect 331496 332172 331548 332178
rect 331496 332114 331548 332120
rect 331968 331770 331996 340054
rect 332692 335708 332744 335714
rect 332692 335650 332744 335656
rect 332600 335640 332652 335646
rect 332600 335582 332652 335588
rect 331956 331764 332008 331770
rect 331956 331706 332008 331712
rect 331862 29608 331918 29617
rect 331862 29543 331918 29552
rect 331876 29345 331904 29543
rect 331862 29336 331918 29345
rect 331862 29271 331918 29280
rect 331404 8356 331456 8362
rect 331404 8298 331456 8304
rect 331312 7880 331364 7886
rect 331312 7822 331364 7828
rect 332612 5234 332640 335582
rect 332704 7954 332732 335650
rect 332796 9178 332824 340054
rect 333072 335646 333100 340054
rect 333244 336932 333296 336938
rect 333244 336874 333296 336880
rect 333060 335640 333112 335646
rect 333060 335582 333112 335588
rect 332784 9172 332836 9178
rect 332784 9114 332836 9120
rect 332692 7948 332744 7954
rect 332692 7890 332744 7896
rect 332600 5228 332652 5234
rect 332600 5170 332652 5176
rect 331220 5160 331272 5166
rect 331220 5102 331272 5108
rect 329840 5092 329892 5098
rect 329840 5034 329892 5040
rect 328736 4956 328788 4962
rect 328736 4898 328788 4904
rect 328460 4820 328512 4826
rect 328460 4762 328512 4768
rect 328472 3738 328500 4762
rect 333256 4146 333284 336874
rect 333440 335714 333468 340054
rect 333428 335708 333480 335714
rect 333428 335650 333480 335656
rect 334072 335708 334124 335714
rect 334072 335650 334124 335656
rect 333980 335640 334032 335646
rect 333980 335582 334032 335588
rect 333886 157720 333942 157729
rect 333886 157655 333942 157664
rect 333900 157457 333928 157655
rect 333886 157448 333942 157457
rect 333886 157383 333942 157392
rect 333612 4956 333664 4962
rect 333612 4898 333664 4904
rect 332416 4140 332468 4146
rect 332416 4082 332468 4088
rect 333244 4140 333296 4146
rect 333244 4082 333296 4088
rect 328460 3732 328512 3738
rect 328460 3674 328512 3680
rect 331220 3732 331272 3738
rect 331220 3674 331272 3680
rect 327724 3120 327776 3126
rect 327724 3062 327776 3068
rect 328828 3120 328880 3126
rect 328828 3062 328880 3068
rect 327632 3052 327684 3058
rect 327632 2994 327684 3000
rect 326528 2916 326580 2922
rect 326528 2858 326580 2864
rect 327644 480 327672 2994
rect 328840 480 328868 3062
rect 330024 2848 330076 2854
rect 330024 2790 330076 2796
rect 330036 480 330064 2790
rect 331232 480 331260 3674
rect 332428 480 332456 4082
rect 333624 480 333652 4898
rect 333992 4622 334020 335582
rect 334084 8022 334112 335650
rect 334176 9246 334204 340054
rect 334544 335646 334572 340054
rect 334912 335714 334940 340054
rect 335268 337136 335320 337142
rect 335268 337078 335320 337084
rect 334900 335708 334952 335714
rect 334900 335650 334952 335656
rect 334532 335640 334584 335646
rect 334532 335582 334584 335588
rect 334164 9240 334216 9246
rect 334164 9182 334216 9188
rect 334072 8016 334124 8022
rect 334072 7958 334124 7964
rect 333980 4616 334032 4622
rect 333980 4558 334032 4564
rect 335280 4146 335308 337078
rect 335360 335640 335412 335646
rect 335360 335582 335412 335588
rect 335372 4554 335400 335582
rect 335464 6594 335492 340054
rect 336016 335646 336044 340054
rect 336096 337680 336148 337686
rect 336096 337622 336148 337628
rect 336004 335640 336056 335646
rect 336004 335582 336056 335588
rect 336108 334506 336136 337622
rect 336016 334478 336136 334506
rect 335452 6588 335504 6594
rect 335452 6530 335504 6536
rect 335360 4548 335412 4554
rect 335360 4490 335412 4496
rect 334716 4140 334768 4146
rect 334716 4082 334768 4088
rect 335268 4140 335320 4146
rect 335268 4082 335320 4088
rect 334728 480 334756 4082
rect 335544 3800 335596 3806
rect 336016 3754 336044 334478
rect 336752 333334 336780 340068
rect 336844 340054 337318 340082
rect 337396 340054 337778 340082
rect 338238 340054 338344 340082
rect 336740 333328 336792 333334
rect 336740 333270 336792 333276
rect 336844 331294 336872 340054
rect 336924 333328 336976 333334
rect 336924 333270 336976 333276
rect 336832 331288 336884 331294
rect 336832 331230 336884 331236
rect 336832 331152 336884 331158
rect 336832 331094 336884 331100
rect 336738 240136 336794 240145
rect 336738 240071 336794 240080
rect 336752 230518 336780 240071
rect 336740 230512 336792 230518
rect 336740 230454 336792 230460
rect 336740 225480 336792 225486
rect 336740 225422 336792 225428
rect 336752 212566 336780 225422
rect 336740 212560 336792 212566
rect 336740 212502 336792 212508
rect 336738 183560 336794 183569
rect 336738 183495 336794 183504
rect 336752 173942 336780 183495
rect 336740 173936 336792 173942
rect 336740 173878 336792 173884
rect 336740 125588 336792 125594
rect 336740 125530 336792 125536
rect 336752 115977 336780 125530
rect 336738 115968 336794 115977
rect 336738 115903 336794 115912
rect 336740 33856 336792 33862
rect 336740 33798 336792 33804
rect 336752 19378 336780 33798
rect 336740 19372 336792 19378
rect 336740 19314 336792 19320
rect 336646 17096 336702 17105
rect 336646 17031 336702 17040
rect 336660 16697 336688 17031
rect 336646 16688 336702 16697
rect 336646 16623 336702 16632
rect 336844 6662 336872 331094
rect 336936 280158 336964 333270
rect 337396 328506 337424 340054
rect 338120 335640 338172 335646
rect 338120 335582 338172 335588
rect 337292 328500 337344 328506
rect 337292 328442 337344 328448
rect 337384 328500 337436 328506
rect 337384 328442 337436 328448
rect 337304 321638 337332 328442
rect 337292 321632 337344 321638
rect 337292 321574 337344 321580
rect 337384 321496 337436 321502
rect 337384 321438 337436 321444
rect 337396 311914 337424 321438
rect 337200 311908 337252 311914
rect 337200 311850 337252 311856
rect 337384 311908 337436 311914
rect 337384 311850 337436 311856
rect 337212 307766 337240 311850
rect 337200 307760 337252 307766
rect 337200 307702 337252 307708
rect 337016 298240 337068 298246
rect 337016 298182 337068 298188
rect 337028 298110 337056 298182
rect 337016 298104 337068 298110
rect 337016 298046 337068 298052
rect 337200 292460 337252 292466
rect 337200 292402 337252 292408
rect 337212 288402 337240 292402
rect 337120 288374 337240 288402
rect 337120 282946 337148 288374
rect 337108 282940 337160 282946
rect 337108 282882 337160 282888
rect 336924 280152 336976 280158
rect 336924 280094 336976 280100
rect 337108 278792 337160 278798
rect 337108 278734 337160 278740
rect 337120 274009 337148 278734
rect 337106 274000 337162 274009
rect 337106 273935 337162 273944
rect 336924 270564 336976 270570
rect 336924 270506 336976 270512
rect 336936 260846 336964 270506
rect 336924 260840 336976 260846
rect 336924 260782 336976 260788
rect 336922 260672 336978 260681
rect 336922 260607 336978 260616
rect 336936 259486 336964 260607
rect 337120 259486 337148 259517
rect 336924 259480 336976 259486
rect 336924 259422 336976 259428
rect 337108 259480 337160 259486
rect 337160 259428 337332 259434
rect 337108 259422 337332 259428
rect 337120 259406 337332 259422
rect 337304 254658 337332 259406
rect 337292 254652 337344 254658
rect 337292 254594 337344 254600
rect 336924 249824 336976 249830
rect 336924 249766 336976 249772
rect 336936 240145 336964 249766
rect 337108 241596 337160 241602
rect 337108 241538 337160 241544
rect 336922 240136 336978 240145
rect 337120 240122 337148 241538
rect 337120 240094 337240 240122
rect 336922 240071 336978 240080
rect 337212 234666 337240 240094
rect 337200 234660 337252 234666
rect 337200 234602 337252 234608
rect 336924 230512 336976 230518
rect 336924 230454 336976 230460
rect 337108 230512 337160 230518
rect 337108 230454 337160 230460
rect 336936 225486 336964 230454
rect 336924 225480 336976 225486
rect 336924 225422 336976 225428
rect 337120 220833 337148 230454
rect 337106 220824 337162 220833
rect 337106 220759 337162 220768
rect 337198 220688 337254 220697
rect 337198 220623 337254 220632
rect 336924 212560 336976 212566
rect 336924 212502 336976 212508
rect 336936 202842 336964 212502
rect 337212 205578 337240 220623
rect 337120 205550 337240 205578
rect 336924 202836 336976 202842
rect 336924 202778 336976 202784
rect 337120 196042 337148 205550
rect 337108 196036 337160 196042
rect 337108 195978 337160 195984
rect 337200 195968 337252 195974
rect 337200 195910 337252 195916
rect 336924 193248 336976 193254
rect 336924 193190 336976 193196
rect 336936 183569 336964 193190
rect 337212 186266 337240 195910
rect 337120 186238 337240 186266
rect 336922 183560 336978 183569
rect 337120 183530 337148 186238
rect 336922 183495 336978 183504
rect 337108 183524 337160 183530
rect 337108 183466 337160 183472
rect 336924 173936 336976 173942
rect 336924 173878 336976 173884
rect 336936 125594 336964 173878
rect 337108 172576 337160 172582
rect 337108 172518 337160 172524
rect 337120 169318 337148 172518
rect 337108 169312 337160 169318
rect 337108 169254 337160 169260
rect 337384 169312 337436 169318
rect 337384 169254 337436 169260
rect 337396 162897 337424 169254
rect 337198 162888 337254 162897
rect 337198 162823 337254 162832
rect 337382 162888 337438 162897
rect 337382 162823 337438 162832
rect 337212 158030 337240 162823
rect 337016 158024 337068 158030
rect 337016 157966 337068 157972
rect 337200 158024 337252 158030
rect 337200 157966 337252 157972
rect 337028 147642 337056 157966
rect 337028 147614 337240 147642
rect 337212 143562 337240 147614
rect 337120 143534 337240 143562
rect 337120 138038 337148 143534
rect 337108 138032 337160 138038
rect 337108 137974 337160 137980
rect 337200 137964 337252 137970
rect 337200 137906 337252 137912
rect 337212 132462 337240 137906
rect 337200 132456 337252 132462
rect 337200 132398 337252 132404
rect 336924 125588 336976 125594
rect 336924 125530 336976 125536
rect 336922 115968 336978 115977
rect 336922 115903 336978 115912
rect 336936 86970 336964 115903
rect 337200 114572 337252 114578
rect 337200 114514 337252 114520
rect 337212 110922 337240 114514
rect 337120 110894 337240 110922
rect 337120 99482 337148 110894
rect 337108 99476 337160 99482
rect 337108 99418 337160 99424
rect 337108 99340 337160 99346
rect 337108 99282 337160 99288
rect 337120 95248 337148 99282
rect 337120 95220 337240 95248
rect 337212 86970 337240 95220
rect 336924 86964 336976 86970
rect 336924 86906 336976 86912
rect 337200 86964 337252 86970
rect 337200 86906 337252 86912
rect 337200 77308 337252 77314
rect 337200 77250 337252 77256
rect 336924 75948 336976 75954
rect 336924 75890 336976 75896
rect 336936 66230 336964 75890
rect 336924 66224 336976 66230
rect 336924 66166 336976 66172
rect 337212 56817 337240 77250
rect 338026 76256 338082 76265
rect 338026 76191 338082 76200
rect 338040 76158 338068 76191
rect 338028 76152 338080 76158
rect 338028 76094 338080 76100
rect 337198 56808 337254 56817
rect 337198 56743 337254 56752
rect 337290 56672 337346 56681
rect 336924 56636 336976 56642
rect 337290 56607 337346 56616
rect 336924 56578 336976 56584
rect 336936 46918 336964 56578
rect 337304 56574 337332 56607
rect 337292 56568 337344 56574
rect 337292 56510 337344 56516
rect 337200 47048 337252 47054
rect 337200 46990 337252 46996
rect 337212 46918 337240 46990
rect 336924 46912 336976 46918
rect 336924 46854 336976 46860
rect 337200 46912 337252 46918
rect 337200 46854 337252 46860
rect 337200 37392 337252 37398
rect 337200 37334 337252 37340
rect 336924 37324 336976 37330
rect 336924 37266 336976 37272
rect 336936 33862 336964 37266
rect 337212 37262 337240 37334
rect 337200 37256 337252 37262
rect 337200 37198 337252 37204
rect 337292 37256 337344 37262
rect 337292 37198 337344 37204
rect 336924 33856 336976 33862
rect 336924 33798 336976 33804
rect 336924 19372 336976 19378
rect 336924 19314 336976 19320
rect 336936 8090 336964 19314
rect 337304 18494 337332 37198
rect 337292 18488 337344 18494
rect 337292 18430 337344 18436
rect 337108 18012 337160 18018
rect 337108 17954 337160 17960
rect 336924 8084 336976 8090
rect 336924 8026 336976 8032
rect 336832 6656 336884 6662
rect 336832 6598 336884 6604
rect 337120 6118 337148 17954
rect 337108 6112 337160 6118
rect 337108 6054 337160 6060
rect 337108 5092 337160 5098
rect 337108 5034 337160 5040
rect 335596 3748 336044 3754
rect 335544 3742 336044 3748
rect 335556 3726 336044 3742
rect 335556 3194 335952 3210
rect 335556 3188 335964 3194
rect 335556 3182 335912 3188
rect 335556 2854 335584 3182
rect 335912 3130 335964 3136
rect 335912 3052 335964 3058
rect 335912 2994 335964 3000
rect 335544 2848 335596 2854
rect 335544 2790 335596 2796
rect 335924 480 335952 2994
rect 337120 480 337148 5034
rect 338132 5030 338160 335582
rect 338316 8158 338344 340054
rect 338408 340054 338790 340082
rect 338960 340054 339250 340082
rect 339604 340054 339710 340082
rect 338304 8152 338356 8158
rect 338304 8094 338356 8100
rect 338408 6730 338436 340054
rect 338764 336932 338816 336938
rect 338764 336874 338816 336880
rect 338396 6724 338448 6730
rect 338396 6666 338448 6672
rect 338120 5024 338172 5030
rect 338120 4966 338172 4972
rect 338776 4146 338804 336874
rect 338960 335646 338988 340054
rect 338948 335640 339000 335646
rect 338948 335582 339000 335588
rect 339500 149728 339552 149734
rect 339500 149670 339552 149676
rect 339512 144945 339540 149670
rect 339498 144936 339554 144945
rect 339498 144871 339554 144880
rect 339604 8226 339632 340054
rect 340248 336802 340276 340068
rect 340708 338162 340736 340068
rect 340984 340054 341182 340082
rect 340328 338156 340380 338162
rect 340328 338098 340380 338104
rect 340696 338156 340748 338162
rect 340696 338098 340748 338104
rect 340236 336796 340288 336802
rect 340236 336738 340288 336744
rect 340340 336734 340368 338098
rect 340788 336932 340840 336938
rect 340788 336874 340840 336880
rect 340328 336728 340380 336734
rect 340328 336670 340380 336676
rect 339776 318844 339828 318850
rect 339776 318786 339828 318792
rect 339788 311930 339816 318786
rect 339696 311902 339816 311930
rect 339696 311846 339724 311902
rect 339684 311840 339736 311846
rect 339684 311782 339736 311788
rect 339868 311840 339920 311846
rect 339868 311782 339920 311788
rect 339880 309126 339908 311782
rect 339868 309120 339920 309126
rect 339868 309062 339920 309068
rect 339868 299940 339920 299946
rect 339868 299882 339920 299888
rect 339880 282946 339908 299882
rect 339684 282940 339736 282946
rect 339684 282882 339736 282888
rect 339868 282940 339920 282946
rect 339868 282882 339920 282888
rect 339696 282826 339724 282882
rect 339696 282798 339816 282826
rect 339788 273306 339816 282798
rect 339788 273278 339908 273306
rect 339880 263634 339908 273278
rect 339684 263628 339736 263634
rect 339684 263570 339736 263576
rect 339868 263628 339920 263634
rect 339868 263570 339920 263576
rect 339696 263514 339724 263570
rect 339696 263486 339816 263514
rect 339788 253994 339816 263486
rect 339788 253966 339908 253994
rect 339880 244322 339908 253966
rect 339684 244316 339736 244322
rect 339684 244258 339736 244264
rect 339868 244316 339920 244322
rect 339868 244258 339920 244264
rect 339696 244202 339724 244258
rect 339696 244174 339816 244202
rect 339788 234682 339816 244174
rect 339788 234654 339908 234682
rect 339880 225010 339908 234654
rect 339684 225004 339736 225010
rect 339684 224946 339736 224952
rect 339868 225004 339920 225010
rect 339868 224946 339920 224952
rect 339696 224890 339724 224946
rect 339696 224862 339816 224890
rect 339788 215370 339816 224862
rect 339788 215342 339908 215370
rect 339880 205698 339908 215342
rect 339684 205692 339736 205698
rect 339684 205634 339736 205640
rect 339868 205692 339920 205698
rect 339868 205634 339920 205640
rect 339696 205578 339724 205634
rect 339696 205550 339816 205578
rect 339788 196058 339816 205550
rect 339788 196030 339908 196058
rect 339880 182186 339908 196030
rect 339880 182158 340000 182186
rect 339972 173874 340000 182158
rect 339684 173868 339736 173874
rect 339684 173810 339736 173816
rect 339960 173868 340012 173874
rect 339960 173810 340012 173816
rect 339696 164234 339724 173810
rect 339696 164206 339816 164234
rect 339788 157434 339816 164206
rect 339788 157406 339908 157434
rect 339880 157162 339908 157406
rect 339788 157134 339908 157162
rect 339788 149734 339816 157134
rect 339776 149728 339828 149734
rect 339776 149670 339828 149676
rect 339682 144936 339738 144945
rect 339682 144871 339738 144880
rect 339696 144838 339724 144871
rect 339684 144832 339736 144838
rect 339684 144774 339736 144780
rect 339868 144832 339920 144838
rect 339868 144774 339920 144780
rect 339880 128382 339908 144774
rect 339684 128376 339736 128382
rect 339868 128376 339920 128382
rect 339736 128324 339816 128330
rect 339684 128318 339816 128324
rect 339868 128318 339920 128324
rect 339696 128302 339816 128318
rect 339788 125594 339816 128302
rect 339776 125588 339828 125594
rect 339776 125530 339828 125536
rect 339776 118652 339828 118658
rect 339776 118594 339828 118600
rect 339788 115954 339816 118594
rect 339788 115926 339908 115954
rect 339880 104922 339908 115926
rect 339776 104916 339828 104922
rect 339776 104858 339828 104864
rect 339868 104916 339920 104922
rect 339868 104858 339920 104864
rect 339788 104786 339816 104858
rect 339776 104780 339828 104786
rect 339776 104722 339828 104728
rect 339960 95260 340012 95266
rect 339960 95202 340012 95208
rect 339972 77314 340000 95202
rect 339776 77308 339828 77314
rect 339776 77250 339828 77256
rect 339960 77308 340012 77314
rect 339960 77250 340012 77256
rect 339788 60738 339816 77250
rect 339696 60722 339816 60738
rect 339684 60716 339816 60722
rect 339736 60710 339816 60716
rect 339868 60716 339920 60722
rect 339684 60658 339736 60664
rect 339868 60658 339920 60664
rect 339880 57934 339908 60658
rect 339868 57928 339920 57934
rect 339868 57870 339920 57876
rect 339776 48340 339828 48346
rect 339776 48282 339828 48288
rect 339788 41426 339816 48282
rect 339696 41398 339816 41426
rect 339696 41290 339724 41398
rect 339696 41262 339816 41290
rect 339788 12458 339816 41262
rect 339696 12430 339816 12458
rect 339592 8220 339644 8226
rect 339592 8162 339644 8168
rect 339696 6526 339724 12430
rect 339684 6520 339736 6526
rect 339684 6462 339736 6468
rect 340800 4146 340828 336874
rect 340984 8294 341012 340054
rect 341628 337550 341656 340068
rect 341720 340054 342194 340082
rect 342364 340054 342654 340082
rect 341616 337544 341668 337550
rect 341616 337486 341668 337492
rect 341720 335594 341748 340054
rect 341800 337272 341852 337278
rect 341800 337214 341852 337220
rect 341168 335566 341748 335594
rect 341168 331226 341196 335566
rect 341812 335458 341840 337214
rect 341536 335430 341840 335458
rect 341156 331220 341208 331226
rect 341156 331162 341208 331168
rect 341340 331220 341392 331226
rect 341340 331162 341392 331168
rect 341352 328438 341380 331162
rect 341340 328432 341392 328438
rect 341340 328374 341392 328380
rect 341432 318844 341484 318850
rect 341432 318786 341484 318792
rect 341444 311914 341472 318786
rect 341248 311908 341300 311914
rect 341248 311850 341300 311856
rect 341432 311908 341484 311914
rect 341432 311850 341484 311856
rect 341260 309126 341288 311850
rect 341248 309120 341300 309126
rect 341248 309062 341300 309068
rect 341156 299532 341208 299538
rect 341156 299474 341208 299480
rect 341168 299418 341196 299474
rect 341246 299432 341302 299441
rect 341168 299390 341246 299418
rect 341246 299367 341302 299376
rect 341246 289912 341302 289921
rect 341246 289847 341302 289856
rect 341260 289814 341288 289847
rect 341248 289808 341300 289814
rect 341248 289750 341300 289756
rect 341156 280220 341208 280226
rect 341156 280162 341208 280168
rect 341168 280106 341196 280162
rect 341246 280120 341302 280129
rect 341168 280078 341246 280106
rect 341246 280055 341302 280064
rect 341246 270600 341302 270609
rect 341246 270535 341302 270544
rect 341260 270502 341288 270535
rect 341248 270496 341300 270502
rect 341248 270438 341300 270444
rect 341156 260908 341208 260914
rect 341156 260850 341208 260856
rect 341168 260794 341196 260850
rect 341246 260808 341302 260817
rect 341168 260766 341246 260794
rect 341246 260743 341302 260752
rect 341246 251288 341302 251297
rect 341246 251223 341302 251232
rect 341260 244390 341288 251223
rect 341248 244384 341300 244390
rect 341248 244326 341300 244332
rect 341156 244248 341208 244254
rect 341156 244190 341208 244196
rect 341168 240145 341196 244190
rect 341154 240136 341210 240145
rect 341154 240071 341210 240080
rect 341430 240136 341486 240145
rect 341430 240071 341486 240080
rect 341444 230518 341472 240071
rect 341248 230512 341300 230518
rect 341248 230454 341300 230460
rect 341432 230512 341484 230518
rect 341432 230454 341484 230460
rect 341260 225078 341288 230454
rect 341248 225072 341300 225078
rect 341248 225014 341300 225020
rect 341156 224936 341208 224942
rect 341156 224878 341208 224884
rect 341168 220794 341196 224878
rect 341156 220788 341208 220794
rect 341156 220730 341208 220736
rect 341156 215280 341208 215286
rect 341156 215222 341208 215228
rect 341168 211154 341196 215222
rect 341168 211126 341288 211154
rect 341260 202910 341288 211126
rect 341156 202904 341208 202910
rect 341154 202872 341156 202881
rect 341248 202904 341300 202910
rect 341208 202872 341210 202881
rect 341248 202846 341300 202852
rect 341430 202872 341486 202881
rect 341154 202807 341210 202816
rect 341430 202807 341486 202816
rect 341444 193254 341472 202807
rect 341248 193248 341300 193254
rect 341248 193190 341300 193196
rect 341432 193248 341484 193254
rect 341432 193190 341484 193196
rect 341260 186266 341288 193190
rect 341168 186238 341288 186266
rect 341168 182170 341196 186238
rect 341156 182164 341208 182170
rect 341156 182106 341208 182112
rect 341248 182164 341300 182170
rect 341248 182106 341300 182112
rect 341260 168994 341288 182106
rect 341168 168966 341288 168994
rect 341168 157434 341196 168966
rect 341168 157406 341380 157434
rect 341352 154442 341380 157406
rect 341168 154414 341380 154442
rect 341168 153202 341196 154414
rect 341156 153196 341208 153202
rect 341156 153138 341208 153144
rect 341340 144900 341392 144906
rect 341340 144842 341392 144848
rect 341352 143562 341380 144842
rect 341260 143534 341380 143562
rect 341260 128450 341288 143534
rect 341248 128444 341300 128450
rect 341248 128386 341300 128392
rect 341248 128308 341300 128314
rect 341248 128250 341300 128256
rect 341260 125594 341288 128250
rect 341248 125588 341300 125594
rect 341248 125530 341300 125536
rect 341156 118652 341208 118658
rect 341156 118594 341208 118600
rect 341168 115954 341196 118594
rect 341168 115938 341288 115954
rect 341168 115932 341300 115938
rect 341168 115926 341248 115932
rect 341248 115874 341300 115880
rect 341260 115843 341288 115874
rect 341156 106344 341208 106350
rect 341156 106286 341208 106292
rect 341168 104854 341196 106286
rect 341156 104848 341208 104854
rect 341156 104790 341208 104796
rect 341156 95260 341208 95266
rect 341156 95202 341208 95208
rect 341168 90438 341196 95202
rect 341156 90432 341208 90438
rect 341156 90374 341208 90380
rect 341064 77308 341116 77314
rect 341064 77250 341116 77256
rect 341076 67658 341104 77250
rect 341064 67652 341116 67658
rect 341064 67594 341116 67600
rect 341156 67652 341208 67658
rect 341156 67594 341208 67600
rect 341168 60722 341196 67594
rect 341156 60716 341208 60722
rect 341156 60658 341208 60664
rect 341340 60716 341392 60722
rect 341340 60658 341392 60664
rect 341352 53122 341380 60658
rect 341260 53094 341380 53122
rect 341260 48346 341288 53094
rect 341248 48340 341300 48346
rect 341248 48282 341300 48288
rect 341432 48340 341484 48346
rect 341432 48282 341484 48288
rect 341444 46918 341472 48282
rect 341432 46912 341484 46918
rect 341432 46854 341484 46860
rect 341248 37324 341300 37330
rect 341248 37266 341300 37272
rect 341260 32298 341288 37266
rect 341248 32292 341300 32298
rect 341248 32234 341300 32240
rect 341248 29096 341300 29102
rect 341168 29044 341248 29050
rect 341168 29038 341300 29044
rect 341168 29022 341288 29038
rect 341168 27606 341196 29022
rect 341156 27600 341208 27606
rect 341156 27542 341208 27548
rect 341248 9716 341300 9722
rect 341248 9658 341300 9664
rect 340972 8288 341024 8294
rect 340972 8230 341024 8236
rect 341260 6458 341288 9658
rect 341248 6452 341300 6458
rect 341248 6394 341300 6400
rect 338764 4140 338816 4146
rect 338764 4082 338816 4088
rect 339500 4140 339552 4146
rect 339500 4082 339552 4088
rect 340788 4140 340840 4146
rect 340788 4082 340840 4088
rect 338304 3732 338356 3738
rect 338304 3674 338356 3680
rect 338316 480 338344 3674
rect 339512 480 339540 4082
rect 341536 3806 341564 335430
rect 342364 6186 342392 340054
rect 342720 337544 342772 337550
rect 342718 337512 342720 337521
rect 342772 337512 342774 337521
rect 342718 337447 342774 337456
rect 342904 337204 342956 337210
rect 342904 337146 342956 337152
rect 342352 6180 342404 6186
rect 342352 6122 342404 6128
rect 342916 3874 342944 337146
rect 343100 336802 343128 340068
rect 343088 336796 343140 336802
rect 343088 336738 343140 336744
rect 343652 6390 343680 340068
rect 344112 337482 344140 340068
rect 344572 337686 344600 340068
rect 345138 340054 345244 340082
rect 344560 337680 344612 337686
rect 344560 337622 344612 337628
rect 344376 337544 344428 337550
rect 344376 337486 344428 337492
rect 344100 337476 344152 337482
rect 344100 337418 344152 337424
rect 344284 336864 344336 336870
rect 344284 336806 344336 336812
rect 343640 6384 343692 6390
rect 343640 6326 343692 6332
rect 342904 3868 342956 3874
rect 342904 3810 342956 3816
rect 343088 3868 343140 3874
rect 343088 3810 343140 3816
rect 341524 3800 341576 3806
rect 341524 3742 341576 3748
rect 341892 3800 341944 3806
rect 341892 3742 341944 3748
rect 340696 3188 340748 3194
rect 340696 3130 340748 3136
rect 340708 480 340736 3130
rect 341904 480 341932 3742
rect 343100 480 343128 3810
rect 344296 3482 344324 336806
rect 344204 3454 344324 3482
rect 344204 2990 344232 3454
rect 344388 3346 344416 337486
rect 345216 6254 345244 340054
rect 345584 337618 345612 340068
rect 345676 340054 346058 340082
rect 345572 337612 345624 337618
rect 345572 337554 345624 337560
rect 345676 336818 345704 340054
rect 345756 337612 345808 337618
rect 345756 337554 345808 337560
rect 345768 337521 345796 337554
rect 345754 337512 345810 337521
rect 345754 337447 345810 337456
rect 345940 336932 345992 336938
rect 345584 336802 345704 336818
rect 345572 336796 345704 336802
rect 345624 336790 345704 336796
rect 345860 336892 345940 336920
rect 345572 336738 345624 336744
rect 345860 331242 345888 336892
rect 345940 336874 345992 336880
rect 345676 331214 345888 331242
rect 345204 6248 345256 6254
rect 345204 6190 345256 6196
rect 345676 4146 345704 331214
rect 346596 5302 346624 340068
rect 347056 337890 347084 340068
rect 347044 337884 347096 337890
rect 347044 337826 347096 337832
rect 347516 337482 347544 340068
rect 347976 340054 348082 340082
rect 347504 337476 347556 337482
rect 347504 337418 347556 337424
rect 347780 87032 347832 87038
rect 347778 87000 347780 87009
rect 347832 87000 347834 87009
rect 347778 86935 347834 86944
rect 347780 29096 347832 29102
rect 347778 29064 347780 29073
rect 347832 29064 347834 29073
rect 347778 28999 347834 29008
rect 347778 16960 347834 16969
rect 347778 16895 347780 16904
rect 347832 16895 347834 16904
rect 347780 16866 347832 16872
rect 347976 5370 348004 340054
rect 348528 338706 348556 340068
rect 348516 338700 348568 338706
rect 348516 338642 348568 338648
rect 348424 337884 348476 337890
rect 348424 337826 348476 337832
rect 347964 5364 348016 5370
rect 347964 5306 348016 5312
rect 346584 5296 346636 5302
rect 346584 5238 346636 5244
rect 345664 4140 345716 4146
rect 345664 4082 345716 4088
rect 347872 4140 347924 4146
rect 347872 4082 347924 4088
rect 344296 3330 344416 3346
rect 344284 3324 344416 3330
rect 344336 3318 344416 3324
rect 344284 3266 344336 3272
rect 346676 3188 346728 3194
rect 346676 3130 346728 3136
rect 344192 2984 344244 2990
rect 344192 2926 344244 2932
rect 344284 2916 344336 2922
rect 344284 2858 344336 2864
rect 344296 480 344324 2858
rect 345480 604 345532 610
rect 345480 546 345532 552
rect 345492 480 345520 546
rect 346688 480 346716 3130
rect 347884 480 347912 4082
rect 348436 3262 348464 337826
rect 348988 337278 349016 340068
rect 349356 340054 349554 340082
rect 349068 337476 349120 337482
rect 349068 337418 349120 337424
rect 348976 337272 349028 337278
rect 348976 337214 349028 337220
rect 349080 4146 349108 337418
rect 349356 5438 349384 340054
rect 350000 337686 350028 340068
rect 350184 340054 350474 340082
rect 350644 340054 351026 340082
rect 349988 337680 350040 337686
rect 349988 337622 350040 337628
rect 350184 337618 350212 340054
rect 350172 337612 350224 337618
rect 350172 337554 350224 337560
rect 350644 6322 350672 340054
rect 351184 337612 351236 337618
rect 351184 337554 351236 337560
rect 350632 6316 350684 6322
rect 350632 6258 350684 6264
rect 349344 5432 349396 5438
rect 349344 5374 349396 5380
rect 351196 4146 351224 337554
rect 351472 336802 351500 340068
rect 351932 337822 351960 340068
rect 352116 340054 352498 340082
rect 351920 337816 351972 337822
rect 351920 337758 351972 337764
rect 351828 337544 351880 337550
rect 351828 337486 351880 337492
rect 351460 336796 351512 336802
rect 351460 336738 351512 336744
rect 351840 4146 351868 337486
rect 352116 5506 352144 340054
rect 352944 337958 352972 340068
rect 352932 337952 352984 337958
rect 352932 337894 352984 337900
rect 353404 337006 353432 340068
rect 353496 340054 353970 340082
rect 353392 337000 353444 337006
rect 353392 336942 353444 336948
rect 352564 336796 352616 336802
rect 352564 336738 352616 336744
rect 352104 5500 352156 5506
rect 352104 5442 352156 5448
rect 352576 4146 352604 336738
rect 352656 16924 352708 16930
rect 352656 16866 352708 16872
rect 352668 16697 352696 16866
rect 352654 16688 352710 16697
rect 352654 16623 352710 16632
rect 353496 4418 353524 340054
rect 354416 338094 354444 340068
rect 354404 338088 354456 338094
rect 354404 338030 354456 338036
rect 354876 337686 354904 340068
rect 354968 340054 355442 340082
rect 354864 337680 354916 337686
rect 354864 337622 354916 337628
rect 353484 4412 353536 4418
rect 353484 4354 353536 4360
rect 354968 4350 354996 340054
rect 355888 338026 355916 340068
rect 356256 340054 356362 340082
rect 356624 340054 356914 340082
rect 355876 338020 355928 338026
rect 355876 337962 355928 337968
rect 355324 337952 355376 337958
rect 355324 337894 355376 337900
rect 354956 4344 355008 4350
rect 354956 4286 355008 4292
rect 349068 4140 349120 4146
rect 349068 4082 349120 4088
rect 351184 4140 351236 4146
rect 351184 4082 351236 4088
rect 351368 4140 351420 4146
rect 351368 4082 351420 4088
rect 351828 4140 351880 4146
rect 351828 4082 351880 4088
rect 351920 4140 351972 4146
rect 351920 4082 351972 4088
rect 352564 4140 352616 4146
rect 352564 4082 352616 4088
rect 350264 3324 350316 3330
rect 350264 3266 350316 3272
rect 348424 3256 348476 3262
rect 348424 3198 348476 3204
rect 349068 3256 349120 3262
rect 349068 3198 349120 3204
rect 349080 480 349108 3198
rect 350276 480 350304 3266
rect 351380 480 351408 4082
rect 351932 2990 351960 4082
rect 355336 3670 355364 337894
rect 355968 337204 356020 337210
rect 355968 337146 356020 337152
rect 355324 3664 355376 3670
rect 355324 3606 355376 3612
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 351920 2984 351972 2990
rect 351920 2926 351972 2932
rect 352564 2984 352616 2990
rect 352564 2926 352616 2932
rect 352576 480 352604 2926
rect 353772 480 353800 3334
rect 355980 2922 356008 337146
rect 356152 332852 356204 332858
rect 356152 332794 356204 332800
rect 356164 4282 356192 332794
rect 356152 4276 356204 4282
rect 356152 4218 356204 4224
rect 356256 3369 356284 340054
rect 356624 332858 356652 340054
rect 356704 337748 356756 337754
rect 356704 337690 356756 337696
rect 356612 332852 356664 332858
rect 356612 332794 356664 332800
rect 356242 3360 356298 3369
rect 356242 3295 356298 3304
rect 356716 3262 356744 337690
rect 357360 336870 357388 340068
rect 357348 336864 357400 336870
rect 357348 336806 357400 336812
rect 357820 336802 357848 340068
rect 358004 340054 358386 340082
rect 357808 336796 357860 336802
rect 357808 336738 357860 336744
rect 358004 331242 358032 340054
rect 358084 338088 358136 338094
rect 358084 338030 358136 338036
rect 357636 331214 358032 331242
rect 357636 331208 357664 331214
rect 357452 331180 357664 331208
rect 357452 323626 357480 331180
rect 357452 323598 357572 323626
rect 357544 311930 357572 323598
rect 357544 311902 357848 311930
rect 357820 302326 357848 311902
rect 357808 302320 357860 302326
rect 357808 302262 357860 302268
rect 357900 302116 357952 302122
rect 357900 302058 357952 302064
rect 357912 292602 357940 302058
rect 357440 292596 357492 292602
rect 357440 292538 357492 292544
rect 357900 292596 357952 292602
rect 357900 292538 357952 292544
rect 357452 282946 357480 292538
rect 357440 282940 357492 282946
rect 357440 282882 357492 282888
rect 357716 282804 357768 282810
rect 357716 282746 357768 282752
rect 357728 273170 357756 282746
rect 357452 273142 357756 273170
rect 357452 263616 357480 273142
rect 357452 263588 357664 263616
rect 357636 263514 357664 263588
rect 357544 263486 357664 263514
rect 357544 253910 357572 263486
rect 357532 253904 357584 253910
rect 357532 253846 357584 253852
rect 357716 253904 357768 253910
rect 357716 253846 357768 253852
rect 357728 241534 357756 253846
rect 357624 241528 357676 241534
rect 357624 241470 357676 241476
rect 357716 241528 357768 241534
rect 357716 241470 357768 241476
rect 357636 234682 357664 241470
rect 357544 234654 357664 234682
rect 357544 234598 357572 234654
rect 357532 234592 357584 234598
rect 357532 234534 357584 234540
rect 357716 234592 357768 234598
rect 357716 234534 357768 234540
rect 357728 231826 357756 234534
rect 357636 231798 357756 231826
rect 357636 212566 357664 231798
rect 357624 212560 357676 212566
rect 357624 212502 357676 212508
rect 357716 212560 357768 212566
rect 357716 212502 357768 212508
rect 357728 205578 357756 212502
rect 357636 205550 357756 205578
rect 357636 196058 357664 205550
rect 357544 196030 357664 196058
rect 357544 195974 357572 196030
rect 357532 195968 357584 195974
rect 357532 195910 357584 195916
rect 357716 195968 357768 195974
rect 357716 195910 357768 195916
rect 357728 180878 357756 195910
rect 357624 180872 357676 180878
rect 357624 180814 357676 180820
rect 357716 180872 357768 180878
rect 357716 180814 357768 180820
rect 357636 176798 357664 180814
rect 357624 176792 357676 176798
rect 357624 176734 357676 176740
rect 357624 176656 357676 176662
rect 357624 176598 357676 176604
rect 357636 167686 357664 176598
rect 357440 167680 357492 167686
rect 357440 167622 357492 167628
rect 357624 167680 357676 167686
rect 357624 167622 357676 167628
rect 357452 162874 357480 167622
rect 357452 162846 357572 162874
rect 357544 162790 357572 162846
rect 357532 162784 357584 162790
rect 357532 162726 357584 162732
rect 357624 162784 357676 162790
rect 357624 162726 357676 162732
rect 357636 153218 357664 162726
rect 357636 153190 357756 153218
rect 357728 147642 357756 153190
rect 357544 147614 357756 147642
rect 357544 140026 357572 147614
rect 357452 139998 357572 140026
rect 357452 125769 357480 139998
rect 357438 125760 357494 125769
rect 357438 125695 357494 125704
rect 357530 125624 357586 125633
rect 357530 125559 357586 125568
rect 357544 114646 357572 125559
rect 357532 114640 357584 114646
rect 357532 114582 357584 114588
rect 357440 114572 357492 114578
rect 357440 114514 357492 114520
rect 357452 114458 357480 114514
rect 357452 114430 357572 114458
rect 357544 104922 357572 114430
rect 357532 104916 357584 104922
rect 357532 104858 357584 104864
rect 357716 104916 357768 104922
rect 357716 104858 357768 104864
rect 357346 87272 357402 87281
rect 357346 87207 357402 87216
rect 357360 87038 357388 87207
rect 357348 87032 357400 87038
rect 357348 86974 357400 86980
rect 357728 80170 357756 104858
rect 357716 80164 357768 80170
rect 357716 80106 357768 80112
rect 357624 80096 357676 80102
rect 357624 80038 357676 80044
rect 357636 72434 357664 80038
rect 357636 72406 357756 72434
rect 357728 56642 357756 72406
rect 357532 56636 357584 56642
rect 357532 56578 357584 56584
rect 357716 56636 357768 56642
rect 357716 56578 357768 56584
rect 357544 56506 357572 56578
rect 357532 56500 357584 56506
rect 357532 56442 357584 56448
rect 357624 46980 357676 46986
rect 357624 46922 357676 46928
rect 357636 46850 357664 46922
rect 357624 46844 357676 46850
rect 357624 46786 357676 46792
rect 357624 37324 357676 37330
rect 357624 37266 357676 37272
rect 357636 32434 357664 37266
rect 357624 32428 357676 32434
rect 357624 32370 357676 32376
rect 357808 32428 357860 32434
rect 357808 32370 357860 32376
rect 357346 29336 357402 29345
rect 357346 29271 357402 29280
rect 357360 29102 357388 29271
rect 357348 29096 357400 29102
rect 357348 29038 357400 29044
rect 357820 27713 357848 32370
rect 357622 27704 357678 27713
rect 357622 27639 357678 27648
rect 357806 27704 357862 27713
rect 357806 27639 357862 27648
rect 357636 27606 357664 27639
rect 357624 27600 357676 27606
rect 357624 27542 357676 27548
rect 357716 18012 357768 18018
rect 357716 17954 357768 17960
rect 357728 4214 357756 17954
rect 357716 4208 357768 4214
rect 357716 4150 357768 4156
rect 358096 3670 358124 338030
rect 358728 337680 358780 337686
rect 358728 337622 358780 337628
rect 358740 328438 358768 337622
rect 358728 328432 358780 328438
rect 358728 328374 358780 328380
rect 358728 318844 358780 318850
rect 358728 318786 358780 318792
rect 358740 317422 358768 318786
rect 358728 317416 358780 317422
rect 358728 317358 358780 317364
rect 358728 307828 358780 307834
rect 358728 307770 358780 307776
rect 358740 298110 358768 307770
rect 358728 298104 358780 298110
rect 358728 298046 358780 298052
rect 358728 280288 358780 280294
rect 358728 280230 358780 280236
rect 358740 278769 358768 280230
rect 358542 278760 358598 278769
rect 358542 278695 358598 278704
rect 358726 278760 358782 278769
rect 358726 278695 358782 278704
rect 358556 269142 358584 278695
rect 358544 269136 358596 269142
rect 358544 269078 358596 269084
rect 358636 269136 358688 269142
rect 358636 269078 358688 269084
rect 358648 260930 358676 269078
rect 358648 260902 358768 260930
rect 358740 259418 358768 260902
rect 358728 259412 358780 259418
rect 358728 259354 358780 259360
rect 358740 240174 358768 240205
rect 358728 240168 358780 240174
rect 358648 240116 358728 240122
rect 358648 240110 358780 240116
rect 358648 240094 358768 240110
rect 358648 230518 358676 240094
rect 358452 230512 358504 230518
rect 358636 230512 358688 230518
rect 358504 230460 358584 230466
rect 358452 230454 358584 230460
rect 358636 230454 358688 230460
rect 358464 230450 358584 230454
rect 358464 230444 358596 230450
rect 358464 230438 358544 230444
rect 358544 230386 358596 230392
rect 358728 220856 358780 220862
rect 358726 220824 358728 220833
rect 358780 220824 358782 220833
rect 358726 220759 358782 220768
rect 358726 211168 358782 211177
rect 358726 211103 358782 211112
rect 358740 201482 358768 211103
rect 358452 201476 358504 201482
rect 358452 201418 358504 201424
rect 358728 201476 358780 201482
rect 358728 201418 358780 201424
rect 358464 191865 358492 201418
rect 358450 191856 358506 191865
rect 358450 191791 358506 191800
rect 358634 191856 358690 191865
rect 358634 191791 358690 191800
rect 358648 183598 358676 191791
rect 358636 183592 358688 183598
rect 358636 183534 358688 183540
rect 358728 183592 358780 183598
rect 358728 183534 358780 183540
rect 358740 182170 358768 183534
rect 358544 182164 358596 182170
rect 358544 182106 358596 182112
rect 358728 182164 358780 182170
rect 358728 182106 358780 182112
rect 358556 172553 358584 182106
rect 358542 172544 358598 172553
rect 358542 172479 358598 172488
rect 358726 172544 358782 172553
rect 358726 172479 358782 172488
rect 358740 162858 358768 172479
rect 358544 162852 358596 162858
rect 358544 162794 358596 162800
rect 358728 162852 358780 162858
rect 358728 162794 358780 162800
rect 358556 153241 358584 162794
rect 358542 153232 358598 153241
rect 358542 153167 358598 153176
rect 358726 153232 358782 153241
rect 358726 153167 358782 153176
rect 358740 135250 358768 153167
rect 358728 135244 358780 135250
rect 358728 135186 358780 135192
rect 358728 125656 358780 125662
rect 358728 125598 358780 125604
rect 358740 114578 358768 125598
rect 358636 114572 358688 114578
rect 358636 114514 358688 114520
rect 358728 114572 358780 114578
rect 358728 114514 358780 114520
rect 358648 106350 358676 114514
rect 358636 106344 358688 106350
rect 358636 106286 358688 106292
rect 358728 106208 358780 106214
rect 358728 106150 358780 106156
rect 358740 104786 358768 106150
rect 358728 104780 358780 104786
rect 358728 104722 358780 104728
rect 358726 87000 358782 87009
rect 358726 86935 358782 86944
rect 358740 85542 358768 86935
rect 358728 85536 358780 85542
rect 358728 85478 358780 85484
rect 358832 77382 358860 340068
rect 358924 340054 359306 340082
rect 359476 340054 359766 340082
rect 358924 77382 358952 340054
rect 359476 337362 359504 340054
rect 359200 337334 359504 337362
rect 359200 327321 359228 337334
rect 359464 337272 359516 337278
rect 359464 337214 359516 337220
rect 359186 327312 359242 327321
rect 359186 327247 359242 327256
rect 359186 327176 359242 327185
rect 359186 327111 359242 327120
rect 359200 327078 359228 327111
rect 359188 327072 359240 327078
rect 359188 327014 359240 327020
rect 359188 317756 359240 317762
rect 359188 317698 359240 317704
rect 359200 307850 359228 317698
rect 359200 307822 359320 307850
rect 359292 299606 359320 307822
rect 359280 299600 359332 299606
rect 359280 299542 359332 299548
rect 359096 299464 359148 299470
rect 359096 299406 359148 299412
rect 359108 298110 359136 299406
rect 359096 298104 359148 298110
rect 359096 298046 359148 298052
rect 359188 288448 359240 288454
rect 359188 288390 359240 288396
rect 359200 280242 359228 288390
rect 359108 280214 359228 280242
rect 359108 280158 359136 280214
rect 359096 280152 359148 280158
rect 359096 280094 359148 280100
rect 359188 280152 359240 280158
rect 359188 280094 359240 280100
rect 359200 263514 359228 280094
rect 359108 263486 359228 263514
rect 359108 253994 359136 263486
rect 359016 253966 359136 253994
rect 359016 253910 359044 253966
rect 359004 253904 359056 253910
rect 359004 253846 359056 253852
rect 359188 253904 359240 253910
rect 359188 253846 359240 253852
rect 359200 241534 359228 253846
rect 359096 241528 359148 241534
rect 359096 241470 359148 241476
rect 359188 241528 359240 241534
rect 359188 241470 359240 241476
rect 359108 234682 359136 241470
rect 359016 234654 359136 234682
rect 359016 234598 359044 234654
rect 359004 234592 359056 234598
rect 359004 234534 359056 234540
rect 359188 234592 359240 234598
rect 359188 234534 359240 234540
rect 359200 222222 359228 234534
rect 359096 222216 359148 222222
rect 359096 222158 359148 222164
rect 359188 222216 359240 222222
rect 359188 222158 359240 222164
rect 359108 212566 359136 222158
rect 359096 212560 359148 212566
rect 359096 212502 359148 212508
rect 359188 212560 359240 212566
rect 359188 212502 359240 212508
rect 359200 205578 359228 212502
rect 359108 205550 359228 205578
rect 359108 196058 359136 205550
rect 359016 196030 359136 196058
rect 359016 195974 359044 196030
rect 359004 195968 359056 195974
rect 359004 195910 359056 195916
rect 359188 195968 359240 195974
rect 359188 195910 359240 195916
rect 359200 183598 359228 195910
rect 359096 183592 359148 183598
rect 359096 183534 359148 183540
rect 359188 183592 359240 183598
rect 359188 183534 359240 183540
rect 359108 157350 359136 183534
rect 359096 157344 359148 157350
rect 359096 157286 359148 157292
rect 359188 157276 359240 157282
rect 359188 157218 359240 157224
rect 359200 147642 359228 157218
rect 359108 147614 359228 147642
rect 359108 140026 359136 147614
rect 359108 139998 359228 140026
rect 359200 128330 359228 139998
rect 359108 128302 359228 128330
rect 359108 124166 359136 128302
rect 359096 124160 359148 124166
rect 359096 124102 359148 124108
rect 359188 124160 359240 124166
rect 359188 124102 359240 124108
rect 359200 106298 359228 124102
rect 359108 106270 359228 106298
rect 359004 104780 359056 104786
rect 359004 104722 359056 104728
rect 359016 87009 359044 104722
rect 359108 101402 359136 106270
rect 359108 101374 359320 101402
rect 359292 99226 359320 101374
rect 359200 99198 359320 99226
rect 359002 87000 359058 87009
rect 359002 86935 359058 86944
rect 359200 80170 359228 99198
rect 359188 80164 359240 80170
rect 359188 80106 359240 80112
rect 359096 80096 359148 80102
rect 359096 80038 359148 80044
rect 358820 77376 358872 77382
rect 358820 77318 358872 77324
rect 358912 77376 358964 77382
rect 358912 77318 358964 77324
rect 358820 77240 358872 77246
rect 358820 77182 358872 77188
rect 358912 77240 358964 77246
rect 358912 77182 358964 77188
rect 358728 67652 358780 67658
rect 358728 67594 358780 67600
rect 358740 66230 358768 67594
rect 358728 66224 358780 66230
rect 358728 66166 358780 66172
rect 358636 56636 358688 56642
rect 358636 56578 358688 56584
rect 358648 48346 358676 56578
rect 358636 48340 358688 48346
rect 358636 48282 358688 48288
rect 358728 48340 358780 48346
rect 358728 48282 358780 48288
rect 358740 46918 358768 48282
rect 358728 46912 358780 46918
rect 358728 46854 358780 46860
rect 358636 37324 358688 37330
rect 358636 37266 358688 37272
rect 358648 29034 358676 37266
rect 358636 29028 358688 29034
rect 358636 28970 358688 28976
rect 358728 29028 358780 29034
rect 358728 28970 358780 28976
rect 358740 27606 358768 28970
rect 358728 27600 358780 27606
rect 358728 27542 358780 27548
rect 358544 9716 358596 9722
rect 358544 9658 358596 9664
rect 358084 3664 358136 3670
rect 358084 3606 358136 3612
rect 356704 3256 356756 3262
rect 356704 3198 356756 3204
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 354956 2916 355008 2922
rect 354956 2858 355008 2864
rect 355968 2916 356020 2922
rect 355968 2858 356020 2864
rect 354968 480 354996 2858
rect 356152 2848 356204 2854
rect 356152 2790 356204 2796
rect 356164 480 356192 2790
rect 357360 480 357388 3198
rect 358556 480 358584 9658
rect 358832 4010 358860 77182
rect 358924 4078 358952 77182
rect 359004 75948 359056 75954
rect 359004 75890 359056 75896
rect 359016 67658 359044 75890
rect 359108 72434 359136 80038
rect 359108 72406 359228 72434
rect 359004 67652 359056 67658
rect 359004 67594 359056 67600
rect 359200 48362 359228 72406
rect 359108 48334 359228 48362
rect 359108 46918 359136 48334
rect 359096 46912 359148 46918
rect 359096 46854 359148 46860
rect 359004 37324 359056 37330
rect 359004 37266 359056 37272
rect 359016 34134 359044 37266
rect 359004 34128 359056 34134
rect 359004 34070 359056 34076
rect 359096 34060 359148 34066
rect 359096 34002 359148 34008
rect 359108 27606 359136 34002
rect 359096 27600 359148 27606
rect 359096 27542 359148 27548
rect 359188 27600 359240 27606
rect 359188 27542 359240 27548
rect 359200 4758 359228 27542
rect 359188 4752 359240 4758
rect 359188 4694 359240 4700
rect 358912 4072 358964 4078
rect 358912 4014 358964 4020
rect 358820 4004 358872 4010
rect 358820 3946 358872 3952
rect 359476 2922 359504 337214
rect 360304 336938 360332 340068
rect 360764 337754 360792 340068
rect 360948 340054 361238 340082
rect 360752 337748 360804 337754
rect 360752 337690 360804 337696
rect 360292 336932 360344 336938
rect 360292 336874 360344 336880
rect 360948 331242 360976 340054
rect 361776 337346 361804 340068
rect 361868 340054 362250 340082
rect 362328 340054 362710 340082
rect 363156 340054 363262 340082
rect 361764 337340 361816 337346
rect 361764 337282 361816 337288
rect 361672 333328 361724 333334
rect 361672 333270 361724 333276
rect 360304 331226 360976 331242
rect 360292 331220 360976 331226
rect 360344 331214 360476 331220
rect 360292 331162 360344 331168
rect 360528 331214 360976 331220
rect 360476 331162 360528 331168
rect 360488 321586 360516 331162
rect 360304 321558 360516 321586
rect 360304 321450 360332 321558
rect 360304 321422 360424 321450
rect 360396 311930 360424 321422
rect 360304 311902 360424 311930
rect 360304 311794 360332 311902
rect 360304 311766 360424 311794
rect 360396 302274 360424 311766
rect 360396 302246 360516 302274
rect 360488 282946 360516 302246
rect 360292 282940 360344 282946
rect 360292 282882 360344 282888
rect 360476 282940 360528 282946
rect 360476 282882 360528 282888
rect 360304 282826 360332 282882
rect 360304 282798 360424 282826
rect 360396 273306 360424 282798
rect 360396 273278 360516 273306
rect 360488 263634 360516 273278
rect 360292 263628 360344 263634
rect 360292 263570 360344 263576
rect 360476 263628 360528 263634
rect 360476 263570 360528 263576
rect 360304 263514 360332 263570
rect 360304 263486 360424 263514
rect 360396 253994 360424 263486
rect 360396 253966 360516 253994
rect 360488 244322 360516 253966
rect 360292 244316 360344 244322
rect 360292 244258 360344 244264
rect 360476 244316 360528 244322
rect 360476 244258 360528 244264
rect 360304 244202 360332 244258
rect 360304 244174 360424 244202
rect 360396 234682 360424 244174
rect 360396 234654 360516 234682
rect 360488 225010 360516 234654
rect 360292 225004 360344 225010
rect 360292 224946 360344 224952
rect 360476 225004 360528 225010
rect 360476 224946 360528 224952
rect 360304 224890 360332 224946
rect 360304 224862 360424 224890
rect 360396 215370 360424 224862
rect 360396 215342 360516 215370
rect 360488 205698 360516 215342
rect 360292 205692 360344 205698
rect 360292 205634 360344 205640
rect 360476 205692 360528 205698
rect 360476 205634 360528 205640
rect 360304 205578 360332 205634
rect 360304 205550 360424 205578
rect 360396 196058 360424 205550
rect 360396 196030 360516 196058
rect 360488 193225 360516 196030
rect 360474 193216 360530 193225
rect 360474 193151 360530 193160
rect 360658 193216 360714 193225
rect 360658 193151 360714 193160
rect 360672 183598 360700 193151
rect 360476 183592 360528 183598
rect 360476 183534 360528 183540
rect 360660 183592 360712 183598
rect 360660 183534 360712 183540
rect 360488 182170 360516 183534
rect 360476 182164 360528 182170
rect 360476 182106 360528 182112
rect 360660 182164 360712 182170
rect 360660 182106 360712 182112
rect 360672 172530 360700 182106
rect 360580 172502 360700 172530
rect 360580 162897 360608 172502
rect 360198 162888 360254 162897
rect 360198 162823 360254 162832
rect 360566 162888 360622 162897
rect 360566 162823 360622 162832
rect 360212 153241 360240 162823
rect 360198 153232 360254 153241
rect 360198 153167 360254 153176
rect 360382 153232 360438 153241
rect 360382 153167 360438 153176
rect 360396 147762 360424 153167
rect 360384 147756 360436 147762
rect 360384 147698 360436 147704
rect 360200 144900 360252 144906
rect 360200 144842 360252 144848
rect 360212 124234 360240 144842
rect 360200 124228 360252 124234
rect 360200 124170 360252 124176
rect 360384 124228 360436 124234
rect 360384 124170 360436 124176
rect 360396 119354 360424 124170
rect 360304 119326 360424 119354
rect 360304 118538 360332 119326
rect 360304 118510 360516 118538
rect 360488 106457 360516 118510
rect 360474 106448 360530 106457
rect 360474 106383 360530 106392
rect 360382 106312 360438 106321
rect 360382 106247 360384 106256
rect 360436 106247 360438 106256
rect 360568 106276 360620 106282
rect 360384 106218 360436 106224
rect 360568 106218 360620 106224
rect 360580 96665 360608 106218
rect 360290 96656 360346 96665
rect 360290 96591 360292 96600
rect 360344 96591 360346 96600
rect 360566 96656 360622 96665
rect 360566 96591 360622 96600
rect 360292 96562 360344 96568
rect 360292 89684 360344 89690
rect 360292 89626 360344 89632
rect 360304 86986 360332 89626
rect 360304 86958 360424 86986
rect 360396 86902 360424 86958
rect 360200 86896 360252 86902
rect 360200 86838 360252 86844
rect 360384 86896 360436 86902
rect 360384 86838 360436 86844
rect 360212 72434 360240 86838
rect 360212 72406 360332 72434
rect 360304 60722 360332 72406
rect 360292 60716 360344 60722
rect 360292 60658 360344 60664
rect 360476 60716 360528 60722
rect 360476 60658 360528 60664
rect 360488 48414 360516 60658
rect 360476 48408 360528 48414
rect 360476 48350 360528 48356
rect 360384 48340 360436 48346
rect 360384 48282 360436 48288
rect 360396 41426 360424 48282
rect 360304 41410 360424 41426
rect 360292 41404 360424 41410
rect 360344 41398 360424 41404
rect 360476 41404 360528 41410
rect 360292 41346 360344 41352
rect 360476 41346 360528 41352
rect 360488 12458 360516 41346
rect 360304 12430 360516 12458
rect 360304 4690 360332 12430
rect 361684 4894 361712 333270
rect 361672 4888 361724 4894
rect 361672 4830 361724 4836
rect 360292 4684 360344 4690
rect 360292 4626 360344 4632
rect 359740 4004 359792 4010
rect 359740 3946 359792 3952
rect 359464 2916 359516 2922
rect 359464 2858 359516 2864
rect 359752 480 359780 3946
rect 360936 3664 360988 3670
rect 360936 3606 360988 3612
rect 360948 480 360976 3606
rect 361868 3466 361896 340054
rect 362224 336864 362276 336870
rect 362224 336806 362276 336812
rect 361856 3460 361908 3466
rect 361856 3402 361908 3408
rect 362132 3188 362184 3194
rect 362132 3130 362184 3136
rect 362144 480 362172 3130
rect 362236 3126 362264 336806
rect 362328 333334 362356 340054
rect 362868 337816 362920 337822
rect 362868 337758 362920 337764
rect 362316 333328 362368 333334
rect 362316 333270 362368 333276
rect 362880 3194 362908 337758
rect 363052 335640 363104 335646
rect 363052 335582 363104 335588
rect 363064 4826 363092 335582
rect 363052 4820 363104 4826
rect 363052 4762 363104 4768
rect 363156 3534 363184 340054
rect 363708 337278 363736 340068
rect 363800 340054 364182 340082
rect 363696 337272 363748 337278
rect 363696 337214 363748 337220
rect 363604 336796 363656 336802
rect 363604 336738 363656 336744
rect 363616 3602 363644 336738
rect 363800 335646 363828 340054
rect 364248 338020 364300 338026
rect 364248 337962 364300 337968
rect 363788 335640 363840 335646
rect 363788 335582 363840 335588
rect 363604 3596 363656 3602
rect 363604 3538 363656 3544
rect 363144 3528 363196 3534
rect 363144 3470 363196 3476
rect 364260 3194 364288 337962
rect 364720 336802 364748 340068
rect 365180 336870 365208 340068
rect 365640 337890 365668 340068
rect 365824 340054 366206 340082
rect 365628 337884 365680 337890
rect 365628 337826 365680 337832
rect 365168 336864 365220 336870
rect 365168 336806 365220 336812
rect 364708 336796 364760 336802
rect 364708 336738 364760 336744
rect 364340 157616 364392 157622
rect 364338 157584 364340 157593
rect 364392 157584 364394 157593
rect 364338 157519 364394 157528
rect 365720 4072 365772 4078
rect 365720 4014 365772 4020
rect 362868 3188 362920 3194
rect 362868 3130 362920 3136
rect 363328 3188 363380 3194
rect 363328 3130 363380 3136
rect 364248 3188 364300 3194
rect 364248 3130 364300 3136
rect 364524 3188 364576 3194
rect 364524 3130 364576 3136
rect 362224 3120 362276 3126
rect 362224 3062 362276 3068
rect 363340 480 363368 3130
rect 364536 480 364564 3130
rect 365732 480 365760 4014
rect 365824 3942 365852 340054
rect 366652 337142 366680 340068
rect 367126 340054 367232 340082
rect 367008 337340 367060 337346
rect 367008 337282 367060 337288
rect 366640 337136 366692 337142
rect 366640 337078 366692 337084
rect 366916 337000 366968 337006
rect 366916 336942 366968 336948
rect 366928 12510 366956 336942
rect 367020 270706 367048 337282
rect 367008 270700 367060 270706
rect 367008 270642 367060 270648
rect 367008 270564 367060 270570
rect 367008 270506 367060 270512
rect 367020 251190 367048 270506
rect 367008 251184 367060 251190
rect 367008 251126 367060 251132
rect 367008 241528 367060 241534
rect 367008 241470 367060 241476
rect 367020 222193 367048 241470
rect 367006 222184 367062 222193
rect 367006 222119 367062 222128
rect 367006 212664 367062 212673
rect 367006 212599 367062 212608
rect 367020 193186 367048 212599
rect 367008 193180 367060 193186
rect 367008 193122 367060 193128
rect 367008 183592 367060 183598
rect 367008 183534 367060 183540
rect 367020 144906 367048 183534
rect 367008 144900 367060 144906
rect 367008 144842 367060 144848
rect 367008 135312 367060 135318
rect 367008 135254 367060 135260
rect 367020 115938 367048 135254
rect 367008 115932 367060 115938
rect 367008 115874 367060 115880
rect 367008 106344 367060 106350
rect 367008 106286 367060 106292
rect 367020 96626 367048 106286
rect 367008 96620 367060 96626
rect 367008 96562 367060 96568
rect 367098 87136 367154 87145
rect 367098 87071 367154 87080
rect 367008 87032 367060 87038
rect 367112 87009 367140 87071
rect 367008 86974 367060 86980
rect 367098 87000 367154 87009
rect 367020 77489 367048 86974
rect 367098 86935 367154 86944
rect 367006 77480 367062 77489
rect 367006 77415 367062 77424
rect 367006 77344 367062 77353
rect 367006 77279 367062 77288
rect 367020 67794 367048 77279
rect 367008 67788 367060 67794
rect 367008 67730 367060 67736
rect 367008 67652 367060 67658
rect 367008 67594 367060 67600
rect 367020 66230 367048 67594
rect 367008 66224 367060 66230
rect 367008 66166 367060 66172
rect 367100 63776 367152 63782
rect 367098 63744 367100 63753
rect 367152 63744 367154 63753
rect 367098 63679 367154 63688
rect 367008 48340 367060 48346
rect 367008 48282 367060 48288
rect 367020 46918 367048 48282
rect 367008 46912 367060 46918
rect 367008 46854 367060 46860
rect 367100 40248 367152 40254
rect 367098 40216 367100 40225
rect 367152 40216 367154 40225
rect 367098 40151 367154 40160
rect 367008 37324 367060 37330
rect 367008 37266 367060 37272
rect 367020 29170 367048 37266
rect 367100 29232 367152 29238
rect 367100 29174 367152 29180
rect 367008 29164 367060 29170
rect 367008 29106 367060 29112
rect 367112 29073 367140 29174
rect 367098 29064 367154 29073
rect 367008 29028 367060 29034
rect 367098 28999 367154 29008
rect 367008 28970 367060 28976
rect 367020 27606 367048 28970
rect 367008 27600 367060 27606
rect 367008 27542 367060 27548
rect 367006 16960 367062 16969
rect 367006 16895 367062 16904
rect 367020 16833 367048 16895
rect 367006 16824 367062 16833
rect 367006 16759 367062 16768
rect 366916 12504 366968 12510
rect 366916 12446 366968 12452
rect 366916 12368 366968 12374
rect 366916 12310 366968 12316
rect 366824 9716 366876 9722
rect 366824 9658 366876 9664
rect 365812 3936 365864 3942
rect 365812 3878 365864 3884
rect 366836 2802 366864 9658
rect 366928 4078 366956 12310
rect 367204 4962 367232 340054
rect 367664 337074 367692 340068
rect 367940 340054 368138 340082
rect 367652 337068 367704 337074
rect 367652 337010 367704 337016
rect 367940 335646 367968 340054
rect 367284 335640 367336 335646
rect 367284 335582 367336 335588
rect 367928 335640 367980 335646
rect 367928 335582 367980 335588
rect 367192 4956 367244 4962
rect 367192 4898 367244 4904
rect 366916 4072 366968 4078
rect 366916 4014 366968 4020
rect 367296 3058 367324 335582
rect 368584 5098 368612 340068
rect 368676 340054 369150 340082
rect 368572 5092 368624 5098
rect 368572 5034 368624 5040
rect 368676 3534 368704 340054
rect 369124 337136 369176 337142
rect 369124 337078 369176 337084
rect 369136 3874 369164 337078
rect 369596 336938 369624 340068
rect 370056 337958 370084 340068
rect 370148 340054 370622 340082
rect 370044 337952 370096 337958
rect 370044 337894 370096 337900
rect 369768 337408 369820 337414
rect 369768 337350 369820 337356
rect 369584 336932 369636 336938
rect 369584 336874 369636 336880
rect 369676 16856 369728 16862
rect 369674 16824 369676 16833
rect 369728 16824 369730 16833
rect 369674 16759 369730 16768
rect 369780 4078 369808 337350
rect 369860 76152 369912 76158
rect 369858 76120 369860 76129
rect 369912 76120 369914 76129
rect 369858 76055 369914 76064
rect 369216 4072 369268 4078
rect 369216 4014 369268 4020
rect 369768 4072 369820 4078
rect 369768 4014 369820 4020
rect 369124 3868 369176 3874
rect 369124 3810 369176 3816
rect 368664 3528 368716 3534
rect 368664 3470 368716 3476
rect 368020 3460 368072 3466
rect 368020 3402 368072 3408
rect 367284 3052 367336 3058
rect 367284 2994 367336 3000
rect 366836 2774 366956 2802
rect 366928 480 366956 2774
rect 368032 480 368060 3402
rect 369228 480 369256 4014
rect 370148 3806 370176 340054
rect 371068 337142 371096 340068
rect 371528 338094 371556 340068
rect 371516 338088 371568 338094
rect 371516 338030 371568 338036
rect 371148 337612 371200 337618
rect 371148 337554 371200 337560
rect 371056 337136 371108 337142
rect 371056 337078 371108 337084
rect 370504 336796 370556 336802
rect 370504 336738 370556 336744
rect 370412 4140 370464 4146
rect 370412 4082 370464 4088
rect 370136 3800 370188 3806
rect 370136 3742 370188 3748
rect 370424 480 370452 4082
rect 370516 3738 370544 336738
rect 371160 4146 371188 337554
rect 372080 337482 372108 340068
rect 372068 337476 372120 337482
rect 372068 337418 372120 337424
rect 372540 336802 372568 340068
rect 373000 337278 373028 340068
rect 373276 340054 373566 340082
rect 374026 340054 374316 340082
rect 372988 337272 373040 337278
rect 372988 337214 373040 337220
rect 372528 336796 372580 336802
rect 372528 336738 372580 336744
rect 373276 328506 373304 340054
rect 373908 337680 373960 337686
rect 373908 337622 373960 337628
rect 372712 328500 372764 328506
rect 372712 328442 372764 328448
rect 373264 328500 373316 328506
rect 373264 328442 373316 328448
rect 372724 318782 372752 328442
rect 372712 318776 372764 318782
rect 372712 318718 372764 318724
rect 372712 309188 372764 309194
rect 372712 309130 372764 309136
rect 372724 299470 372752 309130
rect 372712 299464 372764 299470
rect 372712 299406 372764 299412
rect 372712 289876 372764 289882
rect 372712 289818 372764 289824
rect 372724 280158 372752 289818
rect 372712 280152 372764 280158
rect 372712 280094 372764 280100
rect 372712 270564 372764 270570
rect 372712 270506 372764 270512
rect 372724 260846 372752 270506
rect 372712 260840 372764 260846
rect 372712 260782 372764 260788
rect 372712 251252 372764 251258
rect 372712 251194 372764 251200
rect 372724 241505 372752 251194
rect 372526 241496 372582 241505
rect 372526 241431 372582 241440
rect 372710 241496 372766 241505
rect 372710 241431 372766 241440
rect 372540 231878 372568 241431
rect 372528 231872 372580 231878
rect 372528 231814 372580 231820
rect 372712 231872 372764 231878
rect 372712 231814 372764 231820
rect 372724 222193 372752 231814
rect 372526 222184 372582 222193
rect 372526 222119 372582 222128
rect 372710 222184 372766 222193
rect 372710 222119 372766 222128
rect 372540 212566 372568 222119
rect 372528 212560 372580 212566
rect 372528 212502 372580 212508
rect 372712 212560 372764 212566
rect 372712 212502 372764 212508
rect 372724 202881 372752 212502
rect 372526 202872 372582 202881
rect 372526 202807 372582 202816
rect 372710 202872 372766 202881
rect 372710 202807 372766 202816
rect 372540 193254 372568 202807
rect 372528 193248 372580 193254
rect 372528 193190 372580 193196
rect 372712 193248 372764 193254
rect 372712 193190 372764 193196
rect 372724 176662 372752 193190
rect 372712 176656 372764 176662
rect 372712 176598 372764 176604
rect 372804 176588 372856 176594
rect 372804 176530 372856 176536
rect 372816 173913 372844 176530
rect 372802 173904 372858 173913
rect 372802 173839 372858 173848
rect 372986 173904 373042 173913
rect 372986 173839 373042 173848
rect 373000 164257 373028 173839
rect 372802 164248 372858 164257
rect 372802 164183 372804 164192
rect 372856 164183 372858 164192
rect 372986 164248 373042 164257
rect 372986 164183 373042 164192
rect 372804 164154 372856 164160
rect 373816 157616 373868 157622
rect 373814 157584 373816 157593
rect 373868 157584 373870 157593
rect 373814 157519 373870 157528
rect 372804 157344 372856 157350
rect 372804 157286 372856 157292
rect 372816 138174 372844 157286
rect 372804 138168 372856 138174
rect 372804 138110 372856 138116
rect 372712 135312 372764 135318
rect 372712 135254 372764 135260
rect 372724 118726 372752 135254
rect 372712 118720 372764 118726
rect 372712 118662 372764 118668
rect 372712 118584 372764 118590
rect 372712 118526 372764 118532
rect 372724 106282 372752 118526
rect 372712 106276 372764 106282
rect 372712 106218 372764 106224
rect 372804 106276 372856 106282
rect 372804 106218 372856 106224
rect 372816 80170 372844 106218
rect 372804 80164 372856 80170
rect 372804 80106 372856 80112
rect 372712 80096 372764 80102
rect 372712 80038 372764 80044
rect 372724 70394 372752 80038
rect 372632 70366 372752 70394
rect 372632 70258 372660 70366
rect 372632 70230 372752 70258
rect 372724 51082 372752 70230
rect 372632 51054 372752 51082
rect 372632 50946 372660 51054
rect 372632 50918 372752 50946
rect 372724 31770 372752 50918
rect 372632 31742 372752 31770
rect 372632 31634 372660 31742
rect 372632 31606 372752 31634
rect 372724 12458 372752 31606
rect 372632 12430 372752 12458
rect 371148 4140 371200 4146
rect 371148 4082 371200 4088
rect 372632 4078 372660 12430
rect 372620 4072 372672 4078
rect 372620 4014 372672 4020
rect 371608 3936 371660 3942
rect 371608 3878 371660 3884
rect 370504 3732 370556 3738
rect 370504 3674 370556 3680
rect 371620 480 371648 3878
rect 373920 3874 373948 337622
rect 374092 335640 374144 335646
rect 374092 335582 374144 335588
rect 372804 3868 372856 3874
rect 372804 3810 372856 3816
rect 373908 3868 373960 3874
rect 373908 3810 373960 3816
rect 372816 480 372844 3810
rect 374000 3800 374052 3806
rect 374000 3742 374052 3748
rect 374012 480 374040 3742
rect 374104 2990 374132 335582
rect 374288 3330 374316 340054
rect 374472 337550 374500 340068
rect 374656 340054 375038 340082
rect 374460 337544 374512 337550
rect 374460 337486 374512 337492
rect 374656 335646 374684 340054
rect 375288 337544 375340 337550
rect 375288 337486 375340 337492
rect 374644 335640 374696 335646
rect 374644 335582 374696 335588
rect 375300 3806 375328 337486
rect 375380 96620 375432 96626
rect 375380 96562 375432 96568
rect 375392 87009 375420 96562
rect 375378 87000 375434 87009
rect 375378 86935 375434 86944
rect 375288 3800 375340 3806
rect 375288 3742 375340 3748
rect 375196 3732 375248 3738
rect 375196 3674 375248 3680
rect 374276 3324 374328 3330
rect 374276 3266 374328 3272
rect 374092 2984 374144 2990
rect 374092 2926 374144 2932
rect 375208 480 375236 3674
rect 375484 3398 375512 340068
rect 375944 337754 375972 340068
rect 376128 340054 376510 340082
rect 375932 337748 375984 337754
rect 375932 337690 375984 337696
rect 376024 336796 376076 336802
rect 376024 336738 376076 336744
rect 375656 328500 375708 328506
rect 375656 328442 375708 328448
rect 375668 313970 375696 328442
rect 375576 313942 375696 313970
rect 375576 309233 375604 313942
rect 375562 309224 375618 309233
rect 375562 309159 375618 309168
rect 375746 309224 375802 309233
rect 375746 309159 375802 309168
rect 375760 299470 375788 309159
rect 375748 299464 375800 299470
rect 375748 299406 375800 299412
rect 375656 289876 375708 289882
rect 375656 289818 375708 289824
rect 375668 282962 375696 289818
rect 375576 282934 375696 282962
rect 375576 282826 375604 282934
rect 375576 282798 375696 282826
rect 375668 263650 375696 282798
rect 375576 263622 375696 263650
rect 375576 263514 375604 263622
rect 375576 263486 375696 263514
rect 375668 244338 375696 263486
rect 375576 244310 375696 244338
rect 375576 244202 375604 244310
rect 375576 244174 375696 244202
rect 375668 225026 375696 244174
rect 375576 224998 375696 225026
rect 375576 224890 375604 224998
rect 375576 224862 375696 224890
rect 375668 205714 375696 224862
rect 375576 205686 375696 205714
rect 375576 205578 375604 205686
rect 375576 205550 375696 205578
rect 375668 186402 375696 205550
rect 375576 186374 375696 186402
rect 375576 186266 375604 186374
rect 375576 186238 375788 186266
rect 375760 157434 375788 186238
rect 375576 157406 375788 157434
rect 375576 157298 375604 157406
rect 375576 157270 375696 157298
rect 375668 157162 375696 157270
rect 375668 157134 375788 157162
rect 375760 138106 375788 157134
rect 375748 138100 375800 138106
rect 375748 138042 375800 138048
rect 375656 138032 375708 138038
rect 375656 137974 375708 137980
rect 375668 128466 375696 137974
rect 375576 128438 375696 128466
rect 375576 128330 375604 128438
rect 375576 128302 375696 128330
rect 375668 109070 375696 128302
rect 375656 109064 375708 109070
rect 375656 109006 375708 109012
rect 375564 108996 375616 109002
rect 375564 108938 375616 108944
rect 375576 106321 375604 108938
rect 375562 106312 375618 106321
rect 375562 106247 375618 106256
rect 375746 106312 375802 106321
rect 375746 106247 375802 106256
rect 375760 99346 375788 106247
rect 375564 99340 375616 99346
rect 375564 99282 375616 99288
rect 375748 99340 375800 99346
rect 375748 99282 375800 99288
rect 375576 96626 375604 99282
rect 375564 96620 375616 96626
rect 375564 96562 375616 96568
rect 375654 87000 375710 87009
rect 375654 86935 375710 86944
rect 375668 86902 375696 86935
rect 375564 86896 375616 86902
rect 375564 86838 375616 86844
rect 375656 86896 375708 86902
rect 375656 86838 375708 86844
rect 375576 80152 375604 86838
rect 375576 80124 375696 80152
rect 375668 67590 375696 80124
rect 375656 67584 375708 67590
rect 375656 67526 375708 67532
rect 375656 62008 375708 62014
rect 375656 61950 375708 61956
rect 375668 41426 375696 61950
rect 375576 41398 375696 41426
rect 375576 41290 375604 41398
rect 375576 41262 375696 41290
rect 375668 12458 375696 41262
rect 375576 12430 375696 12458
rect 375472 3392 375524 3398
rect 375472 3334 375524 3340
rect 375576 2854 375604 12430
rect 376036 3262 376064 336738
rect 376128 328506 376156 340054
rect 376956 336802 376984 340068
rect 377416 337822 377444 340068
rect 377508 340054 377890 340082
rect 377404 337816 377456 337822
rect 377404 337758 377456 337764
rect 376944 336796 376996 336802
rect 376944 336738 376996 336744
rect 377508 335594 377536 340054
rect 378048 337000 378100 337006
rect 378048 336942 378100 336948
rect 377680 336796 377732 336802
rect 377680 336738 377732 336744
rect 377140 335566 377536 335594
rect 376116 328500 376168 328506
rect 376116 328442 376168 328448
rect 377140 321638 377168 335566
rect 377692 331242 377720 336738
rect 377416 331214 377720 331242
rect 377128 321632 377180 321638
rect 377128 321574 377180 321580
rect 377220 321428 377272 321434
rect 377220 321370 377272 321376
rect 377232 289882 377260 321370
rect 377128 289876 377180 289882
rect 377128 289818 377180 289824
rect 377220 289876 377272 289882
rect 377220 289818 377272 289824
rect 377140 280158 377168 289818
rect 377128 280152 377180 280158
rect 377128 280094 377180 280100
rect 377128 270564 377180 270570
rect 377128 270506 377180 270512
rect 377140 260846 377168 270506
rect 377128 260840 377180 260846
rect 377128 260782 377180 260788
rect 377128 251252 377180 251258
rect 377128 251194 377180 251200
rect 377140 241505 377168 251194
rect 376942 241496 376998 241505
rect 376942 241431 376998 241440
rect 377126 241496 377182 241505
rect 377126 241431 377182 241440
rect 376956 231878 376984 241431
rect 376944 231872 376996 231878
rect 376944 231814 376996 231820
rect 377128 231872 377180 231878
rect 377128 231814 377180 231820
rect 377140 222193 377168 231814
rect 376942 222184 376998 222193
rect 376942 222119 376998 222128
rect 377126 222184 377182 222193
rect 377126 222119 377182 222128
rect 376956 212566 376984 222119
rect 376944 212560 376996 212566
rect 376944 212502 376996 212508
rect 377128 212560 377180 212566
rect 377128 212502 377180 212508
rect 377140 202881 377168 212502
rect 376942 202872 376998 202881
rect 376942 202807 376998 202816
rect 377126 202872 377182 202881
rect 377126 202807 377182 202816
rect 376956 193254 376984 202807
rect 376944 193248 376996 193254
rect 376944 193190 376996 193196
rect 377128 193248 377180 193254
rect 377128 193190 377180 193196
rect 377140 183569 377168 193190
rect 376942 183560 376998 183569
rect 376942 183495 376998 183504
rect 377126 183560 377182 183569
rect 377126 183495 377182 183504
rect 376956 173942 376984 183495
rect 376944 173936 376996 173942
rect 376944 173878 376996 173884
rect 377036 173936 377088 173942
rect 377036 173878 377088 173884
rect 377048 166954 377076 173878
rect 377048 166926 377168 166954
rect 377140 157350 377168 166926
rect 377128 157344 377180 157350
rect 377128 157286 377180 157292
rect 377220 157276 377272 157282
rect 377220 157218 377272 157224
rect 377232 140078 377260 157218
rect 377220 140072 377272 140078
rect 377220 140014 377272 140020
rect 377128 135312 377180 135318
rect 377128 135254 377180 135260
rect 377140 118726 377168 135254
rect 377128 118720 377180 118726
rect 377128 118662 377180 118668
rect 377128 118584 377180 118590
rect 377128 118526 377180 118532
rect 377140 115938 377168 118526
rect 376944 115932 376996 115938
rect 376944 115874 376996 115880
rect 377128 115932 377180 115938
rect 377128 115874 377180 115880
rect 376956 106457 376984 115874
rect 376942 106448 376998 106457
rect 376942 106383 376998 106392
rect 377126 106448 377182 106457
rect 377126 106383 377182 106392
rect 377140 106264 377168 106383
rect 377048 106236 377168 106264
rect 377048 99414 377076 106236
rect 377036 99408 377088 99414
rect 377036 99350 377088 99356
rect 377128 99340 377180 99346
rect 377128 99282 377180 99288
rect 376666 76256 376722 76265
rect 376666 76191 376722 76200
rect 376680 76158 376708 76191
rect 376668 76152 376720 76158
rect 376668 76094 376720 76100
rect 377140 70514 377168 99282
rect 377128 70508 377180 70514
rect 377128 70450 377180 70456
rect 377128 67652 377180 67658
rect 377128 67594 377180 67600
rect 376666 63880 376722 63889
rect 376666 63815 376722 63824
rect 376680 63782 376708 63815
rect 376668 63776 376720 63782
rect 376668 63718 376720 63724
rect 377140 51762 377168 67594
rect 377140 51734 377260 51762
rect 377232 46986 377260 51734
rect 377220 46980 377272 46986
rect 377220 46922 377272 46928
rect 377312 46980 377364 46986
rect 377312 46922 377364 46928
rect 376666 40352 376722 40361
rect 376666 40287 376722 40296
rect 376680 40254 376708 40287
rect 376668 40248 376720 40254
rect 376668 40190 376720 40196
rect 377324 38622 377352 46922
rect 377128 38616 377180 38622
rect 377128 38558 377180 38564
rect 377312 38616 377364 38622
rect 377312 38558 377364 38564
rect 377140 31822 377168 38558
rect 377128 31816 377180 31822
rect 377128 31758 377180 31764
rect 377128 31680 377180 31686
rect 377128 31622 377180 31628
rect 376666 29336 376722 29345
rect 376666 29271 376722 29280
rect 376680 29238 376708 29271
rect 376668 29232 376720 29238
rect 376668 29174 376720 29180
rect 377140 22166 377168 31622
rect 377128 22160 377180 22166
rect 377128 22102 377180 22108
rect 377036 22092 377088 22098
rect 377036 22034 377088 22040
rect 376666 16960 376722 16969
rect 376666 16895 376722 16904
rect 376680 16862 376708 16895
rect 376668 16856 376720 16862
rect 376668 16798 376720 16804
rect 377048 9625 377076 22034
rect 376758 9616 376814 9625
rect 376758 9551 376814 9560
rect 377034 9616 377090 9625
rect 377034 9551 377090 9560
rect 376772 4078 376800 9551
rect 376760 4072 376812 4078
rect 376760 4014 376812 4020
rect 377416 3670 377444 331214
rect 378060 4146 378088 336942
rect 378428 336802 378456 340068
rect 378888 338094 378916 340068
rect 378876 338088 378928 338094
rect 378876 338030 378928 338036
rect 379348 338026 379376 340068
rect 379716 340054 379914 340082
rect 379336 338020 379388 338026
rect 379336 337962 379388 337968
rect 378416 336796 378468 336802
rect 378416 336738 378468 336744
rect 378508 63912 378560 63918
rect 378506 63880 378508 63889
rect 378560 63880 378562 63889
rect 378506 63815 378562 63824
rect 377588 4140 377640 4146
rect 377588 4082 377640 4088
rect 378048 4140 378100 4146
rect 378048 4082 378100 4088
rect 378784 4140 378836 4146
rect 378784 4082 378836 4088
rect 377404 3664 377456 3670
rect 377404 3606 377456 3612
rect 376024 3256 376076 3262
rect 376024 3198 376076 3204
rect 376392 3052 376444 3058
rect 376392 2994 376444 3000
rect 375564 2848 375616 2854
rect 375564 2790 375616 2796
rect 376404 480 376432 2994
rect 377600 480 377628 4082
rect 378796 480 378824 4082
rect 379716 3466 379744 340054
rect 380360 337958 380388 340068
rect 380348 337952 380400 337958
rect 380348 337894 380400 337900
rect 380820 337346 380848 340068
rect 380808 337340 380860 337346
rect 380808 337282 380860 337288
rect 380808 337136 380860 337142
rect 380808 337078 380860 337084
rect 380164 336796 380216 336802
rect 380164 336738 380216 336744
rect 380176 4418 380204 336738
rect 380164 4412 380216 4418
rect 380164 4354 380216 4360
rect 380820 4146 380848 337078
rect 381372 336802 381400 340068
rect 381832 337482 381860 340068
rect 382292 337618 382320 340068
rect 382280 337612 382332 337618
rect 382280 337554 382332 337560
rect 381820 337476 381872 337482
rect 381820 337418 381872 337424
rect 382188 337000 382240 337006
rect 382188 336942 382240 336948
rect 381636 336864 381688 336870
rect 381636 336806 381688 336812
rect 381360 336796 381412 336802
rect 381360 336738 381412 336744
rect 381544 336796 381596 336802
rect 381544 336738 381596 336744
rect 381556 4826 381584 336738
rect 381544 4820 381596 4826
rect 381544 4762 381596 4768
rect 379980 4140 380032 4146
rect 379980 4082 380032 4088
rect 380808 4140 380860 4146
rect 380808 4082 380860 4088
rect 381176 4140 381228 4146
rect 381176 4082 381228 4088
rect 379704 3460 379756 3466
rect 379704 3402 379756 3408
rect 379992 480 380020 4082
rect 381188 480 381216 4082
rect 381648 3058 381676 336806
rect 382200 4146 382228 336942
rect 382844 336802 382872 340068
rect 383304 337686 383332 340068
rect 383292 337680 383344 337686
rect 383292 337622 383344 337628
rect 383764 337550 383792 340068
rect 383856 340054 384330 340082
rect 383752 337544 383804 337550
rect 383752 337486 383804 337492
rect 382832 336796 382884 336802
rect 382832 336738 382884 336744
rect 382188 4140 382240 4146
rect 382188 4082 382240 4088
rect 383568 4140 383620 4146
rect 383568 4082 383620 4088
rect 382372 4004 382424 4010
rect 382372 3946 382424 3952
rect 381636 3052 381688 3058
rect 381636 2994 381688 3000
rect 382384 480 382412 3946
rect 383580 480 383608 4082
rect 383856 3738 383884 340054
rect 384304 336932 384356 336938
rect 384304 336874 384356 336880
rect 384316 4146 384344 336874
rect 384776 336870 384804 340068
rect 385236 337210 385264 340068
rect 385328 340054 385802 340082
rect 385224 337204 385276 337210
rect 385224 337146 385276 337152
rect 384764 336864 384816 336870
rect 384764 336806 384816 336812
rect 384948 336864 385000 336870
rect 384948 336806 385000 336812
rect 384304 4140 384356 4146
rect 384304 4082 384356 4088
rect 383844 3732 383896 3738
rect 383844 3674 383896 3680
rect 384960 610 384988 336806
rect 385328 3942 385356 340054
rect 386248 337142 386276 340068
rect 386236 337136 386288 337142
rect 386236 337078 386288 337084
rect 386708 337006 386736 340068
rect 386696 337000 386748 337006
rect 386696 336942 386748 336948
rect 386800 325961 386828 340190
rect 387720 336938 387748 340068
rect 387708 336932 387760 336938
rect 387708 336874 387760 336880
rect 388180 336870 388208 340068
rect 388444 337816 388496 337822
rect 388444 337758 388496 337764
rect 388168 336864 388220 336870
rect 388168 336806 388220 336812
rect 387064 336796 387116 336802
rect 387064 336738 387116 336744
rect 386786 325952 386842 325961
rect 386786 325887 386842 325896
rect 386786 325816 386842 325825
rect 386786 325751 386842 325760
rect 386800 325689 386828 325751
rect 386786 325680 386842 325689
rect 386786 325615 386842 325624
rect 386970 325680 387026 325689
rect 386970 325615 387026 325624
rect 386984 316130 387012 325615
rect 386788 316124 386840 316130
rect 386788 316066 386840 316072
rect 386972 316124 387024 316130
rect 386972 316066 387024 316072
rect 386800 315994 386828 316066
rect 386788 315988 386840 315994
rect 386788 315930 386840 315936
rect 386788 302116 386840 302122
rect 386788 302058 386840 302064
rect 386800 293078 386828 302058
rect 386788 293072 386840 293078
rect 386788 293014 386840 293020
rect 386788 282804 386840 282810
rect 386788 282746 386840 282752
rect 386800 278730 386828 282746
rect 386788 278724 386840 278730
rect 386788 278666 386840 278672
rect 386788 263492 386840 263498
rect 386788 263434 386840 263440
rect 386800 254046 386828 263434
rect 386788 254040 386840 254046
rect 386788 253982 386840 253988
rect 386696 253904 386748 253910
rect 386696 253846 386748 253852
rect 386708 244202 386736 253846
rect 386524 244174 386736 244202
rect 386524 234682 386552 244174
rect 386432 234654 386552 234682
rect 386432 231849 386460 234654
rect 386418 231840 386474 231849
rect 386418 231775 386474 231784
rect 386786 231840 386842 231849
rect 386786 231775 386842 231784
rect 386800 222222 386828 231775
rect 386604 222216 386656 222222
rect 386604 222158 386656 222164
rect 386788 222216 386840 222222
rect 386788 222158 386840 222164
rect 386616 215354 386644 222158
rect 386420 215348 386472 215354
rect 386420 215290 386472 215296
rect 386604 215348 386656 215354
rect 386604 215290 386656 215296
rect 386432 212537 386460 215290
rect 386418 212528 386474 212537
rect 386418 212463 386474 212472
rect 386602 212528 386658 212537
rect 386602 212463 386658 212472
rect 386616 202881 386644 212463
rect 386602 202872 386658 202881
rect 386602 202807 386658 202816
rect 386878 202872 386934 202881
rect 386878 202807 386934 202816
rect 386892 193254 386920 202807
rect 386696 193248 386748 193254
rect 386696 193190 386748 193196
rect 386880 193248 386932 193254
rect 386880 193190 386932 193196
rect 386708 186266 386736 193190
rect 386616 186238 386736 186266
rect 386616 183569 386644 186238
rect 386602 183560 386658 183569
rect 386602 183495 386658 183504
rect 386970 183560 387026 183569
rect 386970 183495 387026 183504
rect 386984 173942 387012 183495
rect 386788 173936 386840 173942
rect 386788 173878 386840 173884
rect 386972 173936 387024 173942
rect 386972 173878 387024 173884
rect 386800 166954 386828 173878
rect 386708 166926 386828 166954
rect 386708 164218 386736 166926
rect 386512 164212 386564 164218
rect 386512 164154 386564 164160
rect 386696 164212 386748 164218
rect 386696 164154 386748 164160
rect 386418 157992 386474 158001
rect 386418 157927 386474 157936
rect 386432 157729 386460 157927
rect 386418 157720 386474 157729
rect 386418 157655 386474 157664
rect 386524 154601 386552 164154
rect 386510 154592 386566 154601
rect 386510 154527 386566 154536
rect 386786 154592 386842 154601
rect 386786 154527 386842 154536
rect 386800 147642 386828 154527
rect 386524 147614 386828 147642
rect 386524 144906 386552 147614
rect 386512 144900 386564 144906
rect 386512 144842 386564 144848
rect 386696 144900 386748 144906
rect 386696 144842 386748 144848
rect 386708 135289 386736 144842
rect 386418 135280 386474 135289
rect 386418 135215 386474 135224
rect 386694 135280 386750 135289
rect 386694 135215 386750 135224
rect 386432 128330 386460 135215
rect 386432 128302 386644 128330
rect 386616 115977 386644 128302
rect 386418 115968 386474 115977
rect 386418 115903 386474 115912
rect 386602 115968 386658 115977
rect 386602 115903 386658 115912
rect 386432 109018 386460 115903
rect 386432 108990 386552 109018
rect 386524 106282 386552 108990
rect 386512 106276 386564 106282
rect 386512 106218 386564 106224
rect 386512 99340 386564 99346
rect 386512 99282 386564 99288
rect 386524 96642 386552 99282
rect 386524 96614 386644 96642
rect 386616 89758 386644 96614
rect 386420 89752 386472 89758
rect 386604 89752 386656 89758
rect 386472 89700 386604 89706
rect 386420 89694 386656 89700
rect 386432 89678 386644 89694
rect 386616 79914 386644 89678
rect 386616 79886 386736 79914
rect 386708 77246 386736 79886
rect 386696 77240 386748 77246
rect 386696 77182 386748 77188
rect 386418 76528 386474 76537
rect 386418 76463 386474 76472
rect 386432 76265 386460 76463
rect 386418 76256 386474 76265
rect 386418 76191 386474 76200
rect 386604 67652 386656 67658
rect 386604 67594 386656 67600
rect 386328 63912 386380 63918
rect 386326 63880 386328 63889
rect 386380 63880 386382 63889
rect 386326 63815 386382 63824
rect 386616 60738 386644 67594
rect 386432 60710 386644 60738
rect 386432 51066 386460 60710
rect 386420 51060 386472 51066
rect 386420 51002 386472 51008
rect 386604 51060 386656 51066
rect 386604 51002 386656 51008
rect 386616 41426 386644 51002
rect 386616 41398 386736 41426
rect 386708 37369 386736 41398
rect 386510 37360 386566 37369
rect 386510 37295 386566 37304
rect 386694 37360 386750 37369
rect 386694 37295 386750 37304
rect 386524 31822 386552 37295
rect 386512 31816 386564 31822
rect 386512 31758 386564 31764
rect 386604 31680 386656 31686
rect 386604 31622 386656 31628
rect 386616 26246 386644 31622
rect 386604 26240 386656 26246
rect 386604 26182 386656 26188
rect 386326 17232 386382 17241
rect 386326 17167 386382 17176
rect 386340 16833 386368 17167
rect 386326 16824 386382 16833
rect 386326 16759 386382 16768
rect 386236 16652 386288 16658
rect 386236 16594 386288 16600
rect 386248 12374 386276 16594
rect 386236 12368 386288 12374
rect 386236 12310 386288 12316
rect 386604 12368 386656 12374
rect 386604 12310 386656 12316
rect 385868 4072 385920 4078
rect 385868 4014 385920 4020
rect 385316 3936 385368 3942
rect 385316 3878 385368 3884
rect 384672 604 384724 610
rect 384672 546 384724 552
rect 384948 604 385000 610
rect 384948 546 385000 552
rect 384684 480 384712 546
rect 385880 480 385908 4014
rect 386616 4010 386644 12310
rect 387076 4078 387104 336738
rect 388260 4140 388312 4146
rect 388260 4082 388312 4088
rect 387064 4072 387116 4078
rect 387064 4014 387116 4020
rect 386604 4004 386656 4010
rect 386604 3946 386656 3952
rect 387064 2780 387116 2786
rect 387064 2722 387116 2728
rect 387076 480 387104 2722
rect 388272 480 388300 4082
rect 388456 2854 388484 337758
rect 388732 336802 388760 340068
rect 389192 337822 389220 340068
rect 389284 340054 389666 340082
rect 389836 340054 390218 340082
rect 390572 340054 390678 340082
rect 390848 340054 391138 340082
rect 391690 340054 391888 340082
rect 392150 340054 392440 340082
rect 389180 337816 389232 337822
rect 389180 337758 389232 337764
rect 389284 337668 389312 340054
rect 389836 337770 389864 340054
rect 389100 337640 389312 337668
rect 389376 337742 389864 337770
rect 388720 336796 388772 336802
rect 388720 336738 388772 336744
rect 389100 4146 389128 337640
rect 389088 4140 389140 4146
rect 389088 4082 389140 4088
rect 388444 2848 388496 2854
rect 388444 2790 388496 2796
rect 389376 626 389404 337742
rect 390572 626 390600 340054
rect 390848 3534 390876 340054
rect 391860 337668 391888 340054
rect 391860 337640 392164 337668
rect 390836 3528 390888 3534
rect 390836 3470 390888 3476
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 389376 598 389496 626
rect 390572 598 390692 626
rect 389468 480 389496 598
rect 390664 480 390692 598
rect 391860 480 391888 3470
rect 392136 610 392164 337640
rect 392412 336802 392440 340054
rect 392596 337754 392624 340068
rect 392584 337748 392636 337754
rect 392584 337690 392636 337696
rect 392400 336796 392452 336802
rect 392400 336738 392452 336744
rect 393148 3738 393176 340068
rect 393228 337748 393280 337754
rect 393228 337690 393280 337696
rect 393136 3732 393188 3738
rect 393136 3674 393188 3680
rect 393240 3126 393268 337690
rect 393608 337686 393636 340068
rect 394068 337754 394096 340068
rect 394528 340054 394634 340082
rect 394056 337748 394108 337754
rect 394056 337690 394108 337696
rect 393596 337680 393648 337686
rect 393596 337622 393648 337628
rect 393596 336796 393648 336802
rect 393596 336738 393648 336744
rect 393228 3120 393280 3126
rect 393228 3062 393280 3068
rect 393608 2938 393636 336738
rect 394528 3534 394556 340054
rect 394608 337748 394660 337754
rect 394608 337690 394660 337696
rect 394516 3528 394568 3534
rect 394516 3470 394568 3476
rect 394620 3058 394648 337690
rect 395080 337550 395108 340068
rect 395554 340054 396028 340082
rect 395068 337544 395120 337550
rect 395068 337486 395120 337492
rect 395896 337544 395948 337550
rect 395896 337486 395948 337492
rect 395436 3120 395488 3126
rect 395436 3062 395488 3068
rect 394608 3052 394660 3058
rect 394608 2994 394660 3000
rect 393608 2910 394188 2938
rect 392124 604 392176 610
rect 392124 546 392176 552
rect 393044 604 393096 610
rect 394160 592 394188 2910
rect 394160 564 394280 592
rect 393044 546 393096 552
rect 393056 480 393084 546
rect 394252 480 394280 564
rect 395448 480 395476 3062
rect 395908 2990 395936 337486
rect 396000 3330 396028 340054
rect 396092 337822 396120 340068
rect 396080 337816 396132 337822
rect 396080 337758 396132 337764
rect 396552 337754 396580 340068
rect 396540 337748 396592 337754
rect 396540 337690 396592 337696
rect 397012 337482 397040 340068
rect 397472 338026 397500 340068
rect 397460 338020 397512 338026
rect 397460 337962 397512 337968
rect 398024 337686 398052 340068
rect 398196 337816 398248 337822
rect 398196 337758 398248 337764
rect 398104 337748 398156 337754
rect 398104 337690 398156 337696
rect 397460 337680 397512 337686
rect 397460 337622 397512 337628
rect 398012 337680 398064 337686
rect 398012 337622 398064 337628
rect 397000 337476 397052 337482
rect 397000 337418 397052 337424
rect 396078 157584 396134 157593
rect 396078 157519 396080 157528
rect 396132 157519 396134 157528
rect 396080 157490 396132 157496
rect 396078 76120 396134 76129
rect 396078 76055 396080 76064
rect 396132 76055 396134 76064
rect 396080 76026 396132 76032
rect 396632 3732 396684 3738
rect 396632 3674 396684 3680
rect 395988 3324 396040 3330
rect 395988 3266 396040 3272
rect 395896 2984 395948 2990
rect 395896 2926 395948 2932
rect 396644 480 396672 3674
rect 397472 626 397500 337622
rect 398116 4010 398144 337690
rect 398104 4004 398156 4010
rect 398104 3946 398156 3952
rect 398208 2922 398236 337758
rect 398484 337346 398512 340068
rect 398944 337618 398972 340068
rect 399864 337736 399892 340190
rect 399970 340054 400168 340082
rect 399864 337708 400076 337736
rect 399484 337680 399536 337686
rect 399484 337622 399536 337628
rect 398932 337612 398984 337618
rect 398932 337554 398984 337560
rect 398472 337340 398524 337346
rect 398472 337282 398524 337288
rect 399390 76120 399446 76129
rect 399390 76055 399392 76064
rect 399444 76055 399446 76064
rect 399392 76026 399444 76032
rect 398746 16688 398802 16697
rect 398930 16688 398986 16697
rect 398802 16646 398930 16674
rect 398746 16623 398802 16632
rect 398930 16623 398986 16632
rect 399496 3806 399524 337622
rect 399484 3800 399536 3806
rect 399484 3742 399536 3748
rect 400048 3738 400076 337708
rect 400036 3732 400088 3738
rect 400036 3674 400088 3680
rect 400140 3670 400168 340054
rect 400416 337958 400444 340068
rect 400404 337952 400456 337958
rect 400404 337894 400456 337900
rect 400968 337414 400996 340068
rect 400956 337408 401008 337414
rect 400956 337350 401008 337356
rect 401428 337006 401456 340068
rect 401888 337210 401916 340068
rect 402454 340054 402836 340082
rect 402244 337408 402296 337414
rect 402244 337350 402296 337356
rect 401876 337204 401928 337210
rect 401876 337146 401928 337152
rect 401416 337000 401468 337006
rect 401416 336942 401468 336948
rect 400770 157584 400826 157593
rect 400770 157519 400772 157528
rect 400824 157519 400826 157528
rect 400772 157490 400824 157496
rect 400128 3664 400180 3670
rect 400128 3606 400180 3612
rect 402256 3602 402284 337350
rect 402244 3596 402296 3602
rect 402244 3538 402296 3544
rect 400220 3528 400272 3534
rect 400220 3470 400272 3476
rect 399024 3052 399076 3058
rect 399024 2994 399076 3000
rect 398196 2916 398248 2922
rect 398196 2858 398248 2864
rect 397472 598 397776 626
rect 397748 592 397776 598
rect 397748 564 397868 592
rect 397840 480 397868 564
rect 399036 480 399064 2994
rect 400232 480 400260 3470
rect 402808 3330 402836 340054
rect 402900 3534 402928 340068
rect 403360 338094 403388 340068
rect 403926 340054 404308 340082
rect 403348 338088 403400 338094
rect 403348 338030 403400 338036
rect 403624 338020 403676 338026
rect 403624 337962 403676 337968
rect 402888 3528 402940 3534
rect 402888 3470 402940 3476
rect 403636 3398 403664 337962
rect 404280 3942 404308 340054
rect 404372 337822 404400 340068
rect 404360 337816 404412 337822
rect 404360 337758 404412 337764
rect 404832 337686 404860 340068
rect 405398 340054 405688 340082
rect 404820 337680 404872 337686
rect 404820 337622 404872 337628
rect 405004 337000 405056 337006
rect 405004 336942 405056 336948
rect 404912 4004 404964 4010
rect 404912 3946 404964 3952
rect 404268 3936 404320 3942
rect 404268 3878 404320 3884
rect 403624 3392 403676 3398
rect 403624 3334 403676 3340
rect 402520 3324 402572 3330
rect 402520 3266 402572 3272
rect 402796 3324 402848 3330
rect 402796 3266 402848 3272
rect 401324 2984 401376 2990
rect 401324 2926 401376 2932
rect 401336 480 401364 2926
rect 402532 480 402560 3266
rect 403716 2916 403768 2922
rect 403716 2858 403768 2864
rect 403728 480 403756 2858
rect 404924 480 404952 3946
rect 405016 3126 405044 336942
rect 405660 3194 405688 340054
rect 405844 337550 405872 340068
rect 406304 338026 406332 340068
rect 406870 340054 407068 340082
rect 406292 338020 406344 338026
rect 406292 337962 406344 337968
rect 406384 337612 406436 337618
rect 406384 337554 406436 337560
rect 405832 337544 405884 337550
rect 405832 337486 405884 337492
rect 405924 337476 405976 337482
rect 405924 337418 405976 337424
rect 405648 3188 405700 3194
rect 405648 3130 405700 3136
rect 405004 3120 405056 3126
rect 405004 3062 405056 3068
rect 405936 610 405964 337418
rect 406396 3466 406424 337554
rect 407040 3874 407068 340054
rect 407316 337618 407344 340068
rect 407304 337612 407356 337618
rect 407304 337554 407356 337560
rect 407776 337074 407804 340068
rect 408342 340054 408448 340082
rect 408802 340054 409184 340082
rect 407764 337068 407816 337074
rect 407764 337010 407816 337016
rect 408420 5438 408448 340054
rect 409156 337414 409184 340054
rect 408776 337408 408828 337414
rect 408776 337350 408828 337356
rect 409144 337408 409196 337414
rect 409144 337350 409196 337356
rect 408408 5432 408460 5438
rect 408408 5374 408460 5380
rect 407028 3868 407080 3874
rect 407028 3810 407080 3816
rect 408500 3800 408552 3806
rect 408500 3742 408552 3748
rect 406384 3460 406436 3466
rect 406384 3402 406436 3408
rect 407304 3392 407356 3398
rect 407304 3334 407356 3340
rect 405924 604 405976 610
rect 405924 546 405976 552
rect 406108 604 406160 610
rect 406108 546 406160 552
rect 406120 480 406148 546
rect 407316 480 407344 3334
rect 408512 480 408540 3742
rect 408788 2938 408816 337350
rect 409144 337068 409196 337074
rect 409144 337010 409196 337016
rect 409156 3262 409184 337010
rect 409248 337006 409276 340068
rect 409236 337000 409288 337006
rect 409236 336942 409288 336948
rect 409800 3398 409828 340068
rect 410260 337754 410288 340068
rect 410734 340054 411116 340082
rect 410248 337748 410300 337754
rect 410248 337690 410300 337696
rect 411088 4010 411116 340054
rect 411272 337754 411300 340068
rect 411732 337890 411760 340068
rect 412206 340054 412496 340082
rect 411720 337884 411772 337890
rect 411720 337826 411772 337832
rect 411168 337748 411220 337754
rect 411168 337690 411220 337696
rect 411260 337748 411312 337754
rect 411260 337690 411312 337696
rect 412364 337748 412416 337754
rect 412364 337690 412416 337696
rect 411180 4078 411208 337690
rect 412376 5370 412404 337690
rect 412364 5364 412416 5370
rect 412364 5306 412416 5312
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 411076 4004 411128 4010
rect 411076 3946 411128 3952
rect 412468 3806 412496 340054
rect 412548 337884 412600 337890
rect 412548 337826 412600 337832
rect 412560 3942 412588 337826
rect 412744 337414 412772 340068
rect 413218 340054 413600 340082
rect 413284 337952 413336 337958
rect 413284 337894 413336 337900
rect 412732 337408 412784 337414
rect 412732 337350 412784 337356
rect 412548 3936 412600 3942
rect 412548 3878 412600 3884
rect 412456 3800 412508 3806
rect 412456 3742 412508 3748
rect 412088 3732 412140 3738
rect 412088 3674 412140 3680
rect 410892 3460 410944 3466
rect 410892 3402 410944 3408
rect 409788 3392 409840 3398
rect 409788 3334 409840 3340
rect 409144 3256 409196 3262
rect 409144 3198 409196 3204
rect 408788 2910 409736 2938
rect 409708 480 409736 2910
rect 410904 480 410932 3402
rect 412100 480 412128 3674
rect 413192 3664 413244 3670
rect 413192 3606 413244 3612
rect 413204 3346 413232 3606
rect 413296 3534 413324 337894
rect 413572 337736 413600 340054
rect 413664 337958 413692 340068
rect 413652 337952 413704 337958
rect 413652 337894 413704 337900
rect 414216 337754 414244 340068
rect 414676 338094 414704 340068
rect 414664 338088 414716 338094
rect 414664 338030 414716 338036
rect 414204 337748 414256 337754
rect 413572 337708 413968 337736
rect 413836 337408 413888 337414
rect 413836 337350 413888 337356
rect 413848 5302 413876 337350
rect 413836 5296 413888 5302
rect 413836 5238 413888 5244
rect 413940 3874 413968 337708
rect 414204 337690 414256 337696
rect 415136 337142 415164 340068
rect 415596 337754 415624 340068
rect 416148 337822 416176 340068
rect 416136 337816 416188 337822
rect 416136 337758 416188 337764
rect 415308 337748 415360 337754
rect 415308 337690 415360 337696
rect 415584 337748 415636 337754
rect 415584 337690 415636 337696
rect 416504 337748 416556 337754
rect 416504 337690 416556 337696
rect 415124 337136 415176 337142
rect 415124 337078 415176 337084
rect 414018 76120 414074 76129
rect 414018 76055 414020 76064
rect 414072 76055 414074 76064
rect 414020 76026 414072 76032
rect 415320 5234 415348 337690
rect 415308 5228 415360 5234
rect 415308 5170 415360 5176
rect 416516 5166 416544 337690
rect 416504 5160 416556 5166
rect 416504 5102 416556 5108
rect 413928 3868 413980 3874
rect 413928 3810 413980 3816
rect 415676 3596 415728 3602
rect 415676 3538 415728 3544
rect 413284 3528 413336 3534
rect 413284 3470 413336 3476
rect 414480 3528 414532 3534
rect 414480 3470 414532 3476
rect 413204 3318 413324 3346
rect 413296 480 413324 3318
rect 414492 480 414520 3470
rect 415688 480 415716 3538
rect 416608 2990 416636 340068
rect 416688 337816 416740 337822
rect 416688 337758 416740 337764
rect 416700 3670 416728 337758
rect 417068 337754 417096 340068
rect 417424 338020 417476 338026
rect 417424 337962 417476 337968
rect 417056 337748 417108 337754
rect 417056 337690 417108 337696
rect 416964 337204 417016 337210
rect 416964 337146 417016 337152
rect 416688 3664 416740 3670
rect 416688 3606 416740 3612
rect 416976 3346 417004 337146
rect 417436 3602 417464 337962
rect 417620 337890 417648 340068
rect 417608 337884 417660 337890
rect 417608 337826 417660 337832
rect 417976 337748 418028 337754
rect 417976 337690 418028 337696
rect 417882 157584 417938 157593
rect 417882 157519 417884 157528
rect 417936 157519 417938 157528
rect 417884 157490 417936 157496
rect 417882 63744 417938 63753
rect 417882 63679 417884 63688
rect 417936 63679 417938 63688
rect 417884 63650 417936 63656
rect 417884 40248 417936 40254
rect 417882 40216 417884 40225
rect 417936 40216 417938 40225
rect 417882 40151 417938 40160
rect 417988 5098 418016 337690
rect 417976 5092 418028 5098
rect 417976 5034 418028 5040
rect 418080 3670 418108 340068
rect 418540 336802 418568 340068
rect 419092 337074 419120 340068
rect 419080 337068 419132 337074
rect 419080 337010 419132 337016
rect 419552 336802 419580 340068
rect 420012 336870 420040 340068
rect 420276 337952 420328 337958
rect 420276 337894 420328 337900
rect 420184 337816 420236 337822
rect 420184 337758 420236 337764
rect 420000 336864 420052 336870
rect 420000 336806 420052 336812
rect 418528 336796 418580 336802
rect 418528 336738 418580 336744
rect 419448 336796 419500 336802
rect 419448 336738 419500 336744
rect 419540 336796 419592 336802
rect 419540 336738 419592 336744
rect 418158 157584 418214 157593
rect 418158 157519 418160 157528
rect 418212 157519 418214 157528
rect 418160 157490 418212 157496
rect 418158 63744 418214 63753
rect 418158 63679 418160 63688
rect 418212 63679 418214 63688
rect 418160 63650 418212 63656
rect 419460 5030 419488 336738
rect 419448 5024 419500 5030
rect 419448 4966 419500 4972
rect 420196 4010 420224 337758
rect 420184 4004 420236 4010
rect 420184 3946 420236 3952
rect 418068 3664 418120 3670
rect 418068 3606 418120 3612
rect 417424 3596 417476 3602
rect 417424 3538 417476 3544
rect 418068 3528 418120 3534
rect 418068 3470 418120 3476
rect 416976 3318 418016 3346
rect 416872 3120 416924 3126
rect 416872 3062 416924 3068
rect 416596 2984 416648 2990
rect 416596 2926 416648 2932
rect 416884 480 416912 3062
rect 417988 480 418016 3318
rect 418080 2990 418108 3470
rect 420288 3330 420316 337894
rect 420564 337482 420592 340068
rect 420552 337476 420604 337482
rect 420552 337418 420604 337424
rect 421024 337346 421052 340068
rect 421196 337408 421248 337414
rect 421196 337350 421248 337356
rect 421012 337340 421064 337346
rect 421012 337282 421064 337288
rect 420736 336864 420788 336870
rect 420736 336806 420788 336812
rect 420368 40248 420420 40254
rect 420366 40216 420368 40225
rect 420420 40216 420422 40225
rect 420366 40151 420422 40160
rect 420748 4962 420776 336806
rect 420828 336796 420880 336802
rect 420828 336738 420880 336744
rect 420736 4956 420788 4962
rect 420736 4898 420788 4904
rect 420734 3768 420790 3777
rect 420734 3703 420790 3712
rect 420748 3670 420776 3703
rect 420840 3670 420868 336738
rect 421208 336734 421236 337350
rect 421484 336802 421512 340068
rect 422036 337822 422064 340068
rect 422024 337816 422076 337822
rect 422024 337758 422076 337764
rect 421564 337136 421616 337142
rect 421564 337078 421616 337084
rect 421472 336796 421524 336802
rect 421472 336738 421524 336744
rect 421196 336728 421248 336734
rect 421196 336670 421248 336676
rect 421196 327140 421248 327146
rect 421196 327082 421248 327088
rect 421208 317422 421236 327082
rect 421196 317416 421248 317422
rect 421196 317358 421248 317364
rect 421196 307828 421248 307834
rect 421196 307770 421248 307776
rect 421208 298110 421236 307770
rect 421196 298104 421248 298110
rect 421196 298046 421248 298052
rect 421196 288448 421248 288454
rect 421196 288390 421248 288396
rect 421208 278769 421236 288390
rect 421194 278760 421250 278769
rect 421194 278695 421250 278704
rect 421378 278760 421434 278769
rect 421378 278695 421434 278704
rect 421392 269142 421420 278695
rect 421196 269136 421248 269142
rect 421196 269078 421248 269084
rect 421380 269136 421432 269142
rect 421380 269078 421432 269084
rect 421208 259457 421236 269078
rect 421194 259448 421250 259457
rect 421194 259383 421250 259392
rect 421378 259448 421434 259457
rect 421378 259383 421434 259392
rect 421392 249830 421420 259383
rect 421196 249824 421248 249830
rect 421196 249766 421248 249772
rect 421380 249824 421432 249830
rect 421380 249766 421432 249772
rect 421208 241777 421236 249766
rect 421194 241768 421250 241777
rect 421194 241703 421250 241712
rect 421194 241632 421250 241641
rect 421194 241567 421250 241576
rect 421208 240145 421236 241567
rect 421194 240136 421250 240145
rect 421194 240071 421250 240080
rect 421378 240136 421434 240145
rect 421378 240071 421434 240080
rect 421392 230518 421420 240071
rect 421196 230512 421248 230518
rect 421196 230454 421248 230460
rect 421380 230512 421432 230518
rect 421380 230454 421432 230460
rect 421208 220833 421236 230454
rect 421194 220824 421250 220833
rect 421194 220759 421250 220768
rect 421378 220824 421434 220833
rect 421378 220759 421434 220768
rect 421392 211177 421420 220759
rect 421194 211168 421250 211177
rect 421194 211103 421250 211112
rect 421378 211168 421434 211177
rect 421378 211103 421434 211112
rect 421208 201482 421236 211103
rect 421196 201476 421248 201482
rect 421196 201418 421248 201424
rect 421380 201476 421432 201482
rect 421380 201418 421432 201424
rect 421392 191865 421420 201418
rect 421194 191856 421250 191865
rect 421194 191791 421250 191800
rect 421378 191856 421434 191865
rect 421378 191791 421434 191800
rect 421208 182170 421236 191791
rect 421196 182164 421248 182170
rect 421196 182106 421248 182112
rect 421380 182164 421432 182170
rect 421380 182106 421432 182112
rect 421392 172553 421420 182106
rect 421194 172544 421250 172553
rect 421194 172479 421250 172488
rect 421378 172544 421434 172553
rect 421378 172479 421434 172488
rect 421208 162858 421236 172479
rect 421196 162852 421248 162858
rect 421196 162794 421248 162800
rect 421196 153264 421248 153270
rect 421196 153206 421248 153212
rect 421208 143546 421236 153206
rect 421196 143540 421248 143546
rect 421196 143482 421248 143488
rect 421196 133952 421248 133958
rect 421196 133894 421248 133900
rect 421208 124166 421236 133894
rect 421196 124160 421248 124166
rect 421196 124102 421248 124108
rect 421196 114572 421248 114578
rect 421196 114514 421248 114520
rect 421208 104854 421236 114514
rect 421196 104848 421248 104854
rect 421196 104790 421248 104796
rect 421196 87032 421248 87038
rect 421196 86974 421248 86980
rect 421208 85542 421236 86974
rect 421196 85536 421248 85542
rect 421196 85478 421248 85484
rect 421196 75948 421248 75954
rect 421196 75890 421248 75896
rect 421208 66230 421236 75890
rect 421196 66224 421248 66230
rect 421196 66166 421248 66172
rect 421196 56636 421248 56642
rect 421196 56578 421248 56584
rect 421208 46918 421236 56578
rect 421196 46912 421248 46918
rect 421196 46854 421248 46860
rect 421196 37324 421248 37330
rect 421196 37266 421248 37272
rect 421208 29322 421236 37266
rect 421208 29294 421328 29322
rect 421300 29050 421328 29294
rect 421208 29022 421328 29050
rect 421208 27606 421236 29022
rect 421196 27600 421248 27606
rect 421196 27542 421248 27548
rect 421380 9716 421432 9722
rect 421380 9658 421432 9664
rect 420736 3664 420788 3670
rect 420736 3606 420788 3612
rect 420828 3664 420880 3670
rect 420828 3606 420880 3612
rect 419172 3324 419224 3330
rect 419172 3266 419224 3272
rect 420276 3324 420328 3330
rect 420276 3266 420328 3272
rect 418068 2984 418120 2990
rect 418068 2926 418120 2932
rect 419184 480 419212 3266
rect 421392 2972 421420 9658
rect 421576 3058 421604 337078
rect 422496 337074 422524 340068
rect 422484 337068 422536 337074
rect 422484 337010 422536 337016
rect 422208 336796 422260 336802
rect 422208 336738 422260 336744
rect 422220 4894 422248 336738
rect 423416 335594 423444 340190
rect 423508 337278 423536 340068
rect 423496 337272 423548 337278
rect 423496 337214 423548 337220
rect 423968 336938 423996 340068
rect 424324 337680 424376 337686
rect 424324 337622 424376 337628
rect 423956 336932 424008 336938
rect 423956 336874 424008 336880
rect 423416 335566 423628 335594
rect 423404 76084 423456 76090
rect 423404 76026 423456 76032
rect 423416 75970 423444 76026
rect 423494 75984 423550 75993
rect 423416 75942 423494 75970
rect 423494 75919 423550 75928
rect 422208 4888 422260 4894
rect 422208 4830 422260 4836
rect 423600 4826 423628 335566
rect 423588 4820 423640 4826
rect 423588 4762 423640 4768
rect 424336 4010 424364 337622
rect 424416 337068 424468 337074
rect 424416 337010 424468 337016
rect 423956 4004 424008 4010
rect 423956 3946 424008 3952
rect 424324 4004 424376 4010
rect 424324 3946 424376 3952
rect 422760 3460 422812 3466
rect 422760 3402 422812 3408
rect 421564 3052 421616 3058
rect 421564 2994 421616 3000
rect 421392 2944 421512 2972
rect 421484 2938 421512 2944
rect 420368 2916 420420 2922
rect 421484 2910 421604 2938
rect 420368 2858 420420 2864
rect 420380 480 420408 2858
rect 421576 480 421604 2910
rect 422772 480 422800 3402
rect 423968 480 423996 3946
rect 424428 2922 424456 337010
rect 424888 335594 424916 340190
rect 424980 338026 425008 340068
rect 424968 338020 425020 338026
rect 424968 337962 425020 337968
rect 425440 337754 425468 340068
rect 425914 340054 426388 340082
rect 425428 337748 425480 337754
rect 425428 337690 425480 337696
rect 424888 335566 425008 335594
rect 424980 4214 425008 335566
rect 426360 5778 426388 340054
rect 426452 337686 426480 340068
rect 426440 337680 426492 337686
rect 426440 337622 426492 337628
rect 426440 337544 426492 337550
rect 426440 337486 426492 337492
rect 426452 12442 426480 337486
rect 426912 336870 426940 340068
rect 427386 340054 427768 340082
rect 427084 337612 427136 337618
rect 427084 337554 427136 337560
rect 426900 336864 426952 336870
rect 426900 336806 426952 336812
rect 426440 12436 426492 12442
rect 426440 12378 426492 12384
rect 426348 5772 426400 5778
rect 426348 5714 426400 5720
rect 424968 4208 425020 4214
rect 424968 4150 425020 4156
rect 427096 4010 427124 337554
rect 427544 12436 427596 12442
rect 427544 12378 427596 12384
rect 425152 4004 425204 4010
rect 425152 3946 425204 3952
rect 427084 4004 427136 4010
rect 427084 3946 427136 3952
rect 424416 2916 424468 2922
rect 424416 2858 424468 2864
rect 425164 480 425192 3946
rect 426348 3188 426400 3194
rect 426348 3130 426400 3136
rect 426360 480 426388 3130
rect 427556 480 427584 12378
rect 427740 5846 427768 340054
rect 427924 337618 427952 340068
rect 427912 337612 427964 337618
rect 427912 337554 427964 337560
rect 428384 337006 428412 340068
rect 428858 340054 429148 340082
rect 428464 337748 428516 337754
rect 428464 337690 428516 337696
rect 428372 337000 428424 337006
rect 428372 336942 428424 336948
rect 427728 5840 427780 5846
rect 427728 5782 427780 5788
rect 428476 3738 428504 337690
rect 429120 5982 429148 340054
rect 429396 336802 429424 340068
rect 429870 340054 430160 340082
rect 430330 340054 430436 340082
rect 429844 338088 429896 338094
rect 429844 338030 429896 338036
rect 429384 336796 429436 336802
rect 429384 336738 429436 336744
rect 429108 5976 429160 5982
rect 429108 5918 429160 5924
rect 428464 3732 428516 3738
rect 428464 3674 428516 3680
rect 429856 2990 429884 338030
rect 430132 338026 430160 340054
rect 430120 338020 430172 338026
rect 430120 337962 430172 337968
rect 430408 6118 430436 340054
rect 430868 336802 430896 340068
rect 431328 337958 431356 340068
rect 431316 337952 431368 337958
rect 431316 337894 431368 337900
rect 431224 337204 431276 337210
rect 431224 337146 431276 337152
rect 430488 336796 430540 336802
rect 430488 336738 430540 336744
rect 430856 336796 430908 336802
rect 430856 336738 430908 336744
rect 430396 6112 430448 6118
rect 430396 6054 430448 6060
rect 430500 5914 430528 336738
rect 430488 5908 430540 5914
rect 430488 5850 430540 5856
rect 431132 4004 431184 4010
rect 431132 3946 431184 3952
rect 429936 3460 429988 3466
rect 429936 3402 429988 3408
rect 428740 2984 428792 2990
rect 428740 2926 428792 2932
rect 429844 2984 429896 2990
rect 429844 2926 429896 2932
rect 428752 480 428780 2926
rect 429948 480 429976 3402
rect 431144 480 431172 3946
rect 431236 3262 431264 337146
rect 431316 337000 431368 337006
rect 431316 336942 431368 336948
rect 431224 3256 431276 3262
rect 431224 3198 431276 3204
rect 431328 3126 431356 336942
rect 431788 6866 431816 340068
rect 432340 336802 432368 340068
rect 432800 337482 432828 340068
rect 432788 337476 432840 337482
rect 432788 337418 432840 337424
rect 431868 336796 431920 336802
rect 431868 336738 431920 336744
rect 432328 336796 432380 336802
rect 432328 336738 432380 336744
rect 433156 336796 433208 336802
rect 433156 336738 433208 336744
rect 431776 6860 431828 6866
rect 431776 6802 431828 6808
rect 431880 6050 431908 336738
rect 433168 6798 433196 336738
rect 433156 6792 433208 6798
rect 433156 6734 433208 6740
rect 433260 6594 433288 340068
rect 433524 337204 433576 337210
rect 433524 337146 433576 337152
rect 433248 6588 433300 6594
rect 433248 6530 433300 6536
rect 433536 6526 433564 337146
rect 433720 336802 433748 340068
rect 434272 337210 434300 340068
rect 434260 337204 434312 337210
rect 434260 337146 434312 337152
rect 433984 337136 434036 337142
rect 433984 337078 434036 337084
rect 433708 336796 433760 336802
rect 433708 336738 433760 336744
rect 433524 6520 433576 6526
rect 433524 6462 433576 6468
rect 431868 6044 431920 6050
rect 431868 5986 431920 5992
rect 433524 5432 433576 5438
rect 433524 5374 433576 5380
rect 432328 3188 432380 3194
rect 432328 3130 432380 3136
rect 431316 3120 431368 3126
rect 431316 3062 431368 3068
rect 432340 480 432368 3130
rect 433536 480 433564 5374
rect 433996 4010 434024 337078
rect 434732 336870 434760 340068
rect 434720 336864 434772 336870
rect 434720 336806 434772 336812
rect 435192 336802 435220 340068
rect 435744 337958 435772 340068
rect 435732 337952 435784 337958
rect 435732 337894 435784 337900
rect 436008 336864 436060 336870
rect 436008 336806 436060 336812
rect 434628 336796 434680 336802
rect 434628 336738 434680 336744
rect 435180 336796 435232 336802
rect 435180 336738 435232 336744
rect 435916 336796 435968 336802
rect 435916 336738 435968 336744
rect 434640 6730 434668 336738
rect 434628 6724 434680 6730
rect 434628 6666 434680 6672
rect 435928 6526 435956 336738
rect 436020 6662 436048 336806
rect 436204 336802 436232 340068
rect 436664 337618 436692 340068
rect 436652 337612 436704 337618
rect 436652 337554 436704 337560
rect 437216 337482 437244 340068
rect 437690 340054 438072 340082
rect 438150 340054 438624 340082
rect 437480 337748 437532 337754
rect 437480 337690 437532 337696
rect 437388 337612 437440 337618
rect 437388 337554 437440 337560
rect 437204 337476 437256 337482
rect 437204 337418 437256 337424
rect 436192 336796 436244 336802
rect 436192 336738 436244 336744
rect 437296 336796 437348 336802
rect 437296 336738 437348 336744
rect 437202 157584 437258 157593
rect 437202 157519 437204 157528
rect 437256 157519 437258 157528
rect 437204 157490 437256 157496
rect 437204 87168 437256 87174
rect 437202 87136 437204 87145
rect 437256 87136 437258 87145
rect 437202 87071 437258 87080
rect 437202 76120 437258 76129
rect 437202 76055 437204 76064
rect 437256 76055 437258 76064
rect 437204 76026 437256 76032
rect 437202 63744 437258 63753
rect 437202 63679 437204 63688
rect 437256 63679 437258 63688
rect 437204 63650 437256 63656
rect 437204 40248 437256 40254
rect 437202 40216 437204 40225
rect 437256 40216 437258 40225
rect 437202 40151 437258 40160
rect 437202 29200 437258 29209
rect 437202 29135 437204 29144
rect 437256 29135 437258 29144
rect 437204 29106 437256 29112
rect 437202 16824 437258 16833
rect 437202 16759 437204 16768
rect 437256 16759 437258 16768
rect 437204 16730 437256 16736
rect 436008 6656 436060 6662
rect 436008 6598 436060 6604
rect 434628 6520 434680 6526
rect 434628 6462 434680 6468
rect 435916 6520 435968 6526
rect 435916 6462 435968 6468
rect 433984 4004 434036 4010
rect 433984 3946 434036 3952
rect 434534 3768 434590 3777
rect 434534 3703 434590 3712
rect 434548 3602 434576 3703
rect 434536 3596 434588 3602
rect 434536 3538 434588 3544
rect 434640 480 434668 6462
rect 437308 6458 437336 336738
rect 437296 6452 437348 6458
rect 437296 6394 437348 6400
rect 437400 6390 437428 337554
rect 437492 337482 437520 337690
rect 437480 337476 437532 337482
rect 437480 337418 437532 337424
rect 438044 335510 438072 340054
rect 438124 337408 438176 337414
rect 438124 337350 438176 337356
rect 438032 335504 438084 335510
rect 438032 335446 438084 335452
rect 437478 157584 437534 157593
rect 437478 157519 437480 157528
rect 437532 157519 437534 157528
rect 437480 157490 437532 157496
rect 437480 87168 437532 87174
rect 437478 87136 437480 87145
rect 437532 87136 437534 87145
rect 437478 87071 437534 87080
rect 437478 76120 437534 76129
rect 437478 76055 437480 76064
rect 437532 76055 437534 76064
rect 437480 76026 437532 76032
rect 437478 63744 437534 63753
rect 437478 63679 437480 63688
rect 437532 63679 437534 63688
rect 437480 63650 437532 63656
rect 437480 40248 437532 40254
rect 437478 40216 437480 40225
rect 437532 40216 437534 40225
rect 437478 40151 437534 40160
rect 437478 29200 437534 29209
rect 437478 29135 437480 29144
rect 437532 29135 437534 29144
rect 437480 29106 437532 29112
rect 437478 16824 437534 16833
rect 437478 16759 437480 16768
rect 437532 16759 437534 16768
rect 437480 16730 437532 16736
rect 437388 6384 437440 6390
rect 437388 6326 437440 6332
rect 437480 4140 437532 4146
rect 437480 4082 437532 4088
rect 435824 4004 435876 4010
rect 435824 3946 435876 3952
rect 435836 480 435864 3946
rect 437492 3398 437520 4082
rect 437020 3392 437072 3398
rect 437020 3334 437072 3340
rect 437480 3392 437532 3398
rect 437480 3334 437532 3340
rect 437032 480 437060 3334
rect 438136 2922 438164 337350
rect 438596 335594 438624 340054
rect 438688 337822 438716 340068
rect 438676 337816 438728 337822
rect 438676 337758 438728 337764
rect 439148 336802 439176 340068
rect 439622 340054 440096 340082
rect 439596 337544 439648 337550
rect 439596 337486 439648 337492
rect 439504 336864 439556 336870
rect 439504 336806 439556 336812
rect 439136 336796 439188 336802
rect 439136 336738 439188 336744
rect 438596 335566 438808 335594
rect 438676 335504 438728 335510
rect 438676 335446 438728 335452
rect 438688 6322 438716 335446
rect 438676 6316 438728 6322
rect 438676 6258 438728 6264
rect 438780 6254 438808 335566
rect 438768 6248 438820 6254
rect 438768 6190 438820 6196
rect 439412 4072 439464 4078
rect 439412 4014 439464 4020
rect 438216 3392 438268 3398
rect 438216 3334 438268 3340
rect 438124 2916 438176 2922
rect 438124 2858 438176 2864
rect 438228 480 438256 3334
rect 439424 480 439452 4014
rect 439516 2854 439544 336806
rect 439608 4078 439636 337486
rect 440068 7342 440096 340054
rect 440160 337414 440188 340068
rect 440148 337408 440200 337414
rect 440148 337350 440200 337356
rect 440620 336802 440648 340068
rect 441094 340054 441476 340082
rect 440148 336796 440200 336802
rect 440148 336738 440200 336744
rect 440608 336796 440660 336802
rect 440608 336738 440660 336744
rect 440056 7336 440108 7342
rect 440056 7278 440108 7284
rect 440160 6186 440188 336738
rect 441448 7410 441476 340054
rect 441632 336870 441660 340068
rect 441620 336864 441672 336870
rect 441620 336806 441672 336812
rect 442092 336802 442120 340068
rect 442566 340054 442856 340082
rect 442356 337748 442408 337754
rect 442356 337690 442408 337696
rect 442264 337476 442316 337482
rect 442264 337418 442316 337424
rect 441528 336796 441580 336802
rect 441528 336738 441580 336744
rect 442080 336796 442132 336802
rect 442080 336738 442132 336744
rect 441436 7404 441488 7410
rect 441436 7346 441488 7352
rect 440148 6180 440200 6186
rect 440148 6122 440200 6128
rect 440608 5364 440660 5370
rect 440608 5306 440660 5312
rect 439596 4072 439648 4078
rect 439596 4014 439648 4020
rect 439504 2848 439556 2854
rect 439504 2790 439556 2796
rect 440620 480 440648 5306
rect 441540 4282 441568 336738
rect 441528 4276 441580 4282
rect 441528 4218 441580 4224
rect 441804 3936 441856 3942
rect 441804 3878 441856 3884
rect 441816 480 441844 3878
rect 442276 3670 442304 337418
rect 442264 3664 442316 3670
rect 442264 3606 442316 3612
rect 442368 3262 442396 337690
rect 442828 7478 442856 340054
rect 443104 337618 443132 340068
rect 443092 337612 443144 337618
rect 443092 337554 443144 337560
rect 443564 336802 443592 340068
rect 444038 340054 444236 340082
rect 443644 336864 443696 336870
rect 443644 336806 443696 336812
rect 442908 336796 442960 336802
rect 442908 336738 442960 336744
rect 443552 336796 443604 336802
rect 443552 336738 443604 336744
rect 442816 7472 442868 7478
rect 442816 7414 442868 7420
rect 442920 4350 442948 336738
rect 442908 4344 442960 4350
rect 442908 4286 442960 4292
rect 443000 3800 443052 3806
rect 443000 3742 443052 3748
rect 442356 3256 442408 3262
rect 442356 3198 442408 3204
rect 443012 480 443040 3742
rect 443656 3398 443684 336806
rect 444208 7546 444236 340054
rect 444576 336870 444604 340068
rect 444564 336864 444616 336870
rect 444564 336806 444616 336812
rect 445036 336802 445064 340068
rect 444288 336796 444340 336802
rect 444288 336738 444340 336744
rect 445024 336796 445076 336802
rect 445024 336738 445076 336744
rect 444196 7540 444248 7546
rect 444196 7482 444248 7488
rect 444196 5296 444248 5302
rect 444196 5238 444248 5244
rect 443644 3392 443696 3398
rect 443644 3334 443696 3340
rect 444208 480 444236 5238
rect 444300 4418 444328 336738
rect 445496 8294 445524 340068
rect 446048 337822 446076 340068
rect 446036 337816 446088 337822
rect 446036 337758 446088 337764
rect 445668 336864 445720 336870
rect 445668 336806 445720 336812
rect 445576 336796 445628 336802
rect 445576 336738 445628 336744
rect 445484 8288 445536 8294
rect 445484 8230 445536 8236
rect 445588 4486 445616 336738
rect 445576 4480 445628 4486
rect 445576 4422 445628 4428
rect 444288 4412 444340 4418
rect 444288 4354 444340 4360
rect 445680 3874 445708 336806
rect 446508 336802 446536 340068
rect 446496 336796 446548 336802
rect 446496 336738 446548 336744
rect 446968 8226 446996 340068
rect 447520 336802 447548 340068
rect 447994 340054 448376 340082
rect 447048 336796 447100 336802
rect 447048 336738 447100 336744
rect 447508 336796 447560 336802
rect 447508 336738 447560 336744
rect 448244 336796 448296 336802
rect 448244 336738 448296 336744
rect 446956 8220 447008 8226
rect 446956 8162 447008 8168
rect 447060 4554 447088 336738
rect 448256 8158 448284 336738
rect 448244 8152 448296 8158
rect 448244 8094 448296 8100
rect 447784 5228 447836 5234
rect 447784 5170 447836 5176
rect 447048 4548 447100 4554
rect 447048 4490 447100 4496
rect 445392 3868 445444 3874
rect 445392 3810 445444 3816
rect 445668 3868 445720 3874
rect 445668 3810 445720 3816
rect 445404 480 445432 3810
rect 446588 3324 446640 3330
rect 446588 3266 446640 3272
rect 446600 480 446628 3266
rect 447796 480 447824 5170
rect 448348 4622 448376 340054
rect 448440 336802 448468 340068
rect 448992 337618 449020 340068
rect 449466 340054 449848 340082
rect 448980 337612 449032 337618
rect 448980 337554 449032 337560
rect 449164 337476 449216 337482
rect 449164 337418 449216 337424
rect 448428 336796 448480 336802
rect 448428 336738 448480 336744
rect 448428 336660 448480 336666
rect 448428 336602 448480 336608
rect 448336 4616 448388 4622
rect 448336 4558 448388 4564
rect 448440 4078 448468 336602
rect 448428 4072 448480 4078
rect 448428 4014 448480 4020
rect 448980 2984 449032 2990
rect 448980 2926 449032 2932
rect 448992 480 449020 2926
rect 449176 2922 449204 337418
rect 449820 4690 449848 340054
rect 449912 336802 449940 340068
rect 450464 336870 450492 340068
rect 450938 340054 451136 340082
rect 450452 336864 450504 336870
rect 450452 336806 450504 336812
rect 449900 336796 449952 336802
rect 449900 336738 449952 336744
rect 451004 336796 451056 336802
rect 451004 336738 451056 336744
rect 451016 8090 451044 336738
rect 451004 8084 451056 8090
rect 451004 8026 451056 8032
rect 451108 4758 451136 340054
rect 451188 336864 451240 336870
rect 451188 336806 451240 336812
rect 451096 4752 451148 4758
rect 451096 4694 451148 4700
rect 449808 4684 449860 4690
rect 449808 4626 449860 4632
rect 451200 3738 451228 336806
rect 451384 336802 451412 340068
rect 451844 337958 451872 340068
rect 452410 340054 452608 340082
rect 451832 337952 451884 337958
rect 451832 337894 451884 337900
rect 451372 336796 451424 336802
rect 451372 336738 451424 336744
rect 452476 336796 452528 336802
rect 452476 336738 452528 336744
rect 452488 8022 452516 336738
rect 452476 8016 452528 8022
rect 452476 7958 452528 7964
rect 452580 5506 452608 340054
rect 452856 336802 452884 340068
rect 453316 336870 453344 340068
rect 453304 336864 453356 336870
rect 453304 336806 453356 336812
rect 452844 336796 452896 336802
rect 452844 336738 452896 336744
rect 453764 336796 453816 336802
rect 453764 336738 453816 336744
rect 453776 7954 453804 336738
rect 453764 7948 453816 7954
rect 453764 7890 453816 7896
rect 452568 5500 452620 5506
rect 452568 5442 452620 5448
rect 453868 5438 453896 340068
rect 453948 336864 454000 336870
rect 453948 336806 454000 336812
rect 453856 5432 453908 5438
rect 453856 5374 453908 5380
rect 451280 5160 451332 5166
rect 451280 5102 451332 5108
rect 451188 3732 451240 3738
rect 451188 3674 451240 3680
rect 450176 3052 450228 3058
rect 450176 2994 450228 3000
rect 449164 2916 449216 2922
rect 449164 2858 449216 2864
rect 450188 480 450216 2994
rect 451292 480 451320 5102
rect 453960 3942 453988 336806
rect 454328 336802 454356 340068
rect 454788 338026 454816 340068
rect 454776 338020 454828 338026
rect 454776 337962 454828 337968
rect 454316 336796 454368 336802
rect 454316 336738 454368 336744
rect 455236 336796 455288 336802
rect 455236 336738 455288 336744
rect 454040 87304 454092 87310
rect 454038 87272 454040 87281
rect 454092 87272 454094 87281
rect 454038 87207 454094 87216
rect 455248 7886 455276 336738
rect 455236 7880 455288 7886
rect 455236 7822 455288 7828
rect 455340 5370 455368 340068
rect 455696 337816 455748 337822
rect 455694 337784 455696 337793
rect 455748 337784 455750 337793
rect 455694 337719 455750 337728
rect 455604 337680 455656 337686
rect 455604 337622 455656 337628
rect 455328 5364 455380 5370
rect 455328 5306 455380 5312
rect 454868 5092 454920 5098
rect 454868 5034 454920 5040
rect 453672 3936 453724 3942
rect 453672 3878 453724 3884
rect 453948 3936 454000 3942
rect 453948 3878 454000 3884
rect 452476 604 452528 610
rect 452476 546 452528 552
rect 452488 480 452516 546
rect 453684 480 453712 3878
rect 454880 480 454908 5034
rect 455616 1442 455644 337622
rect 455800 336802 455828 340068
rect 456274 340054 456748 340082
rect 455788 336796 455840 336802
rect 455788 336738 455840 336744
rect 456616 336796 456668 336802
rect 456616 336738 456668 336744
rect 456522 157584 456578 157593
rect 456522 157519 456524 157528
rect 456576 157519 456578 157528
rect 456524 157490 456576 157496
rect 456522 63744 456578 63753
rect 456522 63679 456524 63688
rect 456576 63679 456578 63688
rect 456524 63650 456576 63656
rect 456524 40248 456576 40254
rect 456522 40216 456524 40225
rect 456576 40216 456578 40225
rect 456522 40151 456578 40160
rect 456522 29200 456578 29209
rect 456522 29135 456524 29144
rect 456576 29135 456578 29144
rect 456524 29106 456576 29112
rect 456522 16960 456578 16969
rect 456522 16895 456524 16904
rect 456576 16895 456578 16904
rect 456524 16866 456576 16872
rect 456628 7818 456656 336738
rect 456616 7812 456668 7818
rect 456616 7754 456668 7760
rect 456720 3874 456748 340054
rect 456812 336870 456840 340068
rect 456800 336864 456852 336870
rect 456800 336806 456852 336812
rect 457272 336802 457300 340068
rect 457732 337686 457760 340068
rect 457720 337680 457772 337686
rect 457720 337622 457772 337628
rect 458088 336864 458140 336870
rect 458088 336806 458140 336812
rect 457260 336796 457312 336802
rect 457260 336738 457312 336744
rect 457996 336796 458048 336802
rect 457996 336738 458048 336744
rect 456984 87304 457036 87310
rect 456982 87272 456984 87281
rect 457036 87272 457038 87281
rect 456982 87207 457038 87216
rect 456890 63744 456946 63753
rect 456890 63679 456892 63688
rect 456944 63679 456946 63688
rect 456892 63650 456944 63656
rect 456892 40248 456944 40254
rect 456890 40216 456892 40225
rect 456944 40216 456946 40225
rect 456890 40151 456946 40160
rect 456798 29200 456854 29209
rect 456798 29135 456800 29144
rect 456852 29135 456854 29144
rect 456800 29106 456852 29112
rect 457444 16924 457496 16930
rect 457444 16866 457496 16872
rect 457456 16833 457484 16866
rect 457442 16824 457498 16833
rect 457442 16759 457498 16768
rect 458008 7750 458036 336738
rect 457996 7744 458048 7750
rect 457996 7686 458048 7692
rect 458100 5098 458128 336806
rect 458284 336802 458312 340068
rect 458758 340054 459048 340082
rect 458272 336796 458324 336802
rect 458272 336738 458324 336744
rect 459020 335594 459048 340054
rect 459204 337278 459232 340068
rect 459756 338026 459784 340068
rect 459744 338020 459796 338026
rect 459744 337962 459796 337968
rect 459192 337272 459244 337278
rect 459192 337214 459244 337220
rect 460296 337272 460348 337278
rect 460296 337214 460348 337220
rect 459652 336864 459704 336870
rect 459652 336806 459704 336812
rect 459468 336796 459520 336802
rect 459468 336738 459520 336744
rect 459020 335566 459416 335594
rect 458270 157584 458326 157593
rect 458270 157519 458272 157528
rect 458324 157519 458326 157528
rect 458272 157490 458324 157496
rect 459388 7682 459416 335566
rect 459376 7676 459428 7682
rect 459376 7618 459428 7624
rect 459480 5302 459508 336738
rect 459664 331226 459692 336806
rect 459652 331220 459704 331226
rect 459652 331162 459704 331168
rect 460112 331220 460164 331226
rect 460112 331162 460164 331168
rect 460124 323626 460152 331162
rect 460032 323598 460152 323626
rect 460032 318889 460060 323598
rect 460018 318880 460074 318889
rect 460018 318815 460074 318824
rect 460202 318880 460258 318889
rect 460202 318815 460258 318824
rect 460216 317422 460244 318815
rect 460204 317416 460256 317422
rect 460204 317358 460256 317364
rect 460204 307828 460256 307834
rect 460204 307770 460256 307776
rect 460216 302410 460244 307770
rect 460124 302382 460244 302410
rect 460124 299554 460152 302382
rect 460032 299526 460152 299554
rect 460032 298110 460060 299526
rect 460020 298104 460072 298110
rect 460020 298046 460072 298052
rect 460112 288448 460164 288454
rect 460112 288390 460164 288396
rect 460124 283014 460152 288390
rect 460112 283008 460164 283014
rect 460112 282950 460164 282956
rect 460112 282804 460164 282810
rect 460112 282746 460164 282752
rect 460124 280158 460152 282746
rect 460112 280152 460164 280158
rect 460112 280094 460164 280100
rect 460112 273148 460164 273154
rect 460112 273090 460164 273096
rect 460124 270502 460152 273090
rect 460112 270496 460164 270502
rect 460112 270438 460164 270444
rect 460020 260976 460072 260982
rect 460020 260918 460072 260924
rect 460032 260846 460060 260918
rect 460020 260840 460072 260846
rect 460020 260782 460072 260788
rect 460204 260840 460256 260846
rect 460204 260782 460256 260788
rect 460216 253858 460244 260782
rect 460124 253830 460244 253858
rect 460124 244390 460152 253830
rect 460112 244384 460164 244390
rect 460112 244326 460164 244332
rect 460020 244248 460072 244254
rect 460020 244190 460072 244196
rect 460032 240145 460060 244190
rect 459834 240136 459890 240145
rect 459834 240071 459890 240080
rect 460018 240136 460074 240145
rect 460018 240071 460074 240080
rect 459848 230518 459876 240071
rect 459836 230512 459888 230518
rect 459836 230454 459888 230460
rect 460112 230512 460164 230518
rect 460112 230454 460164 230460
rect 460124 225078 460152 230454
rect 460112 225072 460164 225078
rect 460112 225014 460164 225020
rect 460020 224936 460072 224942
rect 460020 224878 460072 224884
rect 460032 220833 460060 224878
rect 459834 220824 459890 220833
rect 459834 220759 459890 220768
rect 460018 220824 460074 220833
rect 460018 220759 460074 220768
rect 459848 215286 459876 220759
rect 459836 215280 459888 215286
rect 459836 215222 459888 215228
rect 460020 215280 460072 215286
rect 460020 215222 460072 215228
rect 460032 211154 460060 215222
rect 460032 211126 460152 211154
rect 460124 205766 460152 211126
rect 460112 205760 460164 205766
rect 460112 205702 460164 205708
rect 460020 205624 460072 205630
rect 460020 205566 460072 205572
rect 460032 196042 460060 205566
rect 460020 196036 460072 196042
rect 460020 195978 460072 195984
rect 460112 195900 460164 195906
rect 460112 195842 460164 195848
rect 460124 193202 460152 195842
rect 460032 193174 460152 193202
rect 460032 186386 460060 193174
rect 460020 186380 460072 186386
rect 460020 186322 460072 186328
rect 460112 186312 460164 186318
rect 460112 186254 460164 186260
rect 460124 183530 460152 186254
rect 460112 183524 460164 183530
rect 460112 183466 460164 183472
rect 460112 176520 460164 176526
rect 460112 176462 460164 176468
rect 460124 167006 460152 176462
rect 460112 167000 460164 167006
rect 460112 166942 460164 166948
rect 460112 161492 460164 161498
rect 460112 161434 460164 161440
rect 460124 151774 460152 161434
rect 460112 151768 460164 151774
rect 460112 151710 460164 151716
rect 460112 142248 460164 142254
rect 460112 142190 460164 142196
rect 460124 142118 460152 142190
rect 460112 142112 460164 142118
rect 460112 142054 460164 142060
rect 460204 132524 460256 132530
rect 460204 132466 460256 132472
rect 460216 124098 460244 132466
rect 460020 124092 460072 124098
rect 460020 124034 460072 124040
rect 460204 124092 460256 124098
rect 460204 124034 460256 124040
rect 460032 108882 460060 124034
rect 460032 108854 460152 108882
rect 460124 99482 460152 108854
rect 460112 99476 460164 99482
rect 460112 99418 460164 99424
rect 460112 99340 460164 99346
rect 460112 99282 460164 99288
rect 460124 80186 460152 99282
rect 460032 80158 460152 80186
rect 460032 70530 460060 80158
rect 460032 70502 460152 70530
rect 460124 70258 460152 70502
rect 459940 70230 460152 70258
rect 459940 67590 459968 70230
rect 459928 67584 459980 67590
rect 459928 67526 459980 67532
rect 460204 67584 460256 67590
rect 460204 67526 460256 67532
rect 460216 58018 460244 67526
rect 460124 57990 460244 58018
rect 460124 57934 460152 57990
rect 460112 57928 460164 57934
rect 460112 57870 460164 57876
rect 460020 48340 460072 48346
rect 460020 48282 460072 48288
rect 460032 48210 460060 48282
rect 460020 48204 460072 48210
rect 460020 48146 460072 48152
rect 460204 41404 460256 41410
rect 460204 41346 460256 41352
rect 460216 31770 460244 41346
rect 460032 31742 460244 31770
rect 460032 31634 460060 31742
rect 460032 31606 460152 31634
rect 460124 12458 460152 31606
rect 460032 12430 460152 12458
rect 459468 5296 459520 5302
rect 459468 5238 459520 5244
rect 458088 5092 458140 5098
rect 458088 5034 458140 5040
rect 458456 5024 458508 5030
rect 458456 4966 458508 4972
rect 456708 3868 456760 3874
rect 456708 3810 456760 3816
rect 457260 2168 457312 2174
rect 457260 2110 457312 2116
rect 455616 1414 456104 1442
rect 456076 480 456104 1414
rect 457272 480 457300 2110
rect 458468 480 458496 4966
rect 460032 3806 460060 12430
rect 459652 3800 459704 3806
rect 459652 3742 459704 3748
rect 460020 3800 460072 3806
rect 460020 3742 460072 3748
rect 459664 480 459692 3742
rect 460308 2922 460336 337214
rect 460584 335594 460612 340190
rect 460676 337890 460704 340068
rect 460848 338020 460900 338026
rect 460848 337962 460900 337968
rect 460664 337884 460716 337890
rect 460664 337826 460716 337832
rect 460584 335566 460796 335594
rect 460768 7614 460796 335566
rect 460756 7608 460808 7614
rect 460756 7550 460808 7556
rect 460860 5234 460888 337962
rect 461228 336802 461256 340068
rect 461702 340054 461992 340082
rect 462162 340054 462268 340082
rect 461216 336796 461268 336802
rect 461216 336738 461268 336744
rect 461964 336734 461992 340054
rect 462136 336796 462188 336802
rect 462136 336738 462188 336744
rect 461952 336728 462004 336734
rect 461952 336670 462004 336676
rect 460848 5228 460900 5234
rect 460848 5170 460900 5176
rect 462044 5024 462096 5030
rect 462044 4966 462096 4972
rect 460848 3528 460900 3534
rect 460848 3470 460900 3476
rect 460296 2916 460348 2922
rect 460296 2858 460348 2864
rect 460860 480 460888 3470
rect 462056 480 462084 4966
rect 462148 4826 462176 336738
rect 462136 4820 462188 4826
rect 462136 4762 462188 4768
rect 462240 3534 462268 340054
rect 462700 336802 462728 340068
rect 463174 340054 463556 340082
rect 463528 336954 463556 340054
rect 463620 337958 463648 340068
rect 463608 337952 463660 337958
rect 463608 337894 463660 337900
rect 463606 337784 463662 337793
rect 463606 337719 463662 337728
rect 463620 337550 463648 337719
rect 463608 337544 463660 337550
rect 463608 337486 463660 337492
rect 463528 336926 463648 336954
rect 462688 336796 462740 336802
rect 462688 336738 462740 336744
rect 463516 336796 463568 336802
rect 463516 336738 463568 336744
rect 463528 5166 463556 336738
rect 463516 5160 463568 5166
rect 463516 5102 463568 5108
rect 463240 3800 463292 3806
rect 463240 3742 463292 3748
rect 462228 3528 462280 3534
rect 462228 3470 462280 3476
rect 463252 480 463280 3742
rect 463620 3670 463648 336926
rect 463792 336864 463844 336870
rect 463792 336806 463844 336812
rect 463804 321586 463832 336806
rect 464172 336802 464200 340068
rect 464632 337346 464660 340068
rect 465106 340054 465488 340082
rect 465658 340054 465948 340082
rect 466118 340054 466316 340082
rect 464620 337340 464672 337346
rect 464620 337282 464672 337288
rect 464160 336796 464212 336802
rect 464160 336738 464212 336744
rect 464988 336796 465040 336802
rect 464988 336738 465040 336744
rect 463712 321558 463832 321586
rect 463712 316010 463740 321558
rect 463712 315982 463924 316010
rect 463896 306406 463924 315982
rect 463700 306400 463752 306406
rect 463700 306342 463752 306348
rect 463884 306400 463936 306406
rect 463884 306342 463936 306348
rect 463712 302138 463740 306342
rect 463712 302110 463832 302138
rect 463804 292618 463832 302110
rect 463804 292590 463924 292618
rect 463896 292482 463924 292590
rect 463804 292454 463924 292482
rect 463804 282962 463832 292454
rect 463712 282934 463832 282962
rect 463712 282826 463740 282934
rect 463712 282798 463832 282826
rect 463804 275330 463832 282798
rect 463792 275324 463844 275330
rect 463792 275266 463844 275272
rect 463884 270564 463936 270570
rect 463884 270506 463936 270512
rect 463896 263514 463924 270506
rect 463804 263486 463924 263514
rect 463804 260846 463832 263486
rect 463792 260840 463844 260846
rect 463792 260782 463844 260788
rect 463700 251252 463752 251258
rect 463700 251194 463752 251200
rect 463712 244202 463740 251194
rect 463712 244174 463832 244202
rect 463804 234682 463832 244174
rect 463804 234654 464016 234682
rect 463988 231849 464016 234654
rect 463790 231840 463846 231849
rect 463790 231775 463846 231784
rect 463974 231840 464030 231849
rect 463974 231775 464030 231784
rect 463804 222222 463832 231775
rect 463792 222216 463844 222222
rect 463792 222158 463844 222164
rect 464068 222216 464120 222222
rect 464068 222158 464120 222164
rect 464080 215422 464108 222158
rect 464068 215416 464120 215422
rect 464068 215358 464120 215364
rect 463976 215280 464028 215286
rect 463976 215222 464028 215228
rect 463988 212537 464016 215222
rect 463790 212528 463846 212537
rect 463790 212463 463846 212472
rect 463974 212528 464030 212537
rect 463974 212463 464030 212472
rect 463804 202910 463832 212463
rect 463792 202904 463844 202910
rect 463792 202846 463844 202852
rect 464068 202904 464120 202910
rect 464068 202846 464120 202852
rect 464080 196110 464108 202846
rect 464068 196104 464120 196110
rect 464068 196046 464120 196052
rect 463976 195968 464028 195974
rect 463976 195910 464028 195916
rect 463988 193225 464016 195910
rect 463790 193216 463846 193225
rect 463790 193151 463846 193160
rect 463974 193216 464030 193225
rect 463974 193151 464030 193160
rect 463804 183598 463832 193151
rect 463792 183592 463844 183598
rect 463792 183534 463844 183540
rect 464068 183592 464120 183598
rect 464068 183534 464120 183540
rect 464080 176730 464108 183534
rect 463884 176724 463936 176730
rect 463884 176666 463936 176672
rect 464068 176724 464120 176730
rect 464068 176666 464120 176672
rect 463896 157434 463924 176666
rect 463712 157406 463924 157434
rect 463712 157298 463740 157406
rect 463712 157270 463832 157298
rect 463804 147762 463832 157270
rect 463792 147756 463844 147762
rect 463792 147698 463844 147704
rect 463700 144968 463752 144974
rect 463700 144910 463752 144916
rect 463712 138038 463740 144910
rect 463700 138032 463752 138038
rect 463700 137974 463752 137980
rect 463884 137964 463936 137970
rect 463884 137906 463936 137912
rect 463896 132530 463924 137906
rect 463700 132524 463752 132530
rect 463700 132466 463752 132472
rect 463884 132524 463936 132530
rect 463884 132466 463936 132472
rect 463712 132410 463740 132466
rect 463712 132382 463832 132410
rect 463804 122890 463832 132382
rect 463804 122862 463924 122890
rect 463896 111110 463924 122862
rect 463884 111104 463936 111110
rect 463884 111046 463936 111052
rect 464068 111104 464120 111110
rect 464068 111046 464120 111052
rect 464080 106321 464108 111046
rect 463882 106312 463938 106321
rect 463882 106247 463938 106256
rect 464066 106312 464122 106321
rect 464066 106247 464122 106256
rect 463896 99006 463924 106247
rect 463700 99000 463752 99006
rect 463700 98942 463752 98948
rect 463884 99000 463936 99006
rect 463884 98942 463936 98948
rect 463712 89706 463740 98942
rect 463712 89678 463832 89706
rect 463804 89570 463832 89678
rect 463804 89542 463924 89570
rect 463896 70530 463924 89542
rect 463804 70502 463924 70530
rect 463804 70394 463832 70502
rect 463712 70366 463832 70394
rect 463608 3664 463660 3670
rect 463608 3606 463660 3612
rect 463712 610 463740 70366
rect 465000 5098 465028 336738
rect 465460 335646 465488 340054
rect 465448 335640 465500 335646
rect 465448 335582 465500 335588
rect 465920 333010 465948 340054
rect 465920 332982 466224 333010
rect 466090 87544 466146 87553
rect 466090 87479 466146 87488
rect 466104 87145 466132 87479
rect 466090 87136 466146 87145
rect 466090 87071 466146 87080
rect 466090 76528 466146 76537
rect 466090 76463 466146 76472
rect 466104 76129 466132 76463
rect 466090 76120 466146 76129
rect 466090 76055 466146 76064
rect 464988 5092 465040 5098
rect 464988 5034 465040 5040
rect 465632 5024 465684 5030
rect 465632 4966 465684 4972
rect 463700 604 463752 610
rect 463700 546 463752 552
rect 464436 604 464488 610
rect 464436 546 464488 552
rect 464448 480 464476 546
rect 465644 480 465672 4966
rect 466196 4962 466224 332982
rect 466184 4956 466236 4962
rect 466184 4898 466236 4904
rect 466288 3534 466316 340054
rect 466564 337346 466592 340068
rect 467116 337958 467144 340068
rect 467104 337952 467156 337958
rect 467104 337894 467156 337900
rect 467576 337385 467604 340068
rect 468036 337958 468064 340068
rect 468602 340054 468984 340082
rect 467748 337952 467800 337958
rect 467748 337894 467800 337900
rect 468024 337952 468076 337958
rect 468024 337894 468076 337900
rect 467562 337376 467618 337385
rect 466552 337340 466604 337346
rect 467562 337311 467618 337320
rect 466552 337282 466604 337288
rect 466368 335640 466420 335646
rect 466368 335582 466420 335588
rect 466380 3602 466408 335582
rect 467760 4865 467788 337894
rect 468760 8356 468812 8362
rect 468760 8298 468812 8304
rect 467746 4856 467802 4865
rect 467746 4791 467802 4800
rect 466368 3596 466420 3602
rect 466368 3538 466420 3544
rect 466276 3528 466328 3534
rect 466276 3470 466328 3476
rect 467932 3460 467984 3466
rect 467932 3402 467984 3408
rect 466828 2848 466880 2854
rect 466828 2790 466880 2796
rect 466840 480 466868 2790
rect 467944 480 467972 3402
rect 468772 3369 468800 8298
rect 468956 5574 468984 340054
rect 469048 8362 469076 340068
rect 469128 337952 469180 337958
rect 469128 337894 469180 337900
rect 469036 8356 469088 8362
rect 469036 8298 469088 8304
rect 469140 7970 469168 337894
rect 469508 337278 469536 340068
rect 469496 337272 469548 337278
rect 469496 337214 469548 337220
rect 469220 336932 469272 336938
rect 469220 336874 469272 336880
rect 469048 7942 469168 7970
rect 468944 5568 468996 5574
rect 468944 5510 468996 5516
rect 469048 3466 469076 7942
rect 469128 4888 469180 4894
rect 469128 4830 469180 4836
rect 469036 3460 469088 3466
rect 469036 3402 469088 3408
rect 468758 3360 468814 3369
rect 468758 3295 468814 3304
rect 469140 480 469168 4830
rect 469232 1442 469260 336874
rect 469876 182170 469904 581062
rect 469956 580304 470008 580310
rect 469956 580246 470008 580252
rect 469968 252550 469996 580246
rect 470060 299470 470088 581130
rect 470140 579216 470192 579222
rect 470140 579158 470192 579164
rect 470152 322930 470180 579158
rect 470244 346390 470272 581198
rect 470336 393310 470364 581266
rect 470428 416770 470456 581334
rect 470520 440230 470548 581402
rect 471244 579284 471296 579290
rect 471244 579226 471296 579232
rect 470508 440224 470560 440230
rect 470508 440166 470560 440172
rect 470416 416764 470468 416770
rect 470416 416706 470468 416712
rect 471256 405686 471284 579226
rect 471348 499526 471376 583578
rect 471440 546446 471468 583646
rect 580632 583568 580684 583574
rect 580632 583510 580684 583516
rect 580448 583500 580500 583506
rect 580448 583442 580500 583448
rect 580264 583432 580316 583438
rect 580264 583374 580316 583380
rect 580080 581052 580132 581058
rect 580080 580994 580132 581000
rect 580092 580122 580120 580994
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 580242 580212 580751
rect 580172 580236 580224 580242
rect 580172 580178 580224 580184
rect 580092 580094 580212 580122
rect 579804 579148 579856 579154
rect 579804 579090 579856 579096
rect 579712 557524 579764 557530
rect 579712 557466 579764 557472
rect 579724 557297 579752 557466
rect 579710 557288 579766 557297
rect 579710 557223 579766 557232
rect 471428 546440 471480 546446
rect 471428 546382 471480 546388
rect 579712 546440 579764 546446
rect 579712 546382 579764 546388
rect 579724 545601 579752 546382
rect 579710 545592 579766 545601
rect 579710 545527 579766 545536
rect 579712 510604 579764 510610
rect 579712 510546 579764 510552
rect 579724 510377 579752 510546
rect 579710 510368 579766 510377
rect 579710 510303 579766 510312
rect 471336 499520 471388 499526
rect 471336 499462 471388 499468
rect 579712 499520 579764 499526
rect 579712 499462 579764 499468
rect 579724 498681 579752 499462
rect 579710 498672 579766 498681
rect 579710 498607 579766 498616
rect 579712 463684 579764 463690
rect 579712 463626 579764 463632
rect 579724 463457 579752 463626
rect 579710 463448 579766 463457
rect 579710 463383 579766 463392
rect 579816 451761 579844 579090
rect 579988 579080 580040 579086
rect 579988 579022 580040 579028
rect 579896 579012 579948 579018
rect 579896 578954 579948 578960
rect 579802 451752 579858 451761
rect 579802 451687 579858 451696
rect 579804 440224 579856 440230
rect 579804 440166 579856 440172
rect 579816 439929 579844 440166
rect 579802 439920 579858 439929
rect 579802 439855 579858 439864
rect 579804 416764 579856 416770
rect 579804 416706 579856 416712
rect 579816 416537 579844 416706
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 471244 405680 471296 405686
rect 471244 405622 471296 405628
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404841 579844 405622
rect 579802 404832 579858 404841
rect 579802 404767 579858 404776
rect 470324 393304 470376 393310
rect 470324 393246 470376 393252
rect 579804 393304 579856 393310
rect 579804 393246 579856 393252
rect 579816 393009 579844 393246
rect 579802 393000 579858 393009
rect 579802 392935 579858 392944
rect 579908 369617 579936 578954
rect 579894 369608 579950 369617
rect 579894 369543 579950 369552
rect 580000 357921 580028 579022
rect 580080 578944 580132 578950
rect 580080 578886 580132 578892
rect 579986 357912 580042 357921
rect 579986 357847 580042 357856
rect 470232 346384 470284 346390
rect 470232 346326 470284 346332
rect 579988 346384 580040 346390
rect 579988 346326 580040 346332
rect 580000 346089 580028 346326
rect 579986 346080 580042 346089
rect 579986 346015 580042 346024
rect 483020 338088 483072 338094
rect 483018 338056 483020 338065
rect 483388 338088 483440 338094
rect 483072 338056 483074 338065
rect 483018 337991 483074 338000
rect 483386 338056 483388 338065
rect 499580 338088 499632 338094
rect 483440 338056 483442 338065
rect 499580 338030 499632 338036
rect 483386 337991 483442 338000
rect 483018 337920 483074 337929
rect 483018 337855 483020 337864
rect 483072 337855 483074 337864
rect 483386 337920 483442 337929
rect 483386 337855 483388 337864
rect 483020 337826 483072 337832
rect 483440 337855 483442 337864
rect 483388 337826 483440 337832
rect 483018 337784 483074 337793
rect 483018 337719 483020 337728
rect 483072 337719 483074 337728
rect 483386 337784 483442 337793
rect 483386 337719 483388 337728
rect 483020 337690 483072 337696
rect 483440 337719 483442 337728
rect 483388 337690 483440 337696
rect 483018 337648 483074 337657
rect 483018 337583 483020 337592
rect 483072 337583 483074 337592
rect 483478 337648 483534 337657
rect 483478 337583 483480 337592
rect 483020 337554 483072 337560
rect 483532 337583 483534 337592
rect 483480 337554 483532 337560
rect 483112 337544 483164 337550
rect 483296 337544 483348 337550
rect 483164 337492 483296 337498
rect 483112 337486 483348 337492
rect 483124 337470 483336 337486
rect 492680 337204 492732 337210
rect 492680 337146 492732 337152
rect 485780 337136 485832 337142
rect 485780 337078 485832 337084
rect 477592 337068 477644 337074
rect 477592 337010 477644 337016
rect 475384 337000 475436 337006
rect 475384 336942 475436 336948
rect 470600 336864 470652 336870
rect 470600 336806 470652 336812
rect 470612 328438 470640 336806
rect 470600 328432 470652 328438
rect 470600 328374 470652 328380
rect 470140 322924 470192 322930
rect 470140 322866 470192 322872
rect 470600 318844 470652 318850
rect 470600 318786 470652 318792
rect 470612 309126 470640 318786
rect 470600 309120 470652 309126
rect 470600 309062 470652 309068
rect 470600 299532 470652 299538
rect 470600 299474 470652 299480
rect 470048 299464 470100 299470
rect 470048 299406 470100 299412
rect 470612 289814 470640 299474
rect 470600 289808 470652 289814
rect 470600 289750 470652 289756
rect 470600 280220 470652 280226
rect 470600 280162 470652 280168
rect 470612 270502 470640 280162
rect 470600 270496 470652 270502
rect 470600 270438 470652 270444
rect 470600 260908 470652 260914
rect 470600 260850 470652 260856
rect 469956 252544 470008 252550
rect 469956 252486 470008 252492
rect 470612 251190 470640 260850
rect 470600 251184 470652 251190
rect 470600 251126 470652 251132
rect 470600 241528 470652 241534
rect 470600 241470 470652 241476
rect 470612 231849 470640 241470
rect 470414 231840 470470 231849
rect 470414 231775 470470 231784
rect 470598 231840 470654 231849
rect 470598 231775 470654 231784
rect 470428 222222 470456 231775
rect 470416 222216 470468 222222
rect 470416 222158 470468 222164
rect 470600 222216 470652 222222
rect 470600 222158 470652 222164
rect 470612 212537 470640 222158
rect 470414 212528 470470 212537
rect 470414 212463 470470 212472
rect 470598 212528 470654 212537
rect 470598 212463 470654 212472
rect 470428 202910 470456 212463
rect 470416 202904 470468 202910
rect 470416 202846 470468 202852
rect 470600 202904 470652 202910
rect 470600 202846 470652 202852
rect 470612 193225 470640 202846
rect 470414 193216 470470 193225
rect 470414 193151 470470 193160
rect 470598 193216 470654 193225
rect 470598 193151 470654 193160
rect 470428 183598 470456 193151
rect 470416 183592 470468 183598
rect 470416 183534 470468 183540
rect 470600 183592 470652 183598
rect 470600 183534 470652 183540
rect 469864 182164 469916 182170
rect 469864 182106 469916 182112
rect 470612 173913 470640 183534
rect 470414 173904 470470 173913
rect 470414 173839 470470 173848
rect 470598 173904 470654 173913
rect 470598 173839 470654 173848
rect 470428 164257 470456 173839
rect 470414 164248 470470 164257
rect 470414 164183 470470 164192
rect 470598 164248 470654 164257
rect 470598 164183 470654 164192
rect 470612 154562 470640 164183
rect 470416 154556 470468 154562
rect 470416 154498 470468 154504
rect 470600 154556 470652 154562
rect 470600 154498 470652 154504
rect 470428 144945 470456 154498
rect 470414 144936 470470 144945
rect 470414 144871 470470 144880
rect 470598 144936 470654 144945
rect 470598 144871 470654 144880
rect 470612 135250 470640 144871
rect 470416 135244 470468 135250
rect 470416 135186 470468 135192
rect 470600 135244 470652 135250
rect 470600 135186 470652 135192
rect 470428 125633 470456 135186
rect 470414 125624 470470 125633
rect 470414 125559 470470 125568
rect 470598 125624 470654 125633
rect 470598 125559 470654 125568
rect 470612 115938 470640 125559
rect 470600 115932 470652 115938
rect 470600 115874 470652 115880
rect 470600 106344 470652 106350
rect 470600 106286 470652 106292
rect 470612 96626 470640 106286
rect 470600 96620 470652 96626
rect 470600 96562 470652 96568
rect 470600 87032 470652 87038
rect 470600 86974 470652 86980
rect 470612 77246 470640 86974
rect 470600 77240 470652 77246
rect 470600 77182 470652 77188
rect 470600 67652 470652 67658
rect 470600 67594 470652 67600
rect 470612 57934 470640 67594
rect 470600 57928 470652 57934
rect 470600 57870 470652 57876
rect 470600 48340 470652 48346
rect 470600 48282 470652 48288
rect 470612 19310 470640 48282
rect 470600 19304 470652 19310
rect 470600 19246 470652 19252
rect 470600 9716 470652 9722
rect 470600 9658 470652 9664
rect 470612 5642 470640 9658
rect 470600 5636 470652 5642
rect 470600 5578 470652 5584
rect 472716 4208 472768 4214
rect 472716 4150 472768 4156
rect 469232 1414 470364 1442
rect 470336 480 470364 1414
rect 471520 604 471572 610
rect 471520 546 471572 552
rect 471532 480 471560 546
rect 472728 480 472756 4150
rect 475396 3126 475424 336942
rect 476026 29336 476082 29345
rect 476026 29271 476082 29280
rect 476040 29186 476068 29271
rect 476210 29200 476266 29209
rect 476040 29158 476210 29186
rect 476210 29135 476266 29144
rect 475568 16856 475620 16862
rect 475566 16824 475568 16833
rect 475620 16824 475622 16833
rect 475566 16759 475622 16768
rect 476304 5772 476356 5778
rect 476304 5714 476356 5720
rect 475108 3120 475160 3126
rect 475108 3062 475160 3068
rect 475384 3120 475436 3126
rect 475384 3062 475436 3068
rect 473912 2916 473964 2922
rect 473912 2858 473964 2864
rect 473924 480 473952 2858
rect 475120 480 475148 3062
rect 476316 480 476344 5714
rect 477604 3346 477632 337010
rect 482926 76392 482982 76401
rect 482926 76327 482982 76336
rect 482940 76129 482968 76327
rect 482926 76120 482982 76129
rect 482926 76055 482982 76064
rect 482928 16856 482980 16862
rect 482926 16824 482928 16833
rect 482980 16824 482982 16833
rect 482926 16759 482982 16768
rect 483480 5976 483532 5982
rect 483480 5918 483532 5924
rect 479892 5840 479944 5846
rect 479892 5782 479944 5788
rect 477604 3318 478736 3346
rect 477500 3120 477552 3126
rect 477500 3062 477552 3068
rect 477512 480 477540 3062
rect 478708 480 478736 3318
rect 479904 480 479932 5782
rect 482284 3120 482336 3126
rect 482284 3062 482336 3068
rect 481088 2984 481140 2990
rect 481088 2926 481140 2932
rect 481100 480 481128 2926
rect 482296 480 482324 3062
rect 483492 480 483520 5918
rect 484584 5908 484636 5914
rect 484584 5850 484636 5856
rect 484596 480 484624 5850
rect 485792 480 485820 337078
rect 491206 87408 491262 87417
rect 491206 87343 491262 87352
rect 491220 87009 491248 87343
rect 491206 87000 491262 87009
rect 491206 86935 491262 86944
rect 487802 76392 487858 76401
rect 487802 76327 487858 76336
rect 487816 75993 487844 76327
rect 487802 75984 487858 75993
rect 487802 75919 487858 75928
rect 491206 29472 491262 29481
rect 491206 29407 491262 29416
rect 491220 29073 491248 29407
rect 491206 29064 491262 29073
rect 491206 28999 491262 29008
rect 487802 17096 487858 17105
rect 487802 17031 487858 17040
rect 487816 16697 487844 17031
rect 487802 16688 487858 16697
rect 487802 16623 487858 16632
rect 490564 6860 490616 6866
rect 490564 6802 490616 6808
rect 486976 6112 487028 6118
rect 486976 6054 487028 6060
rect 486988 480 487016 6054
rect 488172 6044 488224 6050
rect 488172 5986 488224 5992
rect 488184 480 488212 5986
rect 489368 3052 489420 3058
rect 489368 2994 489420 3000
rect 489380 480 489408 2994
rect 490576 480 490604 6802
rect 491760 6792 491812 6798
rect 491760 6734 491812 6740
rect 491772 480 491800 6734
rect 492692 3482 492720 337146
rect 494612 87168 494664 87174
rect 494612 87110 494664 87116
rect 494624 87009 494652 87110
rect 494610 87000 494666 87009
rect 494610 86935 494666 86944
rect 492772 29096 492824 29102
rect 492770 29064 492772 29073
rect 492824 29064 492826 29073
rect 492770 28999 492826 29008
rect 495348 6724 495400 6730
rect 495348 6666 495400 6672
rect 494152 6588 494204 6594
rect 494152 6530 494204 6536
rect 492692 3454 492996 3482
rect 492968 480 492996 3454
rect 494164 480 494192 6530
rect 495360 480 495388 6666
rect 497740 6656 497792 6662
rect 497740 6598 497792 6604
rect 496544 3256 496596 3262
rect 496544 3198 496596 3204
rect 496556 480 496584 3198
rect 497752 480 497780 6598
rect 498936 6520 498988 6526
rect 498936 6462 498988 6468
rect 498948 480 498976 6462
rect 499592 3482 499620 338030
rect 525064 338020 525116 338026
rect 525064 337962 525116 337968
rect 523684 337884 523736 337890
rect 523684 337826 523736 337832
rect 520924 337816 520976 337822
rect 520924 337758 520976 337764
rect 506480 337748 506532 337754
rect 506480 337690 506532 337696
rect 505744 336796 505796 336802
rect 505744 336738 505796 336744
rect 502246 87272 502302 87281
rect 502246 87207 502302 87216
rect 502260 87174 502288 87207
rect 502248 87168 502300 87174
rect 502248 87110 502300 87116
rect 502246 29336 502302 29345
rect 502246 29271 502302 29280
rect 502260 29102 502288 29271
rect 502248 29096 502300 29102
rect 502248 29038 502300 29044
rect 501236 6452 501288 6458
rect 501236 6394 501288 6400
rect 499592 3454 500172 3482
rect 500144 480 500172 3454
rect 501248 480 501276 6394
rect 502432 6384 502484 6390
rect 502432 6326 502484 6332
rect 502444 480 502472 6326
rect 504824 6316 504876 6322
rect 504824 6258 504876 6264
rect 503628 3324 503680 3330
rect 503628 3266 503680 3272
rect 503640 480 503668 3266
rect 504836 480 504864 6258
rect 505756 3194 505784 336738
rect 506020 6248 506072 6254
rect 506020 6190 506072 6196
rect 505744 3188 505796 3194
rect 505744 3130 505796 3136
rect 506032 480 506060 6190
rect 506492 3482 506520 337690
rect 518164 337612 518216 337618
rect 518164 337554 518216 337560
rect 514024 337544 514076 337550
rect 514024 337486 514076 337492
rect 510620 337408 510672 337414
rect 510620 337350 510672 337356
rect 512642 337376 512698 337385
rect 509884 336864 509936 336870
rect 509884 336806 509936 336812
rect 509608 7336 509660 7342
rect 509608 7278 509660 7284
rect 508412 6180 508464 6186
rect 508412 6122 508464 6128
rect 506492 3454 507256 3482
rect 507228 480 507256 3454
rect 508424 480 508452 6122
rect 509620 480 509648 7278
rect 509896 3058 509924 336806
rect 510632 3482 510660 337350
rect 512642 337311 512698 337320
rect 512000 4276 512052 4282
rect 512000 4218 512052 4224
rect 510632 3454 510844 3482
rect 509884 3052 509936 3058
rect 509884 2994 509936 3000
rect 510816 480 510844 3454
rect 512012 480 512040 4218
rect 512656 3262 512684 337311
rect 513196 7404 513248 7410
rect 513196 7346 513248 7352
rect 512644 3256 512696 3262
rect 512644 3198 512696 3204
rect 513208 480 513236 7346
rect 514036 3398 514064 337486
rect 516784 337476 516836 337482
rect 516784 337418 516836 337424
rect 516796 11778 516824 337418
rect 516704 11750 516824 11778
rect 516704 6934 516732 11750
rect 516784 7472 516836 7478
rect 516784 7414 516836 7420
rect 516692 6928 516744 6934
rect 516692 6870 516744 6876
rect 515588 4344 515640 4350
rect 515588 4286 515640 4292
rect 514024 3392 514076 3398
rect 514024 3334 514076 3340
rect 514392 3324 514444 3330
rect 514392 3266 514444 3272
rect 514404 480 514432 3266
rect 515600 480 515628 4286
rect 516796 480 516824 7414
rect 516876 6928 516928 6934
rect 516876 6870 516928 6876
rect 516888 3330 516916 6870
rect 517888 3392 517940 3398
rect 517888 3334 517940 3340
rect 516876 3324 516928 3330
rect 516876 3266 516928 3272
rect 517900 480 517928 3334
rect 518176 2854 518204 337554
rect 520280 7540 520332 7546
rect 520280 7482 520332 7488
rect 519084 4412 519136 4418
rect 519084 4354 519136 4360
rect 518164 2848 518216 2854
rect 518164 2790 518216 2796
rect 519096 480 519124 4354
rect 520292 480 520320 7482
rect 520936 2990 520964 337758
rect 521016 337680 521068 337686
rect 521016 337622 521068 337628
rect 520924 2984 520976 2990
rect 520924 2926 520976 2932
rect 521028 2922 521056 337622
rect 522672 4480 522724 4486
rect 522672 4422 522724 4428
rect 521476 4140 521528 4146
rect 521476 4082 521528 4088
rect 521016 2916 521068 2922
rect 521016 2858 521068 2864
rect 521488 480 521516 4082
rect 522684 480 522712 4422
rect 523696 3058 523724 337826
rect 523868 8288 523920 8294
rect 523868 8230 523920 8236
rect 523684 3052 523736 3058
rect 523684 2994 523736 3000
rect 523880 480 523908 8230
rect 525076 6882 525104 337962
rect 527824 337952 527876 337958
rect 527824 337894 527876 337900
rect 527456 8220 527508 8226
rect 527456 8162 527508 8168
rect 524984 6854 525104 6882
rect 524984 3126 525012 6854
rect 526260 4548 526312 4554
rect 526260 4490 526312 4496
rect 525064 3392 525116 3398
rect 525064 3334 525116 3340
rect 524972 3120 525024 3126
rect 524972 3062 525024 3068
rect 525076 480 525104 3334
rect 526272 480 526300 4490
rect 527468 480 527496 8162
rect 527836 3398 527864 337894
rect 529204 337340 529256 337346
rect 529204 337282 529256 337288
rect 529216 4146 529244 337282
rect 530584 337272 530636 337278
rect 530584 337214 530636 337220
rect 529848 4616 529900 4622
rect 529848 4558 529900 4564
rect 529204 4140 529256 4146
rect 529204 4082 529256 4088
rect 528652 4072 528704 4078
rect 528652 4014 528704 4020
rect 527824 3392 527876 3398
rect 527824 3334 527876 3340
rect 528664 480 528692 4014
rect 529860 480 529888 4558
rect 530596 4078 530624 337214
rect 579988 322924 580040 322930
rect 579988 322866 580040 322872
rect 580000 322697 580028 322866
rect 579986 322688 580042 322697
rect 579986 322623 580042 322632
rect 580092 310865 580120 578886
rect 580078 310856 580134 310865
rect 580078 310791 580134 310800
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 580184 275777 580212 580094
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 252544 580224 252550
rect 580172 252486 580224 252492
rect 580184 252249 580212 252486
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580276 111489 580304 583374
rect 580356 578604 580408 578610
rect 580356 578546 580408 578552
rect 580368 123185 580396 578546
rect 580460 134881 580488 583442
rect 580540 578672 580592 578678
rect 580540 578614 580592 578620
rect 580552 170105 580580 578614
rect 580644 205329 580672 583510
rect 580908 578876 580960 578882
rect 580908 578818 580960 578824
rect 580724 578808 580776 578814
rect 580724 578750 580776 578756
rect 580736 217025 580764 578750
rect 580816 578740 580868 578746
rect 580816 578682 580868 578688
rect 580828 228857 580856 578682
rect 580920 263945 580948 578818
rect 580906 263936 580962 263945
rect 580906 263871 580962 263880
rect 580814 228848 580870 228857
rect 580814 228783 580870 228792
rect 580722 217016 580778 217025
rect 580722 216951 580778 216960
rect 580630 205320 580686 205329
rect 580630 205255 580686 205264
rect 580538 170096 580594 170105
rect 580538 170031 580594 170040
rect 580446 134872 580502 134881
rect 580446 134807 580502 134816
rect 580354 123176 580410 123185
rect 580354 123111 580410 123120
rect 580262 111480 580318 111489
rect 580262 111415 580318 111424
rect 531044 8152 531096 8158
rect 531044 8094 531096 8100
rect 530584 4072 530636 4078
rect 530584 4014 530636 4020
rect 531056 480 531084 8094
rect 534540 8084 534592 8090
rect 534540 8026 534592 8032
rect 533436 4684 533488 4690
rect 533436 4626 533488 4632
rect 532240 2848 532292 2854
rect 532240 2790 532292 2796
rect 532252 480 532280 2790
rect 533448 480 533476 4626
rect 534552 480 534580 8026
rect 538128 8016 538180 8022
rect 538128 7958 538180 7964
rect 536932 4752 536984 4758
rect 536932 4694 536984 4700
rect 535736 4004 535788 4010
rect 535736 3946 535788 3952
rect 535748 480 535776 3946
rect 536944 480 536972 4694
rect 538140 480 538168 7958
rect 541716 7948 541768 7954
rect 541716 7890 541768 7896
rect 540520 5500 540572 5506
rect 540520 5442 540572 5448
rect 539324 2916 539376 2922
rect 539324 2858 539376 2864
rect 539336 480 539364 2858
rect 540532 480 540560 5442
rect 541728 480 541756 7890
rect 545304 7880 545356 7886
rect 545304 7822 545356 7828
rect 544108 5432 544160 5438
rect 544108 5374 544160 5380
rect 542912 3936 542964 3942
rect 542912 3878 542964 3884
rect 542924 480 542952 3878
rect 544120 480 544148 5374
rect 545316 480 545344 7822
rect 548892 7812 548944 7818
rect 548892 7754 548944 7760
rect 547696 5364 547748 5370
rect 547696 5306 547748 5312
rect 546500 2984 546552 2990
rect 546500 2926 546552 2932
rect 546512 480 546540 2926
rect 547708 480 547736 5306
rect 548904 480 548932 7754
rect 552388 7744 552440 7750
rect 552388 7686 552440 7692
rect 551192 5296 551244 5302
rect 551192 5238 551244 5244
rect 550088 3868 550140 3874
rect 550088 3810 550140 3816
rect 550100 480 550128 3810
rect 551204 480 551232 5238
rect 552400 480 552428 7686
rect 555976 7676 556028 7682
rect 555976 7618 556028 7624
rect 554780 5228 554832 5234
rect 554780 5170 554832 5176
rect 553584 3052 553636 3058
rect 553584 2994 553636 3000
rect 553596 480 553624 2994
rect 554792 480 554820 5170
rect 555988 480 556016 7618
rect 559564 7608 559616 7614
rect 559564 7550 559616 7556
rect 558368 5160 558420 5166
rect 558368 5102 558420 5108
rect 557172 3800 557224 3806
rect 557172 3742 557224 3748
rect 557184 480 557212 3742
rect 558380 480 558408 5102
rect 559576 480 559604 7550
rect 561956 5092 562008 5098
rect 561956 5034 562008 5040
rect 560760 3120 560812 3126
rect 560760 3062 560812 3068
rect 560772 480 560800 3062
rect 561968 480 561996 5034
rect 565544 5024 565596 5030
rect 565544 4966 565596 4972
rect 564348 3732 564400 3738
rect 564348 3674 564400 3680
rect 563152 3188 563204 3194
rect 563152 3130 563204 3136
rect 563164 480 563192 3130
rect 564360 480 564388 3674
rect 565556 480 565584 4966
rect 569040 4956 569092 4962
rect 569040 4898 569092 4904
rect 566740 3664 566792 3670
rect 566740 3606 566792 3612
rect 566752 480 566780 3606
rect 567844 3392 567896 3398
rect 567844 3334 567896 3340
rect 567856 480 567884 3334
rect 569052 480 569080 4898
rect 572628 4888 572680 4894
rect 572628 4830 572680 4836
rect 576214 4856 576270 4865
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 570236 3256 570288 3262
rect 570236 3198 570288 3204
rect 570248 480 570276 3198
rect 571444 480 571472 3538
rect 572640 480 572668 4830
rect 576214 4791 576270 4800
rect 579804 4820 579856 4826
rect 575020 4140 575072 4146
rect 575020 4082 575072 4088
rect 573824 3528 573876 3534
rect 573824 3470 573876 3476
rect 573836 480 573864 3470
rect 575032 480 575060 4082
rect 576228 480 576256 4791
rect 579804 4762 579856 4768
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 577412 3324 577464 3330
rect 577412 3266 577464 3272
rect 577424 480 577452 3266
rect 578620 480 578648 3402
rect 579816 480 579844 4762
rect 582196 4072 582248 4078
rect 582196 4014 582248 4020
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 4014
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 4802 583480 4858 583536
rect 3054 567332 3056 567352
rect 3056 567332 3108 567352
rect 3108 567332 3110 567352
rect 3054 567296 3110 567332
rect 2778 553052 2780 553072
rect 2780 553052 2832 553072
rect 2832 553052 2834 553072
rect 2778 553016 2834 553052
rect 3054 538636 3056 538656
rect 3056 538636 3108 538656
rect 3108 538636 3110 538656
rect 3054 538600 3110 538636
rect 3054 509904 3110 509960
rect 2778 495488 2834 495544
rect 2962 481108 2964 481128
rect 2964 481108 3016 481128
rect 3016 481108 3018 481128
rect 2962 481072 3018 481108
rect 3146 452376 3202 452432
rect 3146 437960 3202 438016
rect 3146 423680 3202 423736
rect 3238 394984 3294 395040
rect 3238 380568 3294 380624
rect 3330 366152 3386 366208
rect 3330 323040 3386 323096
rect 2778 308796 2780 308816
rect 2780 308796 2832 308816
rect 2832 308796 2834 308816
rect 2778 308760 2834 308796
rect 2962 295160 3018 295216
rect 2962 294344 3018 294400
rect 2778 251232 2834 251288
rect 3054 236952 3110 237008
rect 2778 165008 2834 165064
rect 3330 150728 3386 150784
rect 2778 136312 2834 136368
rect 2778 122032 2834 122088
rect 4066 280064 4122 280120
rect 3974 265648 4030 265704
rect 3882 222536 3938 222592
rect 3790 208120 3846 208176
rect 3698 193840 3754 193896
rect 3606 179424 3662 179480
rect 3514 107616 3570 107672
rect 3422 93200 3478 93256
rect 2778 78920 2834 78976
rect 3330 64504 3386 64560
rect 5078 582528 5134 582584
rect 2778 50088 2834 50144
rect 10322 337320 10378 337376
rect 3146 35844 3148 35864
rect 3148 35844 3200 35864
rect 3200 35844 3202 35864
rect 3146 35808 3202 35844
rect 3146 11600 3202 11656
rect 3146 7112 3202 7168
rect 6458 3304 6514 3360
rect 17222 582800 17278 582856
rect 24122 582664 24178 582720
rect 293958 583208 294014 583264
rect 300306 583344 300362 583400
rect 378138 700304 378194 700360
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 460294 583480 460350 583536
rect 420274 583072 420330 583128
rect 426622 582936 426678 582992
rect 449806 582800 449862 582856
rect 447690 582528 447746 582584
rect 462410 582664 462466 582720
rect 468482 579672 468538 579728
rect 231122 579264 231178 579320
rect 232962 579264 233018 579320
rect 235262 579264 235318 579320
rect 237194 579264 237250 579320
rect 239402 579264 239458 579320
rect 241426 579264 241482 579320
rect 249522 579264 249578 579320
rect 466458 579264 466514 579320
rect 51630 6160 51686 6216
rect 57978 337748 58034 337784
rect 57978 337728 57980 337748
rect 57980 337728 58032 337748
rect 58032 337728 58034 337748
rect 67546 337748 67602 337784
rect 67546 337728 67548 337748
rect 67548 337728 67600 337748
rect 67600 337728 67602 337748
rect 132590 8880 132646 8936
rect 129002 7520 129058 7576
rect 208674 4800 208730 4856
rect 231950 337320 232006 337376
rect 232134 153176 232190 153232
rect 232318 153176 232374 153232
rect 232318 48320 232374 48376
rect 232318 47912 232374 47968
rect 232042 3304 232098 3360
rect 236274 309304 236330 309360
rect 236274 309168 236330 309224
rect 236274 270408 236330 270464
rect 236458 260888 236514 260944
rect 236274 251096 236330 251152
rect 236550 251096 236606 251152
rect 236642 232056 236698 232112
rect 236274 231920 236330 231976
rect 236458 222128 236514 222184
rect 236274 212608 236330 212664
rect 236274 212472 236330 212528
rect 236550 212472 236606 212528
rect 236550 202952 236606 203008
rect 236274 193296 236330 193352
rect 236274 193160 236330 193216
rect 236550 193160 236606 193216
rect 236274 154536 236330 154592
rect 236458 154536 236514 154592
rect 236274 135224 236330 135280
rect 236458 135224 236514 135280
rect 236274 115912 236330 115968
rect 236458 115912 236514 115968
rect 236274 96600 236330 96656
rect 236642 96600 236698 96656
rect 239034 135224 239090 135280
rect 239218 135224 239274 135280
rect 239126 96600 239182 96656
rect 239310 96600 239366 96656
rect 240138 29164 240194 29200
rect 240138 29144 240140 29164
rect 240140 29144 240192 29164
rect 240192 29144 240194 29164
rect 244462 259392 244518 259448
rect 244646 259392 244702 259448
rect 244278 241440 244334 241496
rect 244462 241440 244518 241496
rect 244278 222128 244334 222184
rect 244462 222128 244518 222184
rect 244278 202816 244334 202872
rect 244462 202816 244518 202872
rect 244278 154536 244334 154592
rect 244462 154536 244518 154592
rect 244278 135224 244334 135280
rect 244462 135224 244518 135280
rect 247130 144900 247186 144936
rect 247130 144880 247132 144900
rect 247132 144880 247184 144900
rect 247184 144880 247186 144900
rect 247314 144880 247370 144936
rect 249154 334192 249210 334248
rect 249154 328480 249210 328536
rect 249154 322224 249210 322280
rect 249154 317600 249210 317656
rect 249246 298016 249302 298072
rect 249246 288496 249302 288552
rect 249246 288360 249302 288416
rect 249246 278976 249302 279032
rect 249430 277344 249486 277400
rect 249430 267824 249486 267880
rect 249246 212472 249302 212528
rect 249246 205400 249302 205456
rect 249614 202816 249670 202872
rect 249614 196560 249670 196616
rect 249246 191528 249302 191584
rect 249246 182144 249302 182200
rect 249430 180512 249486 180568
rect 249430 173848 249486 173904
rect 249706 29008 249762 29064
rect 250074 288360 250130 288416
rect 250350 288360 250406 288416
rect 250350 154672 250406 154728
rect 250074 154536 250130 154592
rect 250258 135360 250314 135416
rect 250074 135224 250130 135280
rect 249982 6160 250038 6216
rect 251178 87100 251234 87136
rect 251178 87080 251180 87100
rect 251180 87080 251232 87100
rect 251232 87080 251234 87100
rect 251178 27648 251234 27704
rect 251454 241440 251510 241496
rect 251638 241440 251694 241496
rect 251454 222128 251510 222184
rect 251638 222128 251694 222184
rect 251454 202816 251510 202872
rect 251638 202816 251694 202872
rect 251454 183504 251510 183560
rect 251638 183504 251694 183560
rect 251454 154536 251510 154592
rect 251638 154536 251694 154592
rect 251454 48456 251510 48512
rect 251362 48320 251418 48376
rect 251362 27648 251418 27704
rect 259366 17040 259422 17096
rect 259366 16632 259422 16688
rect 259550 280200 259606 280256
rect 259918 280200 259974 280256
rect 259642 202816 259698 202872
rect 259918 202816 259974 202872
rect 259642 164212 259698 164248
rect 259642 164192 259644 164212
rect 259644 164192 259696 164212
rect 259696 164192 259698 164212
rect 259918 164192 259974 164248
rect 260654 87100 260710 87136
rect 260654 87080 260656 87100
rect 260656 87080 260708 87100
rect 260708 87080 260710 87100
rect 260746 63688 260802 63744
rect 260746 63552 260802 63608
rect 262494 247016 262550 247072
rect 262770 246880 262826 246936
rect 262586 125588 262642 125624
rect 262586 125568 262588 125588
rect 262588 125568 262640 125588
rect 262640 125568 262642 125588
rect 262770 125588 262826 125624
rect 262770 125568 262772 125588
rect 262772 125568 262824 125588
rect 262824 125568 262826 125588
rect 263414 63688 263470 63744
rect 263598 63688 263654 63744
rect 264978 182144 265034 182200
rect 265346 219408 265402 219464
rect 265530 219408 265586 219464
rect 265162 211112 265218 211168
rect 265346 211112 265402 211168
rect 265254 182144 265310 182200
rect 267738 278704 267794 278760
rect 267830 278568 267886 278624
rect 267738 248376 267794 248432
rect 268014 248376 268070 248432
rect 266634 211112 266690 211168
rect 266818 211112 266874 211168
rect 267738 209752 267794 209808
rect 267922 209752 267978 209808
rect 267738 182144 267794 182200
rect 267922 182144 267978 182200
rect 266634 173884 266636 173904
rect 266636 173884 266688 173904
rect 266688 173884 266690 173904
rect 266634 173848 266690 173884
rect 266818 173884 266820 173904
rect 266820 173884 266872 173904
rect 266872 173884 266874 173904
rect 266818 173848 266874 173884
rect 266726 135360 266782 135416
rect 266634 135244 266690 135280
rect 266634 135224 266636 135244
rect 266636 135224 266688 135244
rect 266688 135224 266690 135244
rect 267738 125588 267794 125624
rect 267738 125568 267740 125588
rect 267740 125568 267792 125588
rect 267792 125568 267794 125588
rect 267922 125588 267978 125624
rect 267922 125568 267924 125588
rect 267924 125568 267976 125588
rect 267976 125568 267978 125588
rect 266726 116048 266782 116104
rect 266634 115912 266690 115968
rect 270498 325624 270554 325680
rect 270498 125568 270554 125624
rect 270774 325624 270830 325680
rect 270682 314608 270738 314664
rect 270866 314608 270922 314664
rect 270682 220768 270738 220824
rect 270958 220768 271014 220824
rect 270774 209752 270830 209808
rect 270958 209752 271014 209808
rect 270774 180784 270830 180840
rect 271050 180784 271106 180840
rect 270682 125588 270738 125624
rect 270682 125568 270684 125588
rect 270684 125568 270736 125588
rect 270736 125568 270738 125588
rect 270682 106276 270738 106312
rect 270682 106256 270684 106276
rect 270684 106256 270736 106276
rect 270736 106256 270738 106276
rect 270866 106256 270922 106312
rect 271878 229064 271934 229120
rect 272062 269048 272118 269104
rect 272246 269048 272302 269104
rect 272154 259428 272156 259448
rect 272156 259428 272208 259448
rect 272208 259428 272210 259448
rect 272154 259392 272210 259428
rect 272430 259392 272486 259448
rect 272062 229084 272118 229120
rect 272062 229064 272064 229084
rect 272064 229064 272116 229084
rect 272116 229064 272118 229084
rect 272154 202816 272210 202872
rect 272338 202680 272394 202736
rect 272154 183504 272210 183560
rect 272338 183368 272394 183424
rect 273074 63688 273130 63744
rect 273258 63688 273314 63744
rect 273074 40160 273130 40216
rect 273258 40160 273314 40216
rect 278778 29300 278834 29336
rect 278778 29280 278780 29300
rect 278780 29280 278832 29300
rect 278832 29280 278834 29300
rect 278778 16532 278780 16552
rect 278780 16532 278832 16552
rect 278832 16532 278834 16552
rect 278778 16496 278834 16532
rect 281262 29144 281318 29200
rect 282734 40160 282790 40216
rect 282918 40160 282974 40216
rect 283102 7520 283158 7576
rect 284574 278704 284630 278760
rect 284758 278704 284814 278760
rect 284666 220768 284722 220824
rect 284850 220768 284906 220824
rect 284666 201456 284722 201512
rect 284850 201456 284906 201512
rect 284666 193160 284722 193216
rect 284850 193160 284906 193216
rect 285494 157936 285550 157992
rect 285494 157392 285550 157448
rect 284482 8880 284538 8936
rect 285770 202816 285826 202872
rect 286046 261024 286102 261080
rect 285954 260888 286010 260944
rect 286046 249772 286048 249792
rect 286048 249772 286100 249792
rect 286100 249772 286102 249792
rect 286046 249736 286102 249772
rect 285954 249600 286010 249656
rect 285954 222128 286010 222184
rect 286138 222128 286194 222184
rect 285954 220768 286010 220824
rect 286138 220768 286194 220824
rect 285954 202852 285956 202872
rect 285956 202852 286008 202872
rect 286008 202852 286010 202872
rect 285954 202816 286010 202852
rect 285954 172624 286010 172680
rect 286046 172488 286102 172544
rect 285954 122712 286010 122768
rect 286230 122712 286286 122768
rect 285954 38800 286010 38856
rect 285954 38528 286010 38584
rect 288806 258168 288862 258224
rect 288806 258032 288862 258088
rect 288806 201456 288862 201512
rect 288990 201456 289046 201512
rect 288714 64776 288770 64832
rect 288898 64776 288954 64832
rect 290370 219544 290426 219600
rect 290094 219408 290150 219464
rect 290554 16632 290610 16688
rect 291474 306312 291530 306368
rect 291750 306312 291806 306368
rect 291658 219408 291714 219464
rect 292026 219408 292082 219464
rect 291474 164192 291530 164248
rect 291658 164192 291714 164248
rect 295246 87488 295302 87544
rect 295246 86944 295302 87000
rect 295246 75928 295302 75984
rect 295246 75520 295302 75576
rect 295614 275984 295670 276040
rect 295798 275984 295854 276040
rect 295522 247016 295578 247072
rect 295890 247016 295946 247072
rect 296626 87080 296682 87136
rect 296626 86944 296682 87000
rect 296626 29552 296682 29608
rect 296626 29280 296682 29336
rect 298098 29280 298154 29336
rect 298098 28872 298154 28928
rect 298006 16768 298062 16824
rect 298098 16632 298154 16688
rect 301318 317464 301374 317520
rect 301226 317328 301282 317384
rect 301042 241440 301098 241496
rect 301134 241304 301190 241360
rect 301042 222128 301098 222184
rect 301134 221992 301190 222048
rect 301042 202816 301098 202872
rect 301134 202680 301190 202736
rect 301042 144880 301098 144936
rect 301226 144880 301282 144936
rect 301226 66272 301282 66328
rect 301226 66000 301282 66056
rect 306286 76064 306342 76120
rect 306286 75792 306342 75848
rect 306378 40180 306434 40216
rect 306378 40160 306380 40180
rect 306380 40160 306432 40180
rect 306432 40160 306434 40180
rect 306378 28892 306434 28928
rect 306378 28872 306380 28892
rect 306380 28872 306432 28892
rect 306432 28872 306434 28892
rect 307758 337592 307814 337648
rect 306838 124208 306894 124264
rect 307022 124208 307078 124264
rect 306838 103536 306894 103592
rect 307022 103536 307078 103592
rect 307390 3304 307446 3360
rect 310794 193160 310850 193216
rect 311070 193160 311126 193216
rect 310886 153312 310942 153368
rect 310794 153196 310850 153232
rect 310794 153176 310796 153196
rect 310796 153176 310848 153196
rect 310848 153176 310850 153196
rect 310978 116048 311034 116104
rect 310794 115912 310850 115968
rect 310886 45600 310942 45656
rect 311070 45600 311126 45656
rect 312082 4936 312138 4992
rect 315946 87352 316002 87408
rect 315946 87080 316002 87136
rect 315946 40024 316002 40080
rect 315946 28892 316002 28928
rect 315946 28872 315948 28892
rect 315948 28872 316000 28892
rect 316000 28872 316002 28892
rect 315946 4972 315948 4992
rect 315948 4972 316000 4992
rect 316000 4972 316002 4992
rect 315946 4936 316002 4972
rect 314658 4800 314714 4856
rect 317326 337592 317382 337648
rect 317326 29280 317382 29336
rect 317326 28872 317382 28928
rect 317786 115912 317842 115968
rect 317970 115912 318026 115968
rect 320822 16668 320824 16688
rect 320824 16668 320876 16688
rect 320876 16668 320878 16688
rect 320822 16632 320878 16668
rect 322202 29280 322258 29336
rect 322202 29008 322258 29064
rect 323214 288360 323270 288416
rect 323490 288360 323546 288416
rect 323306 269048 323362 269104
rect 323398 268912 323454 268968
rect 323306 211112 323362 211168
rect 323490 211112 323546 211168
rect 323306 193196 323308 193216
rect 323308 193196 323360 193216
rect 323360 193196 323362 193216
rect 323306 193160 323362 193196
rect 323490 193196 323492 193216
rect 323492 193196 323544 193216
rect 323544 193196 323546 193216
rect 323490 193160 323546 193196
rect 324226 157392 324282 157448
rect 324226 157120 324282 157176
rect 323398 116048 323454 116104
rect 323306 115912 323362 115968
rect 325606 298152 325662 298208
rect 324686 269048 324742 269104
rect 324870 269048 324926 269104
rect 324594 183504 324650 183560
rect 324778 183504 324834 183560
rect 324594 144880 324650 144936
rect 324594 144744 324650 144800
rect 325606 16768 325662 16824
rect 325882 298118 325938 298174
rect 325882 296656 325938 296712
rect 326066 296656 326122 296712
rect 325882 240080 325938 240136
rect 326158 240080 326214 240136
rect 325882 144900 325938 144936
rect 325882 144880 325884 144900
rect 325884 144880 325936 144900
rect 325936 144880 325938 144900
rect 326066 144900 326122 144936
rect 326066 144880 326068 144900
rect 326068 144880 326120 144900
rect 326120 144880 326122 144900
rect 327170 230424 327226 230480
rect 327538 230424 327594 230480
rect 327262 212472 327318 212528
rect 327354 212336 327410 212392
rect 327262 145016 327318 145072
rect 327170 144900 327226 144936
rect 327170 144880 327172 144900
rect 327172 144880 327224 144900
rect 327224 144880 327226 144900
rect 328458 87216 328514 87272
rect 328366 87080 328422 87136
rect 328918 75928 328974 75984
rect 329930 103536 329986 103592
rect 330206 315968 330262 316024
rect 330390 315968 330446 316024
rect 330206 249736 330262 249792
rect 330390 249736 330446 249792
rect 330114 103536 330170 103592
rect 330114 28872 330170 28928
rect 330206 28736 330262 28792
rect 331862 29552 331918 29608
rect 331862 29280 331918 29336
rect 333886 157664 333942 157720
rect 333886 157392 333942 157448
rect 336738 240080 336794 240136
rect 336738 183504 336794 183560
rect 336738 115912 336794 115968
rect 336646 17040 336702 17096
rect 336646 16632 336702 16688
rect 337106 273944 337162 274000
rect 336922 260616 336978 260672
rect 336922 240080 336978 240136
rect 337106 220768 337162 220824
rect 337198 220632 337254 220688
rect 336922 183504 336978 183560
rect 337198 162832 337254 162888
rect 337382 162832 337438 162888
rect 336922 115912 336978 115968
rect 338026 76200 338082 76256
rect 337198 56752 337254 56808
rect 337290 56616 337346 56672
rect 339498 144880 339554 144936
rect 339682 144880 339738 144936
rect 341246 299376 341302 299432
rect 341246 289856 341302 289912
rect 341246 280064 341302 280120
rect 341246 270544 341302 270600
rect 341246 260752 341302 260808
rect 341246 251232 341302 251288
rect 341154 240080 341210 240136
rect 341430 240080 341486 240136
rect 341154 202852 341156 202872
rect 341156 202852 341208 202872
rect 341208 202852 341210 202872
rect 341154 202816 341210 202852
rect 341430 202816 341486 202872
rect 342718 337492 342720 337512
rect 342720 337492 342772 337512
rect 342772 337492 342774 337512
rect 342718 337456 342774 337492
rect 345754 337456 345810 337512
rect 347778 86980 347780 87000
rect 347780 86980 347832 87000
rect 347832 86980 347834 87000
rect 347778 86944 347834 86980
rect 347778 29044 347780 29064
rect 347780 29044 347832 29064
rect 347832 29044 347834 29064
rect 347778 29008 347834 29044
rect 347778 16924 347834 16960
rect 347778 16904 347780 16924
rect 347780 16904 347832 16924
rect 347832 16904 347834 16924
rect 352654 16632 352710 16688
rect 356242 3304 356298 3360
rect 357438 125704 357494 125760
rect 357530 125568 357586 125624
rect 357346 87216 357402 87272
rect 357346 29280 357402 29336
rect 357622 27648 357678 27704
rect 357806 27648 357862 27704
rect 358542 278704 358598 278760
rect 358726 278704 358782 278760
rect 358726 220804 358728 220824
rect 358728 220804 358780 220824
rect 358780 220804 358782 220824
rect 358726 220768 358782 220804
rect 358726 211112 358782 211168
rect 358450 191800 358506 191856
rect 358634 191800 358690 191856
rect 358542 172488 358598 172544
rect 358726 172488 358782 172544
rect 358542 153176 358598 153232
rect 358726 153176 358782 153232
rect 358726 86944 358782 87000
rect 359186 327256 359242 327312
rect 359186 327120 359242 327176
rect 359002 86944 359058 87000
rect 360474 193160 360530 193216
rect 360658 193160 360714 193216
rect 360198 162832 360254 162888
rect 360566 162832 360622 162888
rect 360198 153176 360254 153232
rect 360382 153176 360438 153232
rect 360474 106392 360530 106448
rect 360382 106276 360438 106312
rect 360382 106256 360384 106276
rect 360384 106256 360436 106276
rect 360436 106256 360438 106276
rect 360290 96620 360346 96656
rect 360290 96600 360292 96620
rect 360292 96600 360344 96620
rect 360344 96600 360346 96620
rect 360566 96600 360622 96656
rect 364338 157564 364340 157584
rect 364340 157564 364392 157584
rect 364392 157564 364394 157584
rect 364338 157528 364394 157564
rect 367006 222128 367062 222184
rect 367006 212608 367062 212664
rect 367098 87080 367154 87136
rect 367098 86944 367154 87000
rect 367006 77424 367062 77480
rect 367006 77288 367062 77344
rect 367098 63724 367100 63744
rect 367100 63724 367152 63744
rect 367152 63724 367154 63744
rect 367098 63688 367154 63724
rect 367098 40196 367100 40216
rect 367100 40196 367152 40216
rect 367152 40196 367154 40216
rect 367098 40160 367154 40196
rect 367098 29008 367154 29064
rect 367006 16904 367062 16960
rect 367006 16768 367062 16824
rect 369674 16804 369676 16824
rect 369676 16804 369728 16824
rect 369728 16804 369730 16824
rect 369674 16768 369730 16804
rect 369858 76100 369860 76120
rect 369860 76100 369912 76120
rect 369912 76100 369914 76120
rect 369858 76064 369914 76100
rect 372526 241440 372582 241496
rect 372710 241440 372766 241496
rect 372526 222128 372582 222184
rect 372710 222128 372766 222184
rect 372526 202816 372582 202872
rect 372710 202816 372766 202872
rect 372802 173848 372858 173904
rect 372986 173848 373042 173904
rect 372802 164212 372858 164248
rect 372802 164192 372804 164212
rect 372804 164192 372856 164212
rect 372856 164192 372858 164212
rect 372986 164192 373042 164248
rect 373814 157564 373816 157584
rect 373816 157564 373868 157584
rect 373868 157564 373870 157584
rect 373814 157528 373870 157564
rect 375378 86944 375434 87000
rect 375562 309168 375618 309224
rect 375746 309168 375802 309224
rect 375562 106256 375618 106312
rect 375746 106256 375802 106312
rect 375654 86944 375710 87000
rect 376942 241440 376998 241496
rect 377126 241440 377182 241496
rect 376942 222128 376998 222184
rect 377126 222128 377182 222184
rect 376942 202816 376998 202872
rect 377126 202816 377182 202872
rect 376942 183504 376998 183560
rect 377126 183504 377182 183560
rect 376942 106392 376998 106448
rect 377126 106392 377182 106448
rect 376666 76200 376722 76256
rect 376666 63824 376722 63880
rect 376666 40296 376722 40352
rect 376666 29280 376722 29336
rect 376666 16904 376722 16960
rect 376758 9560 376814 9616
rect 377034 9560 377090 9616
rect 378506 63860 378508 63880
rect 378508 63860 378560 63880
rect 378560 63860 378562 63880
rect 378506 63824 378562 63860
rect 386786 325896 386842 325952
rect 386786 325760 386842 325816
rect 386786 325624 386842 325680
rect 386970 325624 387026 325680
rect 386418 231784 386474 231840
rect 386786 231784 386842 231840
rect 386418 212472 386474 212528
rect 386602 212472 386658 212528
rect 386602 202816 386658 202872
rect 386878 202816 386934 202872
rect 386602 183504 386658 183560
rect 386970 183504 387026 183560
rect 386418 157936 386474 157992
rect 386418 157664 386474 157720
rect 386510 154536 386566 154592
rect 386786 154536 386842 154592
rect 386418 135224 386474 135280
rect 386694 135224 386750 135280
rect 386418 115912 386474 115968
rect 386602 115912 386658 115968
rect 386418 76472 386474 76528
rect 386418 76200 386474 76256
rect 386326 63860 386328 63880
rect 386328 63860 386380 63880
rect 386380 63860 386382 63880
rect 386326 63824 386382 63860
rect 386510 37304 386566 37360
rect 386694 37304 386750 37360
rect 386326 17176 386382 17232
rect 386326 16768 386382 16824
rect 396078 157548 396134 157584
rect 396078 157528 396080 157548
rect 396080 157528 396132 157548
rect 396132 157528 396134 157548
rect 396078 76084 396134 76120
rect 396078 76064 396080 76084
rect 396080 76064 396132 76084
rect 396132 76064 396134 76084
rect 399390 76084 399446 76120
rect 399390 76064 399392 76084
rect 399392 76064 399444 76084
rect 399444 76064 399446 76084
rect 398746 16632 398802 16688
rect 398930 16632 398986 16688
rect 400770 157548 400826 157584
rect 400770 157528 400772 157548
rect 400772 157528 400824 157548
rect 400824 157528 400826 157548
rect 414018 76084 414074 76120
rect 414018 76064 414020 76084
rect 414020 76064 414072 76084
rect 414072 76064 414074 76084
rect 417882 157548 417938 157584
rect 417882 157528 417884 157548
rect 417884 157528 417936 157548
rect 417936 157528 417938 157548
rect 417882 63708 417938 63744
rect 417882 63688 417884 63708
rect 417884 63688 417936 63708
rect 417936 63688 417938 63708
rect 417882 40196 417884 40216
rect 417884 40196 417936 40216
rect 417936 40196 417938 40216
rect 417882 40160 417938 40196
rect 418158 157548 418214 157584
rect 418158 157528 418160 157548
rect 418160 157528 418212 157548
rect 418212 157528 418214 157548
rect 418158 63708 418214 63744
rect 418158 63688 418160 63708
rect 418160 63688 418212 63708
rect 418212 63688 418214 63708
rect 420366 40196 420368 40216
rect 420368 40196 420420 40216
rect 420420 40196 420422 40216
rect 420366 40160 420422 40196
rect 420734 3712 420790 3768
rect 421194 278704 421250 278760
rect 421378 278704 421434 278760
rect 421194 259392 421250 259448
rect 421378 259392 421434 259448
rect 421194 241712 421250 241768
rect 421194 241576 421250 241632
rect 421194 240080 421250 240136
rect 421378 240080 421434 240136
rect 421194 220768 421250 220824
rect 421378 220768 421434 220824
rect 421194 211112 421250 211168
rect 421378 211112 421434 211168
rect 421194 191800 421250 191856
rect 421378 191800 421434 191856
rect 421194 172488 421250 172544
rect 421378 172488 421434 172544
rect 423494 75928 423550 75984
rect 437202 157548 437258 157584
rect 437202 157528 437204 157548
rect 437204 157528 437256 157548
rect 437256 157528 437258 157548
rect 437202 87116 437204 87136
rect 437204 87116 437256 87136
rect 437256 87116 437258 87136
rect 437202 87080 437258 87116
rect 437202 76084 437258 76120
rect 437202 76064 437204 76084
rect 437204 76064 437256 76084
rect 437256 76064 437258 76084
rect 437202 63708 437258 63744
rect 437202 63688 437204 63708
rect 437204 63688 437256 63708
rect 437256 63688 437258 63708
rect 437202 40196 437204 40216
rect 437204 40196 437256 40216
rect 437256 40196 437258 40216
rect 437202 40160 437258 40196
rect 437202 29164 437258 29200
rect 437202 29144 437204 29164
rect 437204 29144 437256 29164
rect 437256 29144 437258 29164
rect 437202 16788 437258 16824
rect 437202 16768 437204 16788
rect 437204 16768 437256 16788
rect 437256 16768 437258 16788
rect 434534 3712 434590 3768
rect 437478 157548 437534 157584
rect 437478 157528 437480 157548
rect 437480 157528 437532 157548
rect 437532 157528 437534 157548
rect 437478 87116 437480 87136
rect 437480 87116 437532 87136
rect 437532 87116 437534 87136
rect 437478 87080 437534 87116
rect 437478 76084 437534 76120
rect 437478 76064 437480 76084
rect 437480 76064 437532 76084
rect 437532 76064 437534 76084
rect 437478 63708 437534 63744
rect 437478 63688 437480 63708
rect 437480 63688 437532 63708
rect 437532 63688 437534 63708
rect 437478 40196 437480 40216
rect 437480 40196 437532 40216
rect 437532 40196 437534 40216
rect 437478 40160 437534 40196
rect 437478 29164 437534 29200
rect 437478 29144 437480 29164
rect 437480 29144 437532 29164
rect 437532 29144 437534 29164
rect 437478 16788 437534 16824
rect 437478 16768 437480 16788
rect 437480 16768 437532 16788
rect 437532 16768 437534 16788
rect 454038 87252 454040 87272
rect 454040 87252 454092 87272
rect 454092 87252 454094 87272
rect 454038 87216 454094 87252
rect 455694 337764 455696 337784
rect 455696 337764 455748 337784
rect 455748 337764 455750 337784
rect 455694 337728 455750 337764
rect 456522 157548 456578 157584
rect 456522 157528 456524 157548
rect 456524 157528 456576 157548
rect 456576 157528 456578 157548
rect 456522 63708 456578 63744
rect 456522 63688 456524 63708
rect 456524 63688 456576 63708
rect 456576 63688 456578 63708
rect 456522 40196 456524 40216
rect 456524 40196 456576 40216
rect 456576 40196 456578 40216
rect 456522 40160 456578 40196
rect 456522 29164 456578 29200
rect 456522 29144 456524 29164
rect 456524 29144 456576 29164
rect 456576 29144 456578 29164
rect 456522 16924 456578 16960
rect 456522 16904 456524 16924
rect 456524 16904 456576 16924
rect 456576 16904 456578 16924
rect 456982 87252 456984 87272
rect 456984 87252 457036 87272
rect 457036 87252 457038 87272
rect 456982 87216 457038 87252
rect 456890 63708 456946 63744
rect 456890 63688 456892 63708
rect 456892 63688 456944 63708
rect 456944 63688 456946 63708
rect 456890 40196 456892 40216
rect 456892 40196 456944 40216
rect 456944 40196 456946 40216
rect 456890 40160 456946 40196
rect 456798 29164 456854 29200
rect 456798 29144 456800 29164
rect 456800 29144 456852 29164
rect 456852 29144 456854 29164
rect 457442 16768 457498 16824
rect 458270 157548 458326 157584
rect 458270 157528 458272 157548
rect 458272 157528 458324 157548
rect 458324 157528 458326 157548
rect 460018 318824 460074 318880
rect 460202 318824 460258 318880
rect 459834 240080 459890 240136
rect 460018 240080 460074 240136
rect 459834 220768 459890 220824
rect 460018 220768 460074 220824
rect 463606 337728 463662 337784
rect 463790 231784 463846 231840
rect 463974 231784 464030 231840
rect 463790 212472 463846 212528
rect 463974 212472 464030 212528
rect 463790 193160 463846 193216
rect 463974 193160 464030 193216
rect 463882 106256 463938 106312
rect 464066 106256 464122 106312
rect 466090 87488 466146 87544
rect 466090 87080 466146 87136
rect 466090 76472 466146 76528
rect 466090 76064 466146 76120
rect 467562 337320 467618 337376
rect 467746 4800 467802 4856
rect 468758 3304 468814 3360
rect 580170 580760 580226 580816
rect 579710 557232 579766 557288
rect 579710 545536 579766 545592
rect 579710 510312 579766 510368
rect 579710 498616 579766 498672
rect 579710 463392 579766 463448
rect 579802 451696 579858 451752
rect 579802 439864 579858 439920
rect 579802 416472 579858 416528
rect 579802 404776 579858 404832
rect 579802 392944 579858 393000
rect 579894 369552 579950 369608
rect 579986 357856 580042 357912
rect 579986 346024 580042 346080
rect 483018 338036 483020 338056
rect 483020 338036 483072 338056
rect 483072 338036 483074 338056
rect 483018 338000 483074 338036
rect 483386 338036 483388 338056
rect 483388 338036 483440 338056
rect 483440 338036 483442 338056
rect 483386 338000 483442 338036
rect 483018 337884 483074 337920
rect 483018 337864 483020 337884
rect 483020 337864 483072 337884
rect 483072 337864 483074 337884
rect 483386 337884 483442 337920
rect 483386 337864 483388 337884
rect 483388 337864 483440 337884
rect 483440 337864 483442 337884
rect 483018 337748 483074 337784
rect 483018 337728 483020 337748
rect 483020 337728 483072 337748
rect 483072 337728 483074 337748
rect 483386 337748 483442 337784
rect 483386 337728 483388 337748
rect 483388 337728 483440 337748
rect 483440 337728 483442 337748
rect 483018 337612 483074 337648
rect 483018 337592 483020 337612
rect 483020 337592 483072 337612
rect 483072 337592 483074 337612
rect 483478 337612 483534 337648
rect 483478 337592 483480 337612
rect 483480 337592 483532 337612
rect 483532 337592 483534 337612
rect 470414 231784 470470 231840
rect 470598 231784 470654 231840
rect 470414 212472 470470 212528
rect 470598 212472 470654 212528
rect 470414 193160 470470 193216
rect 470598 193160 470654 193216
rect 470414 173848 470470 173904
rect 470598 173848 470654 173904
rect 470414 164192 470470 164248
rect 470598 164192 470654 164248
rect 470414 144880 470470 144936
rect 470598 144880 470654 144936
rect 470414 125568 470470 125624
rect 470598 125568 470654 125624
rect 476026 29280 476082 29336
rect 476210 29144 476266 29200
rect 475566 16804 475568 16824
rect 475568 16804 475620 16824
rect 475620 16804 475622 16824
rect 475566 16768 475622 16804
rect 482926 76336 482982 76392
rect 482926 76064 482982 76120
rect 482926 16804 482928 16824
rect 482928 16804 482980 16824
rect 482980 16804 482982 16824
rect 482926 16768 482982 16804
rect 491206 87352 491262 87408
rect 491206 86944 491262 87000
rect 487802 76336 487858 76392
rect 487802 75928 487858 75984
rect 491206 29416 491262 29472
rect 491206 29008 491262 29064
rect 487802 17040 487858 17096
rect 487802 16632 487858 16688
rect 494610 86944 494666 87000
rect 492770 29044 492772 29064
rect 492772 29044 492824 29064
rect 492824 29044 492826 29064
rect 492770 29008 492826 29044
rect 502246 87216 502302 87272
rect 502246 29280 502302 29336
rect 512642 337320 512698 337376
rect 579986 322632 580042 322688
rect 580078 310800 580134 310856
rect 579802 299104 579858 299160
rect 580170 275712 580226 275768
rect 580170 252184 580226 252240
rect 580170 181872 580226 181928
rect 580906 263880 580962 263936
rect 580814 228792 580870 228848
rect 580722 216960 580778 217016
rect 580630 205264 580686 205320
rect 580538 170040 580594 170096
rect 580446 134816 580502 134872
rect 580354 123120 580410 123176
rect 580262 111424 580318 111480
rect 576214 4800 576270 4856
rect 580998 3304 581054 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 378133 700362 378199 700365
rect 8109 700360 378199 700362
rect 8109 700304 8114 700360
rect 8170 700304 378138 700360
rect 378194 700304 378199 700360
rect 8109 700302 378199 700304
rect 8109 700299 8175 700302
rect 378133 700299 378199 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect 4797 583538 4863 583541
rect 460289 583538 460355 583541
rect 4797 583536 460355 583538
rect 4797 583480 4802 583536
rect 4858 583480 460294 583536
rect 460350 583480 460355 583536
rect 4797 583478 460355 583480
rect 4797 583475 4863 583478
rect 460289 583475 460355 583478
rect 300301 583402 300367 583405
rect 465942 583402 465948 583404
rect 300301 583400 465948 583402
rect 300301 583344 300306 583400
rect 300362 583344 465948 583400
rect 300301 583342 465948 583344
rect 300301 583339 300367 583342
rect 465942 583340 465948 583342
rect 466012 583340 466018 583404
rect 293953 583266 294019 583269
rect 465758 583266 465764 583268
rect 293953 583264 465764 583266
rect 293953 583208 293958 583264
rect 294014 583208 465764 583264
rect 293953 583206 465764 583208
rect 293953 583203 294019 583206
rect 465758 583204 465764 583206
rect 465828 583204 465834 583268
rect 239438 583068 239444 583132
rect 239508 583130 239514 583132
rect 420269 583130 420335 583133
rect 239508 583128 420335 583130
rect 239508 583072 420274 583128
rect 420330 583072 420335 583128
rect 239508 583070 420335 583072
rect 239508 583068 239514 583070
rect 420269 583067 420335 583070
rect 239254 582932 239260 582996
rect 239324 582994 239330 582996
rect 426617 582994 426683 582997
rect 239324 582992 426683 582994
rect 239324 582936 426622 582992
rect 426678 582936 426683 582992
rect 239324 582934 426683 582936
rect 239324 582932 239330 582934
rect 426617 582931 426683 582934
rect 17217 582858 17283 582861
rect 449801 582858 449867 582861
rect 17217 582856 449867 582858
rect 17217 582800 17222 582856
rect 17278 582800 449806 582856
rect 449862 582800 449867 582856
rect 17217 582798 449867 582800
rect 17217 582795 17283 582798
rect 449801 582795 449867 582798
rect 24117 582722 24183 582725
rect 462405 582722 462471 582725
rect 24117 582720 462471 582722
rect 24117 582664 24122 582720
rect 24178 582664 462410 582720
rect 462466 582664 462471 582720
rect 24117 582662 462471 582664
rect 24117 582659 24183 582662
rect 462405 582659 462471 582662
rect 5073 582586 5139 582589
rect 447685 582586 447751 582589
rect 5073 582584 447751 582586
rect 5073 582528 5078 582584
rect 5134 582528 447690 582584
rect 447746 582528 447751 582584
rect 5073 582526 447751 582528
rect 5073 582523 5139 582526
rect 447685 582523 447751 582526
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 465574 579668 465580 579732
rect 465644 579730 465650 579732
rect 468477 579730 468543 579733
rect 465644 579728 468543 579730
rect 465644 579672 468482 579728
rect 468538 579672 468543 579728
rect 465644 579670 468543 579672
rect 465644 579668 465650 579670
rect 468477 579667 468543 579670
rect 231117 579322 231183 579325
rect 232957 579324 233023 579325
rect 231710 579322 231716 579324
rect 231117 579320 231716 579322
rect 231117 579264 231122 579320
rect 231178 579264 231716 579320
rect 231117 579262 231716 579264
rect 231117 579259 231183 579262
rect 231710 579260 231716 579262
rect 231780 579260 231786 579324
rect 232957 579320 233004 579324
rect 233068 579322 233074 579324
rect 235257 579322 235323 579325
rect 237189 579324 237255 579325
rect 235758 579322 235764 579324
rect 232957 579264 232962 579320
rect 232957 579260 233004 579264
rect 233068 579262 233114 579322
rect 235257 579320 235764 579322
rect 235257 579264 235262 579320
rect 235318 579264 235764 579320
rect 235257 579262 235764 579264
rect 233068 579260 233074 579262
rect 232957 579259 233023 579260
rect 235257 579259 235323 579262
rect 235758 579260 235764 579262
rect 235828 579260 235834 579324
rect 237189 579320 237236 579324
rect 237300 579322 237306 579324
rect 239397 579322 239463 579325
rect 239990 579322 239996 579324
rect 237189 579264 237194 579320
rect 237189 579260 237236 579264
rect 237300 579262 237346 579322
rect 239397 579320 239996 579322
rect 239397 579264 239402 579320
rect 239458 579264 239996 579320
rect 239397 579262 239996 579264
rect 237300 579260 237306 579262
rect 237189 579259 237255 579260
rect 239397 579259 239463 579262
rect 239990 579260 239996 579262
rect 240060 579260 240066 579324
rect 241278 579260 241284 579324
rect 241348 579322 241354 579324
rect 241421 579322 241487 579325
rect 241348 579320 241487 579322
rect 241348 579264 241426 579320
rect 241482 579264 241487 579320
rect 241348 579262 241487 579264
rect 241348 579260 241354 579262
rect 241421 579259 241487 579262
rect 249517 579324 249583 579325
rect 466453 579324 466519 579325
rect 249517 579320 249564 579324
rect 249628 579322 249634 579324
rect 249517 579264 249522 579320
rect 249517 579260 249564 579264
rect 249628 579262 249674 579322
rect 466453 579320 466500 579324
rect 466564 579322 466570 579324
rect 466453 579264 466458 579320
rect 249628 579260 249634 579262
rect 466453 579260 466500 579264
rect 466564 579262 466610 579322
rect 466564 579260 466570 579262
rect 249517 579259 249583 579260
rect 466453 579259 466519 579260
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3049 567354 3115 567357
rect -960 567352 3115 567354
rect -960 567296 3054 567352
rect 3110 567296 3115 567352
rect -960 567294 3115 567296
rect -960 567204 480 567294
rect 3049 567291 3115 567294
rect 579705 557290 579771 557293
rect 583520 557290 584960 557380
rect 579705 557288 584960 557290
rect 579705 557232 579710 557288
rect 579766 557232 584960 557288
rect 579705 557230 584960 557232
rect 579705 557227 579771 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 2773 553074 2839 553077
rect -960 553072 2839 553074
rect -960 553016 2778 553072
rect 2834 553016 2839 553072
rect -960 553014 2839 553016
rect -960 552924 480 553014
rect 2773 553011 2839 553014
rect 579705 545594 579771 545597
rect 583520 545594 584960 545684
rect 579705 545592 584960 545594
rect 579705 545536 579710 545592
rect 579766 545536 584960 545592
rect 579705 545534 584960 545536
rect 579705 545531 579771 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3049 538658 3115 538661
rect -960 538656 3115 538658
rect -960 538600 3054 538656
rect 3110 538600 3115 538656
rect -960 538598 3115 538600
rect -960 538508 480 538598
rect 3049 538595 3115 538598
rect 583520 533898 584960 533988
rect 583342 533838 584960 533898
rect 465942 533020 465948 533084
rect 466012 533082 466018 533084
rect 466012 533022 470610 533082
rect 466012 533020 466018 533022
rect 470550 532946 470610 533022
rect 480302 533022 489930 533082
rect 470550 532886 480178 532946
rect 480118 532810 480178 532886
rect 480302 532810 480362 533022
rect 489870 532946 489930 533022
rect 499622 533022 509250 533082
rect 489870 532886 499498 532946
rect 480118 532750 480362 532810
rect 499438 532810 499498 532886
rect 499622 532810 499682 533022
rect 509190 532946 509250 533022
rect 518942 533022 528570 533082
rect 509190 532886 518818 532946
rect 499438 532750 499682 532810
rect 518758 532810 518818 532886
rect 518942 532810 519002 533022
rect 528510 532946 528570 533022
rect 538262 533022 547890 533082
rect 528510 532886 538138 532946
rect 518758 532750 519002 532810
rect 538078 532810 538138 532886
rect 538262 532810 538322 533022
rect 547830 532946 547890 533022
rect 557582 533022 567210 533082
rect 547830 532886 557458 532946
rect 538078 532750 538322 532810
rect 557398 532810 557458 532886
rect 557582 532810 557642 533022
rect 567150 532946 567210 533022
rect 583342 532946 583402 533838
rect 583520 533748 584960 533838
rect 567150 532886 576778 532946
rect 557398 532750 557642 532810
rect 576718 532810 576778 532886
rect 576902 532886 583402 532946
rect 576902 532810 576962 532886
rect 576718 532750 576962 532810
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579705 510370 579771 510373
rect 583520 510370 584960 510460
rect 579705 510368 584960 510370
rect 579705 510312 579710 510368
rect 579766 510312 584960 510368
rect 579705 510310 584960 510312
rect 579705 510307 579771 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3049 509962 3115 509965
rect -960 509960 3115 509962
rect -960 509904 3054 509960
rect 3110 509904 3115 509960
rect -960 509902 3115 509904
rect -960 509812 480 509902
rect 3049 509899 3115 509902
rect 579705 498674 579771 498677
rect 583520 498674 584960 498764
rect 579705 498672 584960 498674
rect 579705 498616 579710 498672
rect 579766 498616 584960 498672
rect 579705 498614 584960 498616
rect 579705 498611 579771 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 583520 486842 584960 486932
rect 583342 486782 584960 486842
rect 465758 486100 465764 486164
rect 465828 486162 465834 486164
rect 465828 486102 470610 486162
rect 465828 486100 465834 486102
rect 470550 486026 470610 486102
rect 480302 486102 489930 486162
rect 470550 485966 480178 486026
rect 480118 485890 480178 485966
rect 480302 485890 480362 486102
rect 489870 486026 489930 486102
rect 499622 486102 509250 486162
rect 489870 485966 499498 486026
rect 480118 485830 480362 485890
rect 499438 485890 499498 485966
rect 499622 485890 499682 486102
rect 509190 486026 509250 486102
rect 518942 486102 528570 486162
rect 509190 485966 518818 486026
rect 499438 485830 499682 485890
rect 518758 485890 518818 485966
rect 518942 485890 519002 486102
rect 528510 486026 528570 486102
rect 538262 486102 547890 486162
rect 528510 485966 538138 486026
rect 518758 485830 519002 485890
rect 538078 485890 538138 485966
rect 538262 485890 538322 486102
rect 547830 486026 547890 486102
rect 557582 486102 567210 486162
rect 547830 485966 557458 486026
rect 538078 485830 538322 485890
rect 557398 485890 557458 485966
rect 557582 485890 557642 486102
rect 567150 486026 567210 486102
rect 583342 486026 583402 486782
rect 583520 486692 584960 486782
rect 567150 485966 576778 486026
rect 557398 485830 557642 485890
rect 576718 485890 576778 485966
rect 576902 485966 583402 486026
rect 576902 485890 576962 485966
rect 576718 485830 576962 485890
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579705 463450 579771 463453
rect 583520 463450 584960 463540
rect 579705 463448 584960 463450
rect 579705 463392 579710 463448
rect 579766 463392 584960 463448
rect 579705 463390 584960 463392
rect 579705 463387 579771 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3141 452434 3207 452437
rect -960 452432 3207 452434
rect -960 452376 3146 452432
rect 3202 452376 3207 452432
rect -960 452374 3207 452376
rect -960 452284 480 452374
rect 3141 452371 3207 452374
rect 579797 451754 579863 451757
rect 583520 451754 584960 451844
rect 579797 451752 584960 451754
rect 579797 451696 579802 451752
rect 579858 451696 584960 451752
rect 579797 451694 584960 451696
rect 579797 451691 579863 451694
rect 583520 451604 584960 451694
rect 579797 439922 579863 439925
rect 583520 439922 584960 440012
rect 579797 439920 584960 439922
rect 579797 439864 579802 439920
rect 579858 439864 584960 439920
rect 579797 439862 584960 439864
rect 579797 439859 579863 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3141 423738 3207 423741
rect -960 423736 3207 423738
rect -960 423680 3146 423736
rect 3202 423680 3207 423736
rect -960 423678 3207 423680
rect -960 423588 480 423678
rect 3141 423675 3207 423678
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579797 404834 579863 404837
rect 583520 404834 584960 404924
rect 579797 404832 584960 404834
rect 579797 404776 579802 404832
rect 579858 404776 584960 404832
rect 579797 404774 584960 404776
rect 579797 404771 579863 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3233 395042 3299 395045
rect -960 395040 3299 395042
rect -960 394984 3238 395040
rect 3294 394984 3299 395040
rect -960 394982 3299 394984
rect -960 394892 480 394982
rect 3233 394979 3299 394982
rect 579797 393002 579863 393005
rect 583520 393002 584960 393092
rect 579797 393000 584960 393002
rect 579797 392944 579802 393000
rect 579858 392944 584960 393000
rect 579797 392942 584960 392944
rect 579797 392939 579863 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 579889 369610 579955 369613
rect 583520 369610 584960 369700
rect 579889 369608 584960 369610
rect 579889 369552 579894 369608
rect 579950 369552 584960 369608
rect 579889 369550 584960 369552
rect 579889 369547 579955 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3325 366210 3391 366213
rect -960 366208 3391 366210
rect -960 366152 3330 366208
rect 3386 366152 3391 366208
rect -960 366150 3391 366152
rect -960 366060 480 366150
rect 3325 366147 3391 366150
rect 579981 357914 580047 357917
rect 583520 357914 584960 358004
rect 579981 357912 584960 357914
rect 579981 357856 579986 357912
rect 580042 357856 584960 357912
rect 579981 357854 584960 357856
rect 579981 357851 580047 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579981 346082 580047 346085
rect 583520 346082 584960 346172
rect 579981 346080 584960 346082
rect 579981 346024 579986 346080
rect 580042 346024 584960 346080
rect 579981 346022 584960 346024
rect 579981 346019 580047 346022
rect 583520 345932 584960 346022
rect 239438 338058 239444 338060
rect 614 337998 239444 338058
rect -960 337514 480 337604
rect 614 337514 674 337998
rect 239438 337996 239444 337998
rect 239508 337996 239514 338060
rect 483013 338058 483079 338061
rect 483381 338058 483447 338061
rect 483013 338056 483447 338058
rect 483013 338000 483018 338056
rect 483074 338000 483386 338056
rect 483442 338000 483447 338056
rect 483013 337998 483447 338000
rect 483013 337995 483079 337998
rect 483381 337995 483447 337998
rect 483013 337922 483079 337925
rect 483381 337922 483447 337925
rect 483013 337920 483447 337922
rect 483013 337864 483018 337920
rect 483074 337864 483386 337920
rect 483442 337864 483447 337920
rect 483013 337862 483447 337864
rect 483013 337859 483079 337862
rect 483381 337859 483447 337862
rect 57973 337786 58039 337789
rect 67541 337786 67607 337789
rect 57973 337784 67607 337786
rect 57973 337728 57978 337784
rect 58034 337728 67546 337784
rect 67602 337728 67607 337784
rect 57973 337726 67607 337728
rect 57973 337723 58039 337726
rect 67541 337723 67607 337726
rect 455689 337786 455755 337789
rect 463601 337786 463667 337789
rect 455689 337784 463667 337786
rect 455689 337728 455694 337784
rect 455750 337728 463606 337784
rect 463662 337728 463667 337784
rect 455689 337726 463667 337728
rect 455689 337723 455755 337726
rect 463601 337723 463667 337726
rect 483013 337786 483079 337789
rect 483381 337786 483447 337789
rect 483013 337784 483447 337786
rect 483013 337728 483018 337784
rect 483074 337728 483386 337784
rect 483442 337728 483447 337784
rect 483013 337726 483447 337728
rect 483013 337723 483079 337726
rect 483381 337723 483447 337726
rect 307753 337650 307819 337653
rect 317321 337650 317387 337653
rect 307753 337648 317387 337650
rect 307753 337592 307758 337648
rect 307814 337592 317326 337648
rect 317382 337592 317387 337648
rect 307753 337590 317387 337592
rect 307753 337587 307819 337590
rect 317321 337587 317387 337590
rect 483013 337650 483079 337653
rect 483473 337650 483539 337653
rect 483013 337648 483539 337650
rect 483013 337592 483018 337648
rect 483074 337592 483478 337648
rect 483534 337592 483539 337648
rect 483013 337590 483539 337592
rect 483013 337587 483079 337590
rect 483473 337587 483539 337590
rect -960 337454 674 337514
rect 342713 337514 342779 337517
rect 345749 337514 345815 337517
rect 342713 337512 345815 337514
rect 342713 337456 342718 337512
rect 342774 337456 345754 337512
rect 345810 337456 345815 337512
rect 342713 337454 345815 337456
rect -960 337364 480 337454
rect 342713 337451 342779 337454
rect 345749 337451 345815 337454
rect 10317 337378 10383 337381
rect 231945 337378 232011 337381
rect 10317 337376 232011 337378
rect 10317 337320 10322 337376
rect 10378 337320 231950 337376
rect 232006 337320 232011 337376
rect 10317 337318 232011 337320
rect 10317 337315 10383 337318
rect 231945 337315 232011 337318
rect 467557 337378 467623 337381
rect 512637 337378 512703 337381
rect 467557 337376 512703 337378
rect 467557 337320 467562 337376
rect 467618 337320 512642 337376
rect 512698 337320 512703 337376
rect 467557 337318 512703 337320
rect 467557 337315 467623 337318
rect 512637 337315 512703 337318
rect 249149 334250 249215 334253
rect 249374 334250 249380 334252
rect 249149 334248 249380 334250
rect 249149 334192 249154 334248
rect 249210 334192 249380 334248
rect 249149 334190 249380 334192
rect 249149 334187 249215 334190
rect 249374 334188 249380 334190
rect 249444 334188 249450 334252
rect 583520 334236 584960 334476
rect 249149 328538 249215 328541
rect 249149 328536 249258 328538
rect 249149 328480 249154 328536
rect 249210 328504 249258 328536
rect 249374 328504 249380 328506
rect 249210 328480 249380 328504
rect 249149 328475 249380 328480
rect 249198 328444 249380 328475
rect 249374 328442 249380 328444
rect 249444 328442 249450 328506
rect 359181 327314 359247 327317
rect 359046 327312 359247 327314
rect 359046 327256 359186 327312
rect 359242 327256 359247 327312
rect 359046 327254 359247 327256
rect 359046 327178 359106 327254
rect 359181 327251 359247 327254
rect 359181 327178 359247 327181
rect 359046 327176 359247 327178
rect 359046 327120 359186 327176
rect 359242 327120 359247 327176
rect 359046 327118 359247 327120
rect 359181 327115 359247 327118
rect 386781 325954 386847 325957
rect 386646 325952 386847 325954
rect 386646 325896 386786 325952
rect 386842 325896 386847 325952
rect 386646 325894 386847 325896
rect 386646 325818 386706 325894
rect 386781 325891 386847 325894
rect 386781 325818 386847 325821
rect 386646 325816 386847 325818
rect 386646 325760 386786 325816
rect 386842 325760 386847 325816
rect 386646 325758 386847 325760
rect 386781 325755 386847 325758
rect 270493 325682 270559 325685
rect 270769 325682 270835 325685
rect 270493 325680 270835 325682
rect 270493 325624 270498 325680
rect 270554 325624 270774 325680
rect 270830 325624 270835 325680
rect 270493 325622 270835 325624
rect 270493 325619 270559 325622
rect 270769 325619 270835 325622
rect 386781 325682 386847 325685
rect 386965 325682 387031 325685
rect 386781 325680 387031 325682
rect 386781 325624 386786 325680
rect 386842 325624 386970 325680
rect 387026 325624 387031 325680
rect 386781 325622 387031 325624
rect 386781 325619 386847 325622
rect 386965 325619 387031 325622
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 579981 322690 580047 322693
rect 583520 322690 584960 322780
rect 579981 322688 584960 322690
rect 579981 322632 579986 322688
rect 580042 322632 584960 322688
rect 579981 322630 584960 322632
rect 579981 322627 580047 322630
rect 583520 322540 584960 322630
rect 249149 322282 249215 322285
rect 249374 322282 249380 322284
rect 249149 322280 249380 322282
rect 249149 322224 249154 322280
rect 249210 322224 249380 322280
rect 249149 322222 249380 322224
rect 249149 322219 249215 322222
rect 249374 322220 249380 322222
rect 249444 322220 249450 322284
rect 460013 318882 460079 318885
rect 460197 318882 460263 318885
rect 460013 318880 460263 318882
rect 460013 318824 460018 318880
rect 460074 318824 460202 318880
rect 460258 318824 460263 318880
rect 460013 318822 460263 318824
rect 460013 318819 460079 318822
rect 460197 318819 460263 318822
rect 249149 317658 249215 317661
rect 249014 317656 249215 317658
rect 249014 317600 249154 317656
rect 249210 317600 249215 317656
rect 249014 317598 249215 317600
rect 249014 317524 249074 317598
rect 249149 317595 249215 317598
rect 249006 317460 249012 317524
rect 249076 317460 249082 317524
rect 301313 317522 301379 317525
rect 301086 317520 301379 317522
rect 301086 317464 301318 317520
rect 301374 317464 301379 317520
rect 301086 317462 301379 317464
rect 301086 317386 301146 317462
rect 301313 317459 301379 317462
rect 301221 317386 301287 317389
rect 301086 317384 301287 317386
rect 301086 317328 301226 317384
rect 301282 317328 301287 317384
rect 301086 317326 301287 317328
rect 301221 317323 301287 317326
rect 330201 316026 330267 316029
rect 330385 316026 330451 316029
rect 330201 316024 330451 316026
rect 330201 315968 330206 316024
rect 330262 315968 330390 316024
rect 330446 315968 330451 316024
rect 330201 315966 330451 315968
rect 330201 315963 330267 315966
rect 330385 315963 330451 315966
rect 270677 314666 270743 314669
rect 270861 314666 270927 314669
rect 270677 314664 270927 314666
rect 270677 314608 270682 314664
rect 270738 314608 270866 314664
rect 270922 314608 270927 314664
rect 270677 314606 270927 314608
rect 270677 314603 270743 314606
rect 270861 314603 270927 314606
rect 580073 310858 580139 310861
rect 583520 310858 584960 310948
rect 580073 310856 584960 310858
rect 580073 310800 580078 310856
rect 580134 310800 584960 310856
rect 580073 310798 584960 310800
rect 580073 310795 580139 310798
rect 583520 310708 584960 310798
rect 236269 309362 236335 309365
rect 236134 309360 236335 309362
rect 236134 309304 236274 309360
rect 236330 309304 236335 309360
rect 236134 309302 236335 309304
rect 236134 309226 236194 309302
rect 236269 309299 236335 309302
rect 236269 309226 236335 309229
rect 236134 309224 236335 309226
rect 236134 309168 236274 309224
rect 236330 309168 236335 309224
rect 236134 309166 236335 309168
rect 236269 309163 236335 309166
rect 249006 309164 249012 309228
rect 249076 309164 249082 309228
rect 375557 309226 375623 309229
rect 375741 309226 375807 309229
rect 375557 309224 375807 309226
rect 375557 309168 375562 309224
rect 375618 309168 375746 309224
rect 375802 309168 375807 309224
rect 375557 309166 375807 309168
rect 249014 308954 249074 309164
rect 375557 309163 375623 309166
rect 375741 309163 375807 309166
rect 249190 308954 249196 308956
rect -960 308818 480 308908
rect 249014 308894 249196 308954
rect 249190 308892 249196 308894
rect 249260 308892 249266 308956
rect 2773 308818 2839 308821
rect -960 308816 2839 308818
rect -960 308760 2778 308816
rect 2834 308760 2839 308816
rect -960 308758 2839 308760
rect -960 308668 480 308758
rect 2773 308755 2839 308758
rect 291469 306370 291535 306373
rect 291745 306370 291811 306373
rect 291469 306368 291811 306370
rect 291469 306312 291474 306368
rect 291530 306312 291750 306368
rect 291806 306312 291811 306368
rect 291469 306310 291811 306312
rect 291469 306307 291535 306310
rect 291745 306307 291811 306310
rect 249190 302228 249196 302292
rect 249260 302228 249266 302292
rect 249198 302156 249258 302228
rect 249190 302092 249196 302156
rect 249260 302092 249266 302156
rect 341241 299434 341307 299437
rect 341374 299434 341380 299436
rect 341241 299432 341380 299434
rect 341241 299376 341246 299432
rect 341302 299376 341380 299432
rect 341241 299374 341380 299376
rect 341241 299371 341307 299374
rect 341374 299372 341380 299374
rect 341444 299372 341450 299436
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 325601 298210 325667 298213
rect 325601 298208 325802 298210
rect 325601 298152 325606 298208
rect 325662 298176 325802 298208
rect 325877 298176 325943 298179
rect 325662 298174 325943 298176
rect 325662 298152 325882 298174
rect 325601 298150 325882 298152
rect 325601 298147 325667 298150
rect 325742 298118 325882 298150
rect 325938 298118 325943 298174
rect 325742 298116 325943 298118
rect 325877 298113 325943 298116
rect 249241 298076 249307 298077
rect 249190 298074 249196 298076
rect 249150 298014 249196 298074
rect 249260 298072 249307 298076
rect 249302 298016 249307 298072
rect 249190 298012 249196 298014
rect 249260 298012 249307 298016
rect 249241 298011 249307 298012
rect 325877 296714 325943 296717
rect 326061 296714 326127 296717
rect 325877 296712 326127 296714
rect 325877 296656 325882 296712
rect 325938 296656 326066 296712
rect 326122 296656 326127 296712
rect 325877 296654 326127 296656
rect 325877 296651 325943 296654
rect 326061 296651 326127 296654
rect 2957 295218 3023 295221
rect 239254 295218 239260 295220
rect 2957 295216 239260 295218
rect 2957 295160 2962 295216
rect 3018 295160 239260 295216
rect 2957 295158 239260 295160
rect 2957 295155 3023 295158
rect 239254 295156 239260 295158
rect 239324 295156 239330 295220
rect -960 294402 480 294492
rect 2957 294402 3023 294405
rect -960 294400 3023 294402
rect -960 294344 2962 294400
rect 3018 294344 3023 294400
rect -960 294342 3023 294344
rect -960 294252 480 294342
rect 2957 294339 3023 294342
rect 341241 289914 341307 289917
rect 341374 289914 341380 289916
rect 341241 289912 341380 289914
rect 341241 289856 341246 289912
rect 341302 289856 341380 289912
rect 341241 289854 341380 289856
rect 341241 289851 341307 289854
rect 341374 289852 341380 289854
rect 341444 289852 341450 289916
rect 249241 288554 249307 288557
rect 249374 288554 249380 288556
rect 249241 288552 249380 288554
rect 249241 288496 249246 288552
rect 249302 288496 249380 288552
rect 249241 288494 249380 288496
rect 249241 288491 249307 288494
rect 249374 288492 249380 288494
rect 249444 288492 249450 288556
rect 249241 288418 249307 288421
rect 249374 288418 249380 288420
rect 249241 288416 249380 288418
rect 249241 288360 249246 288416
rect 249302 288360 249380 288416
rect 249241 288358 249380 288360
rect 249241 288355 249307 288358
rect 249374 288356 249380 288358
rect 249444 288356 249450 288420
rect 250069 288418 250135 288421
rect 250345 288418 250411 288421
rect 250069 288416 250411 288418
rect 250069 288360 250074 288416
rect 250130 288360 250350 288416
rect 250406 288360 250411 288416
rect 250069 288358 250411 288360
rect 250069 288355 250135 288358
rect 250345 288355 250411 288358
rect 323209 288418 323275 288421
rect 323485 288418 323551 288421
rect 323209 288416 323551 288418
rect 323209 288360 323214 288416
rect 323270 288360 323490 288416
rect 323546 288360 323551 288416
rect 323209 288358 323551 288360
rect 323209 288355 323275 288358
rect 323485 288355 323551 288358
rect 583520 287316 584960 287556
rect 259545 280258 259611 280261
rect 259913 280258 259979 280261
rect 259545 280256 259979 280258
rect -960 280122 480 280212
rect 259545 280200 259550 280256
rect 259606 280200 259918 280256
rect 259974 280200 259979 280256
rect 259545 280198 259979 280200
rect 259545 280195 259611 280198
rect 259913 280195 259979 280198
rect 4061 280122 4127 280125
rect -960 280120 4127 280122
rect -960 280064 4066 280120
rect 4122 280064 4127 280120
rect -960 280062 4127 280064
rect -960 279972 480 280062
rect 4061 280059 4127 280062
rect 341241 280122 341307 280125
rect 341374 280122 341380 280124
rect 341241 280120 341380 280122
rect 341241 280064 341246 280120
rect 341302 280064 341380 280120
rect 341241 280062 341380 280064
rect 341241 280059 341307 280062
rect 341374 280060 341380 280062
rect 341444 280060 341450 280124
rect 249241 279036 249307 279037
rect 249190 279034 249196 279036
rect 249150 278974 249196 279034
rect 249260 279032 249307 279036
rect 249302 278976 249307 279032
rect 249190 278972 249196 278974
rect 249260 278972 249307 278976
rect 249241 278971 249307 278972
rect 267733 278762 267799 278765
rect 284569 278762 284635 278765
rect 284753 278762 284819 278765
rect 267733 278760 267842 278762
rect 267733 278704 267738 278760
rect 267794 278704 267842 278760
rect 267733 278699 267842 278704
rect 284569 278760 284819 278762
rect 284569 278704 284574 278760
rect 284630 278704 284758 278760
rect 284814 278704 284819 278760
rect 284569 278702 284819 278704
rect 284569 278699 284635 278702
rect 284753 278699 284819 278702
rect 358537 278762 358603 278765
rect 358721 278762 358787 278765
rect 358537 278760 358787 278762
rect 358537 278704 358542 278760
rect 358598 278704 358726 278760
rect 358782 278704 358787 278760
rect 358537 278702 358787 278704
rect 358537 278699 358603 278702
rect 358721 278699 358787 278702
rect 421189 278762 421255 278765
rect 421373 278762 421439 278765
rect 421189 278760 421439 278762
rect 421189 278704 421194 278760
rect 421250 278704 421378 278760
rect 421434 278704 421439 278760
rect 421189 278702 421439 278704
rect 421189 278699 421255 278702
rect 421373 278699 421439 278702
rect 267782 278629 267842 278699
rect 267782 278624 267891 278629
rect 267782 278568 267830 278624
rect 267886 278568 267891 278624
rect 267782 278566 267891 278568
rect 267825 278563 267891 278566
rect 249190 277340 249196 277404
rect 249260 277402 249266 277404
rect 249425 277402 249491 277405
rect 249260 277400 249491 277402
rect 249260 277344 249430 277400
rect 249486 277344 249491 277400
rect 249260 277342 249491 277344
rect 249260 277340 249266 277342
rect 249425 277339 249491 277342
rect 295609 276042 295675 276045
rect 295793 276042 295859 276045
rect 295609 276040 295859 276042
rect 295609 275984 295614 276040
rect 295670 275984 295798 276040
rect 295854 275984 295859 276040
rect 295609 275982 295859 275984
rect 295609 275979 295675 275982
rect 295793 275979 295859 275982
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 336958 273940 336964 274004
rect 337028 274002 337034 274004
rect 337101 274002 337167 274005
rect 337028 274000 337167 274002
rect 337028 273944 337106 274000
rect 337162 273944 337167 274000
rect 337028 273942 337167 273944
rect 337028 273940 337034 273942
rect 337101 273939 337167 273942
rect 341241 270602 341307 270605
rect 341374 270602 341380 270604
rect 341241 270600 341380 270602
rect 341241 270544 341246 270600
rect 341302 270544 341380 270600
rect 341241 270542 341380 270544
rect 341241 270539 341307 270542
rect 341374 270540 341380 270542
rect 341444 270540 341450 270604
rect 236269 270468 236335 270469
rect 236269 270466 236316 270468
rect 236224 270464 236316 270466
rect 236224 270408 236274 270464
rect 236224 270406 236316 270408
rect 236269 270404 236316 270406
rect 236380 270404 236386 270468
rect 236269 270403 236335 270404
rect 272057 269106 272123 269109
rect 272241 269106 272307 269109
rect 272057 269104 272307 269106
rect 272057 269048 272062 269104
rect 272118 269048 272246 269104
rect 272302 269048 272307 269104
rect 272057 269046 272307 269048
rect 272057 269043 272123 269046
rect 272241 269043 272307 269046
rect 323301 269106 323367 269109
rect 324681 269106 324747 269109
rect 324865 269106 324931 269109
rect 323301 269104 323410 269106
rect 323301 269048 323306 269104
rect 323362 269048 323410 269104
rect 323301 269043 323410 269048
rect 324681 269104 324931 269106
rect 324681 269048 324686 269104
rect 324742 269048 324870 269104
rect 324926 269048 324931 269104
rect 324681 269046 324931 269048
rect 324681 269043 324747 269046
rect 324865 269043 324931 269046
rect 323350 268973 323410 269043
rect 323350 268968 323459 268973
rect 323350 268912 323398 268968
rect 323454 268912 323459 268968
rect 323350 268910 323459 268912
rect 323393 268907 323459 268910
rect 249425 267884 249491 267885
rect 249374 267820 249380 267884
rect 249444 267882 249491 267884
rect 249444 267880 249536 267882
rect 249486 267824 249536 267880
rect 249444 267822 249536 267824
rect 249444 267820 249491 267822
rect 249425 267819 249491 267820
rect -960 265706 480 265796
rect 3969 265706 4035 265709
rect -960 265704 4035 265706
rect -960 265648 3974 265704
rect 4030 265648 4035 265704
rect -960 265646 4035 265648
rect -960 265556 480 265646
rect 3969 265643 4035 265646
rect 580901 263938 580967 263941
rect 583520 263938 584960 264028
rect 580901 263936 584960 263938
rect 580901 263880 580906 263936
rect 580962 263880 584960 263936
rect 580901 263878 584960 263880
rect 580901 263875 580967 263878
rect 249374 263802 249380 263804
rect 249198 263742 249380 263802
rect 249198 263532 249258 263742
rect 249374 263740 249380 263742
rect 249444 263740 249450 263804
rect 583520 263788 584960 263878
rect 249190 263468 249196 263532
rect 249260 263468 249266 263532
rect 286041 261082 286107 261085
rect 285814 261080 286107 261082
rect 285814 261024 286046 261080
rect 286102 261024 286107 261080
rect 285814 261022 286107 261024
rect 236310 260884 236316 260948
rect 236380 260946 236386 260948
rect 236453 260946 236519 260949
rect 236380 260944 236519 260946
rect 236380 260888 236458 260944
rect 236514 260888 236519 260944
rect 236380 260886 236519 260888
rect 285814 260946 285874 261022
rect 286041 261019 286107 261022
rect 285949 260946 286015 260949
rect 285814 260944 286015 260946
rect 285814 260888 285954 260944
rect 286010 260888 286015 260944
rect 285814 260886 286015 260888
rect 236380 260884 236386 260886
rect 236453 260883 236519 260886
rect 285949 260883 286015 260886
rect 341241 260810 341307 260813
rect 341374 260810 341380 260812
rect 341241 260808 341380 260810
rect 341241 260752 341246 260808
rect 341302 260752 341380 260808
rect 341241 260750 341380 260752
rect 341241 260747 341307 260750
rect 341374 260748 341380 260750
rect 341444 260748 341450 260812
rect 336917 260676 336983 260677
rect 336917 260672 336964 260676
rect 337028 260674 337034 260676
rect 336917 260616 336922 260672
rect 336917 260612 336964 260616
rect 337028 260614 337074 260674
rect 337028 260612 337034 260614
rect 336917 260611 336983 260612
rect 244457 259450 244523 259453
rect 244641 259450 244707 259453
rect 244457 259448 244707 259450
rect 244457 259392 244462 259448
rect 244518 259392 244646 259448
rect 244702 259392 244707 259448
rect 244457 259390 244707 259392
rect 244457 259387 244523 259390
rect 244641 259387 244707 259390
rect 272149 259450 272215 259453
rect 272425 259450 272491 259453
rect 272149 259448 272491 259450
rect 272149 259392 272154 259448
rect 272210 259392 272430 259448
rect 272486 259392 272491 259448
rect 272149 259390 272491 259392
rect 272149 259387 272215 259390
rect 272425 259387 272491 259390
rect 421189 259450 421255 259453
rect 421373 259450 421439 259453
rect 421189 259448 421439 259450
rect 421189 259392 421194 259448
rect 421250 259392 421378 259448
rect 421434 259392 421439 259448
rect 421189 259390 421439 259392
rect 421189 259387 421255 259390
rect 421373 259387 421439 259390
rect 288801 258226 288867 258229
rect 288758 258224 288867 258226
rect 288758 258168 288806 258224
rect 288862 258168 288867 258224
rect 288758 258163 288867 258168
rect 288758 258093 288818 258163
rect 288758 258088 288867 258093
rect 288758 258032 288806 258088
rect 288862 258032 288867 258088
rect 288758 258030 288867 258032
rect 288801 258027 288867 258030
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 2773 251290 2839 251293
rect -960 251288 2839 251290
rect -960 251232 2778 251288
rect 2834 251232 2839 251288
rect -960 251230 2839 251232
rect -960 251140 480 251230
rect 2773 251227 2839 251230
rect 341241 251290 341307 251293
rect 341374 251290 341380 251292
rect 341241 251288 341380 251290
rect 341241 251232 341246 251288
rect 341302 251232 341380 251288
rect 341241 251230 341380 251232
rect 341241 251227 341307 251230
rect 341374 251228 341380 251230
rect 341444 251228 341450 251292
rect 236269 251154 236335 251157
rect 236545 251154 236611 251157
rect 236269 251152 236611 251154
rect 236269 251096 236274 251152
rect 236330 251096 236550 251152
rect 236606 251096 236611 251152
rect 236269 251094 236611 251096
rect 236269 251091 236335 251094
rect 236545 251091 236611 251094
rect 286041 249794 286107 249797
rect 285998 249792 286107 249794
rect 285998 249736 286046 249792
rect 286102 249736 286107 249792
rect 285998 249731 286107 249736
rect 330201 249794 330267 249797
rect 330385 249794 330451 249797
rect 330201 249792 330451 249794
rect 330201 249736 330206 249792
rect 330262 249736 330390 249792
rect 330446 249736 330451 249792
rect 330201 249734 330451 249736
rect 330201 249731 330267 249734
rect 330385 249731 330451 249734
rect 285998 249661 286058 249731
rect 285949 249656 286058 249661
rect 285949 249600 285954 249656
rect 286010 249600 286058 249656
rect 285949 249598 286058 249600
rect 285949 249595 286015 249598
rect 267733 248434 267799 248437
rect 268009 248434 268075 248437
rect 267733 248432 268075 248434
rect 267733 248376 267738 248432
rect 267794 248376 268014 248432
rect 268070 248376 268075 248432
rect 267733 248374 268075 248376
rect 267733 248371 267799 248374
rect 268009 248371 268075 248374
rect 262489 247074 262555 247077
rect 295517 247074 295583 247077
rect 295885 247074 295951 247077
rect 262489 247072 262874 247074
rect 262489 247016 262494 247072
rect 262550 247016 262874 247072
rect 262489 247014 262874 247016
rect 262489 247011 262555 247014
rect 262814 246941 262874 247014
rect 295517 247072 295951 247074
rect 295517 247016 295522 247072
rect 295578 247016 295890 247072
rect 295946 247016 295951 247072
rect 295517 247014 295951 247016
rect 295517 247011 295583 247014
rect 295885 247011 295951 247014
rect 262765 246936 262874 246941
rect 262765 246880 262770 246936
rect 262826 246880 262874 246936
rect 262765 246878 262874 246880
rect 262765 246875 262831 246878
rect 249374 241906 249380 241908
rect 249198 241846 249380 241906
rect 249198 241772 249258 241846
rect 249374 241844 249380 241846
rect 249444 241844 249450 241908
rect 249190 241708 249196 241772
rect 249260 241708 249266 241772
rect 421189 241770 421255 241773
rect 421054 241768 421255 241770
rect 421054 241712 421194 241768
rect 421250 241712 421255 241768
rect 421054 241710 421255 241712
rect 421054 241634 421114 241710
rect 421189 241707 421255 241710
rect 421189 241634 421255 241637
rect 421054 241632 421255 241634
rect 421054 241576 421194 241632
rect 421250 241576 421255 241632
rect 421054 241574 421255 241576
rect 421189 241571 421255 241574
rect 244273 241498 244339 241501
rect 244457 241498 244523 241501
rect 244273 241496 244523 241498
rect 244273 241440 244278 241496
rect 244334 241440 244462 241496
rect 244518 241440 244523 241496
rect 244273 241438 244523 241440
rect 244273 241435 244339 241438
rect 244457 241435 244523 241438
rect 249190 241436 249196 241500
rect 249260 241436 249266 241500
rect 251449 241498 251515 241501
rect 251633 241498 251699 241501
rect 251449 241496 251699 241498
rect 251449 241440 251454 241496
rect 251510 241440 251638 241496
rect 251694 241440 251699 241496
rect 251449 241438 251699 241440
rect 249198 240954 249258 241436
rect 251449 241435 251515 241438
rect 251633 241435 251699 241438
rect 301037 241498 301103 241501
rect 372521 241498 372587 241501
rect 372705 241498 372771 241501
rect 301037 241496 301146 241498
rect 301037 241440 301042 241496
rect 301098 241440 301146 241496
rect 301037 241435 301146 241440
rect 372521 241496 372771 241498
rect 372521 241440 372526 241496
rect 372582 241440 372710 241496
rect 372766 241440 372771 241496
rect 372521 241438 372771 241440
rect 372521 241435 372587 241438
rect 372705 241435 372771 241438
rect 376937 241498 377003 241501
rect 377121 241498 377187 241501
rect 376937 241496 377187 241498
rect 376937 241440 376942 241496
rect 376998 241440 377126 241496
rect 377182 241440 377187 241496
rect 376937 241438 377187 241440
rect 376937 241435 377003 241438
rect 377121 241435 377187 241438
rect 301086 241365 301146 241435
rect 301086 241360 301195 241365
rect 301086 241304 301134 241360
rect 301190 241304 301195 241360
rect 301086 241302 301195 241304
rect 301129 241299 301195 241302
rect 249374 240954 249380 240956
rect 249198 240894 249380 240954
rect 249374 240892 249380 240894
rect 249444 240892 249450 240956
rect 583520 240396 584960 240636
rect 325877 240138 325943 240141
rect 326153 240138 326219 240141
rect 325877 240136 326219 240138
rect 325877 240080 325882 240136
rect 325938 240080 326158 240136
rect 326214 240080 326219 240136
rect 325877 240078 326219 240080
rect 325877 240075 325943 240078
rect 326153 240075 326219 240078
rect 336733 240138 336799 240141
rect 336917 240138 336983 240141
rect 336733 240136 336983 240138
rect 336733 240080 336738 240136
rect 336794 240080 336922 240136
rect 336978 240080 336983 240136
rect 336733 240078 336983 240080
rect 336733 240075 336799 240078
rect 336917 240075 336983 240078
rect 341149 240138 341215 240141
rect 341425 240138 341491 240141
rect 341149 240136 341491 240138
rect 341149 240080 341154 240136
rect 341210 240080 341430 240136
rect 341486 240080 341491 240136
rect 341149 240078 341491 240080
rect 341149 240075 341215 240078
rect 341425 240075 341491 240078
rect 421189 240138 421255 240141
rect 421373 240138 421439 240141
rect 421189 240136 421439 240138
rect 421189 240080 421194 240136
rect 421250 240080 421378 240136
rect 421434 240080 421439 240136
rect 421189 240078 421439 240080
rect 421189 240075 421255 240078
rect 421373 240075 421439 240078
rect 459829 240138 459895 240141
rect 460013 240138 460079 240141
rect 459829 240136 460079 240138
rect 459829 240080 459834 240136
rect 459890 240080 460018 240136
rect 460074 240080 460079 240136
rect 459829 240078 460079 240080
rect 459829 240075 459895 240078
rect 460013 240075 460079 240078
rect -960 237010 480 237100
rect 3049 237010 3115 237013
rect -960 237008 3115 237010
rect -960 236952 3054 237008
rect 3110 236952 3115 237008
rect -960 236950 3115 236952
rect -960 236860 480 236950
rect 3049 236947 3115 236950
rect 236637 232114 236703 232117
rect 236134 232112 236703 232114
rect 236134 232056 236642 232112
rect 236698 232056 236703 232112
rect 236134 232054 236703 232056
rect 236134 231978 236194 232054
rect 236637 232051 236703 232054
rect 236269 231978 236335 231981
rect 236134 231976 236335 231978
rect 236134 231920 236274 231976
rect 236330 231920 236335 231976
rect 236134 231918 236335 231920
rect 236269 231915 236335 231918
rect 386413 231842 386479 231845
rect 386781 231842 386847 231845
rect 386413 231840 386847 231842
rect 386413 231784 386418 231840
rect 386474 231784 386786 231840
rect 386842 231784 386847 231840
rect 386413 231782 386847 231784
rect 386413 231779 386479 231782
rect 386781 231779 386847 231782
rect 463785 231842 463851 231845
rect 463969 231842 464035 231845
rect 463785 231840 464035 231842
rect 463785 231784 463790 231840
rect 463846 231784 463974 231840
rect 464030 231784 464035 231840
rect 463785 231782 464035 231784
rect 463785 231779 463851 231782
rect 463969 231779 464035 231782
rect 470409 231842 470475 231845
rect 470593 231842 470659 231845
rect 470409 231840 470659 231842
rect 470409 231784 470414 231840
rect 470470 231784 470598 231840
rect 470654 231784 470659 231840
rect 470409 231782 470659 231784
rect 470409 231779 470475 231782
rect 470593 231779 470659 231782
rect 327165 230482 327231 230485
rect 327533 230482 327599 230485
rect 327165 230480 327599 230482
rect 327165 230424 327170 230480
rect 327226 230424 327538 230480
rect 327594 230424 327599 230480
rect 327165 230422 327599 230424
rect 327165 230419 327231 230422
rect 327533 230419 327599 230422
rect 271873 229122 271939 229125
rect 272057 229122 272123 229125
rect 271873 229120 272123 229122
rect 271873 229064 271878 229120
rect 271934 229064 272062 229120
rect 272118 229064 272123 229120
rect 271873 229062 272123 229064
rect 271873 229059 271939 229062
rect 272057 229059 272123 229062
rect 580809 228850 580875 228853
rect 583520 228850 584960 228940
rect 580809 228848 584960 228850
rect 580809 228792 580814 228848
rect 580870 228792 584960 228848
rect 580809 228790 584960 228792
rect 580809 228787 580875 228790
rect 583520 228700 584960 228790
rect 249374 224980 249380 225044
rect 249444 224980 249450 225044
rect 249382 224770 249442 224980
rect 249558 224770 249564 224772
rect 249382 224710 249564 224770
rect 249558 224708 249564 224710
rect 249628 224708 249634 224772
rect -960 222594 480 222684
rect 3877 222594 3943 222597
rect -960 222592 3943 222594
rect -960 222536 3882 222592
rect 3938 222536 3943 222592
rect -960 222534 3943 222536
rect -960 222444 480 222534
rect 3877 222531 3943 222534
rect 236453 222186 236519 222189
rect 244273 222186 244339 222189
rect 244457 222186 244523 222189
rect 236453 222184 236562 222186
rect 236453 222128 236458 222184
rect 236514 222128 236562 222184
rect 236453 222123 236562 222128
rect 244273 222184 244523 222186
rect 244273 222128 244278 222184
rect 244334 222128 244462 222184
rect 244518 222128 244523 222184
rect 244273 222126 244523 222128
rect 244273 222123 244339 222126
rect 244457 222123 244523 222126
rect 251449 222186 251515 222189
rect 251633 222186 251699 222189
rect 251449 222184 251699 222186
rect 251449 222128 251454 222184
rect 251510 222128 251638 222184
rect 251694 222128 251699 222184
rect 251449 222126 251699 222128
rect 251449 222123 251515 222126
rect 251633 222123 251699 222126
rect 285949 222186 286015 222189
rect 286133 222186 286199 222189
rect 285949 222184 286199 222186
rect 285949 222128 285954 222184
rect 286010 222128 286138 222184
rect 286194 222128 286199 222184
rect 285949 222126 286199 222128
rect 285949 222123 286015 222126
rect 286133 222123 286199 222126
rect 301037 222186 301103 222189
rect 367001 222188 367067 222189
rect 366950 222186 366956 222188
rect 301037 222184 301146 222186
rect 301037 222128 301042 222184
rect 301098 222128 301146 222184
rect 301037 222123 301146 222128
rect 366910 222126 366956 222186
rect 367020 222184 367067 222188
rect 367062 222128 367067 222184
rect 366950 222124 366956 222126
rect 367020 222124 367067 222128
rect 367001 222123 367067 222124
rect 372521 222186 372587 222189
rect 372705 222186 372771 222189
rect 372521 222184 372771 222186
rect 372521 222128 372526 222184
rect 372582 222128 372710 222184
rect 372766 222128 372771 222184
rect 372521 222126 372771 222128
rect 372521 222123 372587 222126
rect 372705 222123 372771 222126
rect 376937 222186 377003 222189
rect 377121 222186 377187 222189
rect 376937 222184 377187 222186
rect 376937 222128 376942 222184
rect 376998 222128 377126 222184
rect 377182 222128 377187 222184
rect 376937 222126 377187 222128
rect 376937 222123 377003 222126
rect 377121 222123 377187 222126
rect 236310 221988 236316 222052
rect 236380 222050 236386 222052
rect 236502 222050 236562 222123
rect 236380 221990 236562 222050
rect 301086 222053 301146 222123
rect 301086 222048 301195 222053
rect 301086 221992 301134 222048
rect 301190 221992 301195 222048
rect 301086 221990 301195 221992
rect 236380 221988 236386 221990
rect 301129 221987 301195 221990
rect 270677 220826 270743 220829
rect 270953 220826 271019 220829
rect 270677 220824 271019 220826
rect 270677 220768 270682 220824
rect 270738 220768 270958 220824
rect 271014 220768 271019 220824
rect 270677 220766 271019 220768
rect 270677 220763 270743 220766
rect 270953 220763 271019 220766
rect 284661 220826 284727 220829
rect 284845 220826 284911 220829
rect 284661 220824 284911 220826
rect 284661 220768 284666 220824
rect 284722 220768 284850 220824
rect 284906 220768 284911 220824
rect 284661 220766 284911 220768
rect 284661 220763 284727 220766
rect 284845 220763 284911 220766
rect 285949 220826 286015 220829
rect 286133 220826 286199 220829
rect 285949 220824 286199 220826
rect 285949 220768 285954 220824
rect 286010 220768 286138 220824
rect 286194 220768 286199 220824
rect 285949 220766 286199 220768
rect 285949 220763 286015 220766
rect 286133 220763 286199 220766
rect 337101 220826 337167 220829
rect 358721 220826 358787 220829
rect 358854 220826 358860 220828
rect 337101 220824 337210 220826
rect 337101 220768 337106 220824
rect 337162 220768 337210 220824
rect 337101 220763 337210 220768
rect 358721 220824 358860 220826
rect 358721 220768 358726 220824
rect 358782 220768 358860 220824
rect 358721 220766 358860 220768
rect 358721 220763 358787 220766
rect 358854 220764 358860 220766
rect 358924 220764 358930 220828
rect 421189 220826 421255 220829
rect 421373 220826 421439 220829
rect 421189 220824 421439 220826
rect 421189 220768 421194 220824
rect 421250 220768 421378 220824
rect 421434 220768 421439 220824
rect 421189 220766 421439 220768
rect 421189 220763 421255 220766
rect 421373 220763 421439 220766
rect 459829 220826 459895 220829
rect 460013 220826 460079 220829
rect 459829 220824 460079 220826
rect 459829 220768 459834 220824
rect 459890 220768 460018 220824
rect 460074 220768 460079 220824
rect 459829 220766 460079 220768
rect 459829 220763 459895 220766
rect 460013 220763 460079 220766
rect 337150 220693 337210 220763
rect 337150 220688 337259 220693
rect 337150 220632 337198 220688
rect 337254 220632 337259 220688
rect 337150 220630 337259 220632
rect 337193 220627 337259 220630
rect 290365 219602 290431 219605
rect 290046 219600 290431 219602
rect 290046 219544 290370 219600
rect 290426 219544 290431 219600
rect 290046 219542 290431 219544
rect 290046 219469 290106 219542
rect 290365 219539 290431 219542
rect 265341 219466 265407 219469
rect 265525 219466 265591 219469
rect 265341 219464 265591 219466
rect 265341 219408 265346 219464
rect 265402 219408 265530 219464
rect 265586 219408 265591 219464
rect 265341 219406 265591 219408
rect 290046 219464 290155 219469
rect 290046 219408 290094 219464
rect 290150 219408 290155 219464
rect 290046 219406 290155 219408
rect 265341 219403 265407 219406
rect 265525 219403 265591 219406
rect 290089 219403 290155 219406
rect 291653 219466 291719 219469
rect 292021 219466 292087 219469
rect 291653 219464 292087 219466
rect 291653 219408 291658 219464
rect 291714 219408 292026 219464
rect 292082 219408 292087 219464
rect 291653 219406 292087 219408
rect 291653 219403 291719 219406
rect 292021 219403 292087 219406
rect 249190 217364 249196 217428
rect 249260 217426 249266 217428
rect 249558 217426 249564 217428
rect 249260 217366 249564 217426
rect 249260 217364 249266 217366
rect 249558 217364 249564 217366
rect 249628 217364 249634 217428
rect 580717 217018 580783 217021
rect 583520 217018 584960 217108
rect 580717 217016 584960 217018
rect 580717 216960 580722 217016
rect 580778 216960 584960 217016
rect 580717 216958 584960 216960
rect 580717 216955 580783 216958
rect 583520 216868 584960 216958
rect 236269 212668 236335 212669
rect 367001 212668 367067 212669
rect 236269 212666 236316 212668
rect 236224 212664 236316 212666
rect 236224 212608 236274 212664
rect 236224 212606 236316 212608
rect 236269 212604 236316 212606
rect 236380 212604 236386 212668
rect 366950 212666 366956 212668
rect 366910 212606 366956 212666
rect 367020 212664 367067 212668
rect 367062 212608 367067 212664
rect 366950 212604 366956 212606
rect 367020 212604 367067 212608
rect 236269 212603 236335 212604
rect 367001 212603 367067 212604
rect 236269 212530 236335 212533
rect 236545 212530 236611 212533
rect 249241 212532 249307 212533
rect 249190 212530 249196 212532
rect 236269 212528 236611 212530
rect 236269 212472 236274 212528
rect 236330 212472 236550 212528
rect 236606 212472 236611 212528
rect 236269 212470 236611 212472
rect 249150 212470 249196 212530
rect 249260 212528 249307 212532
rect 327257 212530 327323 212533
rect 249302 212472 249307 212528
rect 236269 212467 236335 212470
rect 236545 212467 236611 212470
rect 249190 212468 249196 212470
rect 249260 212468 249307 212472
rect 249241 212467 249307 212468
rect 327214 212528 327323 212530
rect 327214 212472 327262 212528
rect 327318 212472 327323 212528
rect 327214 212467 327323 212472
rect 386413 212530 386479 212533
rect 386597 212530 386663 212533
rect 386413 212528 386663 212530
rect 386413 212472 386418 212528
rect 386474 212472 386602 212528
rect 386658 212472 386663 212528
rect 386413 212470 386663 212472
rect 386413 212467 386479 212470
rect 386597 212467 386663 212470
rect 463785 212530 463851 212533
rect 463969 212530 464035 212533
rect 463785 212528 464035 212530
rect 463785 212472 463790 212528
rect 463846 212472 463974 212528
rect 464030 212472 464035 212528
rect 463785 212470 464035 212472
rect 463785 212467 463851 212470
rect 463969 212467 464035 212470
rect 470409 212530 470475 212533
rect 470593 212530 470659 212533
rect 470409 212528 470659 212530
rect 470409 212472 470414 212528
rect 470470 212472 470598 212528
rect 470654 212472 470659 212528
rect 470409 212470 470659 212472
rect 470409 212467 470475 212470
rect 470593 212467 470659 212470
rect 327214 212394 327274 212467
rect 327349 212394 327415 212397
rect 327214 212392 327415 212394
rect 327214 212336 327354 212392
rect 327410 212336 327415 212392
rect 327214 212334 327415 212336
rect 327349 212331 327415 212334
rect 265157 211170 265223 211173
rect 265341 211170 265407 211173
rect 265157 211168 265407 211170
rect 265157 211112 265162 211168
rect 265218 211112 265346 211168
rect 265402 211112 265407 211168
rect 265157 211110 265407 211112
rect 265157 211107 265223 211110
rect 265341 211107 265407 211110
rect 266629 211170 266695 211173
rect 266813 211170 266879 211173
rect 266629 211168 266879 211170
rect 266629 211112 266634 211168
rect 266690 211112 266818 211168
rect 266874 211112 266879 211168
rect 266629 211110 266879 211112
rect 266629 211107 266695 211110
rect 266813 211107 266879 211110
rect 323301 211170 323367 211173
rect 323485 211170 323551 211173
rect 323301 211168 323551 211170
rect 323301 211112 323306 211168
rect 323362 211112 323490 211168
rect 323546 211112 323551 211168
rect 323301 211110 323551 211112
rect 323301 211107 323367 211110
rect 323485 211107 323551 211110
rect 358721 211170 358787 211173
rect 358854 211170 358860 211172
rect 358721 211168 358860 211170
rect 358721 211112 358726 211168
rect 358782 211112 358860 211168
rect 358721 211110 358860 211112
rect 358721 211107 358787 211110
rect 358854 211108 358860 211110
rect 358924 211108 358930 211172
rect 421189 211170 421255 211173
rect 421373 211170 421439 211173
rect 421189 211168 421439 211170
rect 421189 211112 421194 211168
rect 421250 211112 421378 211168
rect 421434 211112 421439 211168
rect 421189 211110 421439 211112
rect 421189 211107 421255 211110
rect 421373 211107 421439 211110
rect 267733 209810 267799 209813
rect 267917 209810 267983 209813
rect 267733 209808 267983 209810
rect 267733 209752 267738 209808
rect 267794 209752 267922 209808
rect 267978 209752 267983 209808
rect 267733 209750 267983 209752
rect 267733 209747 267799 209750
rect 267917 209747 267983 209750
rect 270769 209810 270835 209813
rect 270953 209810 271019 209813
rect 270769 209808 271019 209810
rect 270769 209752 270774 209808
rect 270830 209752 270958 209808
rect 271014 209752 271019 209808
rect 270769 209750 271019 209752
rect 270769 209747 270835 209750
rect 270953 209747 271019 209750
rect -960 208178 480 208268
rect 3785 208178 3851 208181
rect -960 208176 3851 208178
rect -960 208120 3790 208176
rect 3846 208120 3851 208176
rect -960 208118 3851 208120
rect -960 208028 480 208118
rect 3785 208115 3851 208118
rect 249241 205458 249307 205461
rect 249558 205458 249564 205460
rect 249241 205456 249564 205458
rect 249241 205400 249246 205456
rect 249302 205400 249564 205456
rect 249241 205398 249564 205400
rect 249241 205395 249307 205398
rect 249558 205396 249564 205398
rect 249628 205396 249634 205460
rect 580625 205322 580691 205325
rect 583520 205322 584960 205412
rect 580625 205320 584960 205322
rect 580625 205264 580630 205320
rect 580686 205264 584960 205320
rect 580625 205262 584960 205264
rect 580625 205259 580691 205262
rect 583520 205172 584960 205262
rect 236545 203010 236611 203013
rect 236502 203008 236611 203010
rect 236502 202952 236550 203008
rect 236606 202952 236611 203008
rect 236502 202947 236611 202952
rect 236310 202812 236316 202876
rect 236380 202874 236386 202876
rect 236502 202874 236562 202947
rect 236380 202814 236562 202874
rect 244273 202874 244339 202877
rect 244457 202874 244523 202877
rect 249609 202876 249675 202877
rect 244273 202872 244523 202874
rect 244273 202816 244278 202872
rect 244334 202816 244462 202872
rect 244518 202816 244523 202872
rect 244273 202814 244523 202816
rect 236380 202812 236386 202814
rect 244273 202811 244339 202814
rect 244457 202811 244523 202814
rect 249558 202812 249564 202876
rect 249628 202874 249675 202876
rect 251449 202874 251515 202877
rect 251633 202874 251699 202877
rect 249628 202872 249720 202874
rect 249670 202816 249720 202872
rect 249628 202814 249720 202816
rect 251449 202872 251699 202874
rect 251449 202816 251454 202872
rect 251510 202816 251638 202872
rect 251694 202816 251699 202872
rect 251449 202814 251699 202816
rect 249628 202812 249675 202814
rect 249609 202811 249675 202812
rect 251449 202811 251515 202814
rect 251633 202811 251699 202814
rect 259637 202874 259703 202877
rect 259913 202874 259979 202877
rect 272149 202874 272215 202877
rect 259637 202872 259979 202874
rect 259637 202816 259642 202872
rect 259698 202816 259918 202872
rect 259974 202816 259979 202872
rect 259637 202814 259979 202816
rect 259637 202811 259703 202814
rect 259913 202811 259979 202814
rect 272014 202872 272215 202874
rect 272014 202816 272154 202872
rect 272210 202816 272215 202872
rect 272014 202814 272215 202816
rect 272014 202738 272074 202814
rect 272149 202811 272215 202814
rect 285765 202874 285831 202877
rect 285949 202874 286015 202877
rect 285765 202872 286015 202874
rect 285765 202816 285770 202872
rect 285826 202816 285954 202872
rect 286010 202816 286015 202872
rect 285765 202814 286015 202816
rect 285765 202811 285831 202814
rect 285949 202811 286015 202814
rect 301037 202874 301103 202877
rect 341149 202874 341215 202877
rect 341425 202874 341491 202877
rect 301037 202872 301146 202874
rect 301037 202816 301042 202872
rect 301098 202816 301146 202872
rect 301037 202811 301146 202816
rect 341149 202872 341491 202874
rect 341149 202816 341154 202872
rect 341210 202816 341430 202872
rect 341486 202816 341491 202872
rect 341149 202814 341491 202816
rect 341149 202811 341215 202814
rect 341425 202811 341491 202814
rect 372521 202874 372587 202877
rect 372705 202874 372771 202877
rect 372521 202872 372771 202874
rect 372521 202816 372526 202872
rect 372582 202816 372710 202872
rect 372766 202816 372771 202872
rect 372521 202814 372771 202816
rect 372521 202811 372587 202814
rect 372705 202811 372771 202814
rect 376937 202874 377003 202877
rect 377121 202874 377187 202877
rect 376937 202872 377187 202874
rect 376937 202816 376942 202872
rect 376998 202816 377126 202872
rect 377182 202816 377187 202872
rect 376937 202814 377187 202816
rect 376937 202811 377003 202814
rect 377121 202811 377187 202814
rect 386597 202874 386663 202877
rect 386873 202874 386939 202877
rect 386597 202872 386939 202874
rect 386597 202816 386602 202872
rect 386658 202816 386878 202872
rect 386934 202816 386939 202872
rect 386597 202814 386939 202816
rect 386597 202811 386663 202814
rect 386873 202811 386939 202814
rect 301086 202741 301146 202811
rect 272333 202738 272399 202741
rect 272014 202736 272399 202738
rect 272014 202680 272338 202736
rect 272394 202680 272399 202736
rect 272014 202678 272399 202680
rect 301086 202736 301195 202741
rect 301086 202680 301134 202736
rect 301190 202680 301195 202736
rect 301086 202678 301195 202680
rect 272333 202675 272399 202678
rect 301129 202675 301195 202678
rect 284661 201514 284727 201517
rect 284845 201514 284911 201517
rect 284661 201512 284911 201514
rect 284661 201456 284666 201512
rect 284722 201456 284850 201512
rect 284906 201456 284911 201512
rect 284661 201454 284911 201456
rect 284661 201451 284727 201454
rect 284845 201451 284911 201454
rect 288801 201514 288867 201517
rect 288985 201514 289051 201517
rect 288801 201512 289051 201514
rect 288801 201456 288806 201512
rect 288862 201456 288990 201512
rect 289046 201456 289051 201512
rect 288801 201454 289051 201456
rect 288801 201451 288867 201454
rect 288985 201451 289051 201454
rect 249374 196556 249380 196620
rect 249444 196618 249450 196620
rect 249609 196618 249675 196621
rect 249444 196616 249675 196618
rect 249444 196560 249614 196616
rect 249670 196560 249675 196616
rect 249444 196558 249675 196560
rect 249444 196556 249450 196558
rect 249609 196555 249675 196558
rect -960 193898 480 193988
rect 3693 193898 3759 193901
rect -960 193896 3759 193898
rect -960 193840 3698 193896
rect 3754 193840 3759 193896
rect -960 193838 3759 193840
rect -960 193748 480 193838
rect 3693 193835 3759 193838
rect 583520 193476 584960 193716
rect 236269 193356 236335 193357
rect 236269 193354 236316 193356
rect 236224 193352 236316 193354
rect 236224 193296 236274 193352
rect 236224 193294 236316 193296
rect 236269 193292 236316 193294
rect 236380 193292 236386 193356
rect 236269 193291 236335 193292
rect 236269 193218 236335 193221
rect 236545 193218 236611 193221
rect 236269 193216 236611 193218
rect 236269 193160 236274 193216
rect 236330 193160 236550 193216
rect 236606 193160 236611 193216
rect 236269 193158 236611 193160
rect 236269 193155 236335 193158
rect 236545 193155 236611 193158
rect 284661 193218 284727 193221
rect 284845 193218 284911 193221
rect 284661 193216 284911 193218
rect 284661 193160 284666 193216
rect 284722 193160 284850 193216
rect 284906 193160 284911 193216
rect 284661 193158 284911 193160
rect 284661 193155 284727 193158
rect 284845 193155 284911 193158
rect 310789 193218 310855 193221
rect 311065 193218 311131 193221
rect 310789 193216 311131 193218
rect 310789 193160 310794 193216
rect 310850 193160 311070 193216
rect 311126 193160 311131 193216
rect 310789 193158 311131 193160
rect 310789 193155 310855 193158
rect 311065 193155 311131 193158
rect 323301 193218 323367 193221
rect 323485 193218 323551 193221
rect 323301 193216 323551 193218
rect 323301 193160 323306 193216
rect 323362 193160 323490 193216
rect 323546 193160 323551 193216
rect 323301 193158 323551 193160
rect 323301 193155 323367 193158
rect 323485 193155 323551 193158
rect 360469 193218 360535 193221
rect 360653 193218 360719 193221
rect 360469 193216 360719 193218
rect 360469 193160 360474 193216
rect 360530 193160 360658 193216
rect 360714 193160 360719 193216
rect 360469 193158 360719 193160
rect 360469 193155 360535 193158
rect 360653 193155 360719 193158
rect 463785 193218 463851 193221
rect 463969 193218 464035 193221
rect 463785 193216 464035 193218
rect 463785 193160 463790 193216
rect 463846 193160 463974 193216
rect 464030 193160 464035 193216
rect 463785 193158 464035 193160
rect 463785 193155 463851 193158
rect 463969 193155 464035 193158
rect 470409 193218 470475 193221
rect 470593 193218 470659 193221
rect 470409 193216 470659 193218
rect 470409 193160 470414 193216
rect 470470 193160 470598 193216
rect 470654 193160 470659 193216
rect 470409 193158 470659 193160
rect 470409 193155 470475 193158
rect 470593 193155 470659 193158
rect 358445 191858 358511 191861
rect 358629 191858 358695 191861
rect 358445 191856 358695 191858
rect 249374 191824 249380 191826
rect 249198 191764 249380 191824
rect 249198 191589 249258 191764
rect 249374 191762 249380 191764
rect 249444 191762 249450 191826
rect 358445 191800 358450 191856
rect 358506 191800 358634 191856
rect 358690 191800 358695 191856
rect 358445 191798 358695 191800
rect 358445 191795 358511 191798
rect 358629 191795 358695 191798
rect 421189 191858 421255 191861
rect 421373 191858 421439 191861
rect 421189 191856 421439 191858
rect 421189 191800 421194 191856
rect 421250 191800 421378 191856
rect 421434 191800 421439 191856
rect 421189 191798 421439 191800
rect 421189 191795 421255 191798
rect 421373 191795 421439 191798
rect 249198 191584 249307 191589
rect 249198 191528 249246 191584
rect 249302 191528 249307 191584
rect 249198 191526 249307 191528
rect 249241 191523 249307 191526
rect 251449 183562 251515 183565
rect 251633 183562 251699 183565
rect 272149 183562 272215 183565
rect 251449 183560 251699 183562
rect 251449 183504 251454 183560
rect 251510 183504 251638 183560
rect 251694 183504 251699 183560
rect 251449 183502 251699 183504
rect 251449 183499 251515 183502
rect 251633 183499 251699 183502
rect 272014 183560 272215 183562
rect 272014 183504 272154 183560
rect 272210 183504 272215 183560
rect 272014 183502 272215 183504
rect 272014 183426 272074 183502
rect 272149 183499 272215 183502
rect 324589 183562 324655 183565
rect 324773 183562 324839 183565
rect 324589 183560 324839 183562
rect 324589 183504 324594 183560
rect 324650 183504 324778 183560
rect 324834 183504 324839 183560
rect 324589 183502 324839 183504
rect 324589 183499 324655 183502
rect 324773 183499 324839 183502
rect 336733 183562 336799 183565
rect 336917 183562 336983 183565
rect 336733 183560 336983 183562
rect 336733 183504 336738 183560
rect 336794 183504 336922 183560
rect 336978 183504 336983 183560
rect 336733 183502 336983 183504
rect 336733 183499 336799 183502
rect 336917 183499 336983 183502
rect 376937 183562 377003 183565
rect 377121 183562 377187 183565
rect 376937 183560 377187 183562
rect 376937 183504 376942 183560
rect 376998 183504 377126 183560
rect 377182 183504 377187 183560
rect 376937 183502 377187 183504
rect 376937 183499 377003 183502
rect 377121 183499 377187 183502
rect 386597 183562 386663 183565
rect 386965 183562 387031 183565
rect 386597 183560 387031 183562
rect 386597 183504 386602 183560
rect 386658 183504 386970 183560
rect 387026 183504 387031 183560
rect 386597 183502 387031 183504
rect 386597 183499 386663 183502
rect 386965 183499 387031 183502
rect 272333 183426 272399 183429
rect 272014 183424 272399 183426
rect 272014 183368 272338 183424
rect 272394 183368 272399 183424
rect 272014 183366 272399 183368
rect 272333 183363 272399 183366
rect 249241 182204 249307 182205
rect 249190 182202 249196 182204
rect 249150 182142 249196 182202
rect 249260 182200 249307 182204
rect 249302 182144 249307 182200
rect 249190 182140 249196 182142
rect 249260 182140 249307 182144
rect 249241 182139 249307 182140
rect 264973 182202 265039 182205
rect 265249 182202 265315 182205
rect 264973 182200 265315 182202
rect 264973 182144 264978 182200
rect 265034 182144 265254 182200
rect 265310 182144 265315 182200
rect 264973 182142 265315 182144
rect 264973 182139 265039 182142
rect 265249 182139 265315 182142
rect 267733 182202 267799 182205
rect 267917 182202 267983 182205
rect 267733 182200 267983 182202
rect 267733 182144 267738 182200
rect 267794 182144 267922 182200
rect 267978 182144 267983 182200
rect 267733 182142 267983 182144
rect 267733 182139 267799 182142
rect 267917 182139 267983 182142
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect 270769 180842 270835 180845
rect 271045 180842 271111 180845
rect 270769 180840 271111 180842
rect 270769 180784 270774 180840
rect 270830 180784 271050 180840
rect 271106 180784 271111 180840
rect 270769 180782 271111 180784
rect 270769 180779 270835 180782
rect 271045 180779 271111 180782
rect 249190 180644 249196 180708
rect 249260 180644 249266 180708
rect 249198 180570 249258 180644
rect 249425 180570 249491 180573
rect 249198 180568 249491 180570
rect 249198 180512 249430 180568
rect 249486 180512 249491 180568
rect 249198 180510 249491 180512
rect 249425 180507 249491 180510
rect -960 179482 480 179572
rect 3601 179482 3667 179485
rect -960 179480 3667 179482
rect -960 179424 3606 179480
rect 3662 179424 3667 179480
rect -960 179422 3667 179424
rect -960 179332 480 179422
rect 3601 179419 3667 179422
rect 249425 173906 249491 173909
rect 249742 173906 249748 173908
rect 249425 173904 249748 173906
rect 249425 173848 249430 173904
rect 249486 173848 249748 173904
rect 249425 173846 249748 173848
rect 249425 173843 249491 173846
rect 249742 173844 249748 173846
rect 249812 173844 249818 173908
rect 266629 173906 266695 173909
rect 266813 173906 266879 173909
rect 266629 173904 266879 173906
rect 266629 173848 266634 173904
rect 266690 173848 266818 173904
rect 266874 173848 266879 173904
rect 266629 173846 266879 173848
rect 266629 173843 266695 173846
rect 266813 173843 266879 173846
rect 372797 173906 372863 173909
rect 372981 173906 373047 173909
rect 372797 173904 373047 173906
rect 372797 173848 372802 173904
rect 372858 173848 372986 173904
rect 373042 173848 373047 173904
rect 372797 173846 373047 173848
rect 372797 173843 372863 173846
rect 372981 173843 373047 173846
rect 470409 173906 470475 173909
rect 470593 173906 470659 173909
rect 470409 173904 470659 173906
rect 470409 173848 470414 173904
rect 470470 173848 470598 173904
rect 470654 173848 470659 173904
rect 470409 173846 470659 173848
rect 470409 173843 470475 173846
rect 470593 173843 470659 173846
rect 285949 172682 286015 172685
rect 285949 172680 286058 172682
rect 285949 172624 285954 172680
rect 286010 172624 286058 172680
rect 285949 172619 286058 172624
rect 285998 172549 286058 172619
rect 285998 172544 286107 172549
rect 285998 172488 286046 172544
rect 286102 172488 286107 172544
rect 285998 172486 286107 172488
rect 286041 172483 286107 172486
rect 358537 172546 358603 172549
rect 358721 172546 358787 172549
rect 358537 172544 358787 172546
rect 358537 172488 358542 172544
rect 358598 172488 358726 172544
rect 358782 172488 358787 172544
rect 358537 172486 358787 172488
rect 358537 172483 358603 172486
rect 358721 172483 358787 172486
rect 421189 172546 421255 172549
rect 421373 172546 421439 172549
rect 421189 172544 421439 172546
rect 421189 172488 421194 172544
rect 421250 172488 421378 172544
rect 421434 172488 421439 172544
rect 421189 172486 421439 172488
rect 421189 172483 421255 172486
rect 421373 172483 421439 172486
rect 580533 170098 580599 170101
rect 583520 170098 584960 170188
rect 580533 170096 584960 170098
rect 580533 170040 580538 170096
rect 580594 170040 584960 170096
rect 580533 170038 584960 170040
rect 580533 170035 580599 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 249374 164188 249380 164252
rect 249444 164250 249450 164252
rect 249742 164250 249748 164252
rect 249444 164190 249748 164250
rect 249444 164188 249450 164190
rect 249742 164188 249748 164190
rect 249812 164188 249818 164252
rect 259637 164250 259703 164253
rect 259913 164250 259979 164253
rect 259637 164248 259979 164250
rect 259637 164192 259642 164248
rect 259698 164192 259918 164248
rect 259974 164192 259979 164248
rect 259637 164190 259979 164192
rect 259637 164187 259703 164190
rect 259913 164187 259979 164190
rect 291469 164250 291535 164253
rect 291653 164250 291719 164253
rect 291469 164248 291719 164250
rect 291469 164192 291474 164248
rect 291530 164192 291658 164248
rect 291714 164192 291719 164248
rect 291469 164190 291719 164192
rect 291469 164187 291535 164190
rect 291653 164187 291719 164190
rect 372797 164250 372863 164253
rect 372981 164250 373047 164253
rect 372797 164248 373047 164250
rect 372797 164192 372802 164248
rect 372858 164192 372986 164248
rect 373042 164192 373047 164248
rect 372797 164190 373047 164192
rect 372797 164187 372863 164190
rect 372981 164187 373047 164190
rect 470409 164250 470475 164253
rect 470593 164250 470659 164253
rect 470409 164248 470659 164250
rect 470409 164192 470414 164248
rect 470470 164192 470598 164248
rect 470654 164192 470659 164248
rect 470409 164190 470659 164192
rect 470409 164187 470475 164190
rect 470593 164187 470659 164190
rect 337193 162890 337259 162893
rect 337377 162890 337443 162893
rect 337193 162888 337443 162890
rect 337193 162832 337198 162888
rect 337254 162832 337382 162888
rect 337438 162832 337443 162888
rect 337193 162830 337443 162832
rect 337193 162827 337259 162830
rect 337377 162827 337443 162830
rect 360193 162890 360259 162893
rect 360561 162890 360627 162893
rect 360193 162888 360627 162890
rect 360193 162832 360198 162888
rect 360254 162832 360566 162888
rect 360622 162832 360627 162888
rect 360193 162830 360627 162832
rect 360193 162827 360259 162830
rect 360561 162827 360627 162830
rect 583520 158402 584960 158492
rect 583342 158342 584960 158402
rect 276054 157932 276060 157996
rect 276124 157994 276130 157996
rect 285489 157994 285555 157997
rect 276124 157992 285555 157994
rect 276124 157936 285494 157992
rect 285550 157936 285555 157992
rect 276124 157934 285555 157936
rect 276124 157932 276130 157934
rect 285489 157931 285555 157934
rect 386413 157994 386479 157997
rect 395838 157994 395844 157996
rect 386413 157992 395844 157994
rect 386413 157936 386418 157992
rect 386474 157936 395844 157992
rect 386413 157934 395844 157936
rect 386413 157931 386479 157934
rect 395838 157932 395844 157934
rect 395908 157932 395914 157996
rect 276054 157722 276060 157724
rect 269254 157662 276060 157722
rect 269254 157586 269314 157662
rect 276054 157660 276060 157662
rect 276124 157660 276130 157724
rect 333881 157722 333947 157725
rect 386413 157722 386479 157725
rect 333881 157720 334082 157722
rect 333881 157664 333886 157720
rect 333942 157664 334082 157720
rect 333881 157662 334082 157664
rect 333881 157659 333947 157662
rect 253614 157526 254410 157586
rect 249374 157388 249380 157452
rect 249444 157450 249450 157452
rect 253614 157450 253674 157526
rect 249444 157390 253674 157450
rect 254350 157450 254410 157526
rect 256190 157526 264346 157586
rect 256190 157450 256250 157526
rect 254350 157390 256250 157450
rect 264286 157450 264346 157526
rect 269070 157526 269314 157586
rect 269070 157450 269130 157526
rect 264286 157390 269130 157450
rect 285489 157450 285555 157453
rect 314694 157450 314700 157452
rect 285489 157448 305010 157450
rect 285489 157392 285494 157448
rect 285550 157392 305010 157448
rect 285489 157390 305010 157392
rect 249444 157388 249450 157390
rect 285489 157387 285555 157390
rect 304950 157178 305010 157390
rect 308998 157390 314700 157450
rect 308998 157178 309058 157390
rect 314694 157388 314700 157390
rect 314764 157388 314770 157452
rect 324221 157450 324287 157453
rect 333881 157450 333947 157453
rect 324221 157448 333947 157450
rect 324221 157392 324226 157448
rect 324282 157392 333886 157448
rect 333942 157392 333947 157448
rect 324221 157390 333947 157392
rect 334022 157450 334082 157662
rect 346350 157662 360946 157722
rect 346350 157450 346410 157662
rect 360886 157586 360946 157662
rect 375238 157720 386479 157722
rect 375238 157664 386418 157720
rect 386474 157664 386479 157720
rect 375238 157662 386479 157664
rect 364333 157586 364399 157589
rect 360886 157584 364399 157586
rect 360886 157528 364338 157584
rect 364394 157528 364399 157584
rect 360886 157526 364399 157528
rect 364333 157523 364399 157526
rect 373809 157586 373875 157589
rect 375238 157586 375298 157662
rect 386413 157659 386479 157662
rect 470550 157662 480178 157722
rect 373809 157584 375298 157586
rect 373809 157528 373814 157584
rect 373870 157528 375298 157584
rect 373809 157526 375298 157528
rect 373809 157523 373875 157526
rect 395838 157524 395844 157588
rect 395908 157586 395914 157588
rect 396073 157586 396139 157589
rect 395908 157584 396139 157586
rect 395908 157528 396078 157584
rect 396134 157528 396139 157584
rect 395908 157526 396139 157528
rect 395908 157524 395914 157526
rect 396073 157523 396139 157526
rect 400765 157586 400831 157589
rect 417877 157586 417943 157589
rect 400765 157584 405658 157586
rect 400765 157528 400770 157584
rect 400826 157528 405658 157584
rect 400765 157526 405658 157528
rect 400765 157523 400831 157526
rect 334022 157390 346410 157450
rect 405598 157450 405658 157526
rect 408542 157584 417943 157586
rect 408542 157528 417882 157584
rect 417938 157528 417943 157584
rect 408542 157526 417943 157528
rect 408542 157450 408602 157526
rect 417877 157523 417943 157526
rect 418153 157586 418219 157589
rect 437197 157586 437263 157589
rect 418153 157584 424978 157586
rect 418153 157528 418158 157584
rect 418214 157528 424978 157584
rect 418153 157526 424978 157528
rect 418153 157523 418219 157526
rect 405598 157390 408602 157450
rect 424918 157450 424978 157526
rect 427862 157584 437263 157586
rect 427862 157528 437202 157584
rect 437258 157528 437263 157584
rect 427862 157526 437263 157528
rect 427862 157450 427922 157526
rect 437197 157523 437263 157526
rect 437473 157586 437539 157589
rect 456517 157586 456583 157589
rect 437473 157584 444298 157586
rect 437473 157528 437478 157584
rect 437534 157528 444298 157584
rect 437473 157526 444298 157528
rect 437473 157523 437539 157526
rect 424918 157390 427922 157450
rect 444238 157450 444298 157526
rect 447182 157584 456583 157586
rect 447182 157528 456522 157584
rect 456578 157528 456583 157584
rect 447182 157526 456583 157528
rect 447182 157450 447242 157526
rect 456517 157523 456583 157526
rect 458265 157586 458331 157589
rect 458265 157584 463618 157586
rect 458265 157528 458270 157584
rect 458326 157528 463618 157584
rect 458265 157526 463618 157528
rect 458265 157523 458331 157526
rect 444238 157390 447242 157450
rect 463558 157450 463618 157526
rect 470550 157450 470610 157662
rect 463558 157390 470610 157450
rect 480118 157450 480178 157662
rect 480302 157662 489930 157722
rect 480302 157450 480362 157662
rect 489870 157586 489930 157662
rect 499622 157662 509250 157722
rect 489870 157526 499498 157586
rect 480118 157390 480362 157450
rect 499438 157450 499498 157526
rect 499622 157450 499682 157662
rect 509190 157586 509250 157662
rect 518942 157662 528570 157722
rect 509190 157526 518818 157586
rect 499438 157390 499682 157450
rect 518758 157450 518818 157526
rect 518942 157450 519002 157662
rect 528510 157586 528570 157662
rect 538262 157662 547890 157722
rect 528510 157526 538138 157586
rect 518758 157390 519002 157450
rect 538078 157450 538138 157526
rect 538262 157450 538322 157662
rect 547830 157586 547890 157662
rect 557582 157662 567210 157722
rect 547830 157526 557458 157586
rect 538078 157390 538322 157450
rect 557398 157450 557458 157526
rect 557582 157450 557642 157662
rect 567150 157586 567210 157662
rect 583342 157586 583402 158342
rect 583520 158252 584960 158342
rect 567150 157526 576778 157586
rect 557398 157390 557642 157450
rect 576718 157450 576778 157526
rect 576902 157526 583402 157586
rect 576902 157450 576962 157526
rect 576718 157390 576962 157450
rect 324221 157387 324287 157390
rect 333881 157387 333947 157390
rect 304950 157118 309058 157178
rect 314694 157116 314700 157180
rect 314764 157178 314770 157180
rect 324221 157178 324287 157181
rect 314764 157176 324287 157178
rect 314764 157120 324226 157176
rect 324282 157120 324287 157176
rect 314764 157118 324287 157120
rect 314764 157116 314770 157118
rect 324221 157115 324287 157118
rect 250345 154730 250411 154733
rect 249934 154728 250411 154730
rect 249934 154672 250350 154728
rect 250406 154672 250411 154728
rect 249934 154670 250411 154672
rect 236269 154594 236335 154597
rect 236453 154594 236519 154597
rect 236269 154592 236519 154594
rect 236269 154536 236274 154592
rect 236330 154536 236458 154592
rect 236514 154536 236519 154592
rect 236269 154534 236519 154536
rect 236269 154531 236335 154534
rect 236453 154531 236519 154534
rect 244273 154594 244339 154597
rect 244457 154594 244523 154597
rect 244273 154592 244523 154594
rect 244273 154536 244278 154592
rect 244334 154536 244462 154592
rect 244518 154536 244523 154592
rect 244273 154534 244523 154536
rect 249934 154594 249994 154670
rect 250345 154667 250411 154670
rect 250069 154594 250135 154597
rect 249934 154592 250135 154594
rect 249934 154536 250074 154592
rect 250130 154536 250135 154592
rect 249934 154534 250135 154536
rect 244273 154531 244339 154534
rect 244457 154531 244523 154534
rect 250069 154531 250135 154534
rect 251449 154594 251515 154597
rect 251633 154594 251699 154597
rect 251449 154592 251699 154594
rect 251449 154536 251454 154592
rect 251510 154536 251638 154592
rect 251694 154536 251699 154592
rect 251449 154534 251699 154536
rect 251449 154531 251515 154534
rect 251633 154531 251699 154534
rect 386505 154594 386571 154597
rect 386781 154594 386847 154597
rect 386505 154592 386847 154594
rect 386505 154536 386510 154592
rect 386566 154536 386786 154592
rect 386842 154536 386847 154592
rect 386505 154534 386847 154536
rect 386505 154531 386571 154534
rect 386781 154531 386847 154534
rect 310881 153370 310947 153373
rect 310838 153368 310947 153370
rect 310838 153312 310886 153368
rect 310942 153312 310947 153368
rect 310838 153307 310947 153312
rect 310838 153237 310898 153307
rect 232129 153234 232195 153237
rect 232313 153234 232379 153237
rect 232129 153232 232379 153234
rect 232129 153176 232134 153232
rect 232190 153176 232318 153232
rect 232374 153176 232379 153232
rect 232129 153174 232379 153176
rect 232129 153171 232195 153174
rect 232313 153171 232379 153174
rect 310789 153232 310898 153237
rect 310789 153176 310794 153232
rect 310850 153176 310898 153232
rect 310789 153174 310898 153176
rect 358537 153234 358603 153237
rect 358721 153234 358787 153237
rect 358537 153232 358787 153234
rect 358537 153176 358542 153232
rect 358598 153176 358726 153232
rect 358782 153176 358787 153232
rect 358537 153174 358787 153176
rect 310789 153171 310855 153174
rect 358537 153171 358603 153174
rect 358721 153171 358787 153174
rect 360193 153234 360259 153237
rect 360377 153234 360443 153237
rect 360193 153232 360443 153234
rect 360193 153176 360198 153232
rect 360254 153176 360382 153232
rect 360438 153176 360443 153232
rect 360193 153174 360443 153176
rect 360193 153171 360259 153174
rect 360377 153171 360443 153174
rect -960 150786 480 150876
rect 3325 150786 3391 150789
rect -960 150784 3391 150786
rect -960 150728 3330 150784
rect 3386 150728 3391 150784
rect -960 150726 3391 150728
rect -960 150636 480 150726
rect 3325 150723 3391 150726
rect 583520 146556 584960 146796
rect 327257 145074 327323 145077
rect 327214 145072 327323 145074
rect 327214 145016 327262 145072
rect 327318 145016 327323 145072
rect 327214 145011 327323 145016
rect 327214 144941 327274 145011
rect 247125 144938 247191 144941
rect 247309 144938 247375 144941
rect 247125 144936 247375 144938
rect 247125 144880 247130 144936
rect 247186 144880 247314 144936
rect 247370 144880 247375 144936
rect 247125 144878 247375 144880
rect 247125 144875 247191 144878
rect 247309 144875 247375 144878
rect 301037 144938 301103 144941
rect 301221 144938 301287 144941
rect 324589 144938 324655 144941
rect 301037 144936 301287 144938
rect 301037 144880 301042 144936
rect 301098 144880 301226 144936
rect 301282 144880 301287 144936
rect 301037 144878 301287 144880
rect 301037 144875 301103 144878
rect 301221 144875 301287 144878
rect 324454 144936 324655 144938
rect 324454 144880 324594 144936
rect 324650 144880 324655 144936
rect 324454 144878 324655 144880
rect 324454 144802 324514 144878
rect 324589 144875 324655 144878
rect 325877 144938 325943 144941
rect 326061 144938 326127 144941
rect 325877 144936 326127 144938
rect 325877 144880 325882 144936
rect 325938 144880 326066 144936
rect 326122 144880 326127 144936
rect 325877 144878 326127 144880
rect 325877 144875 325943 144878
rect 326061 144875 326127 144878
rect 327165 144936 327274 144941
rect 327165 144880 327170 144936
rect 327226 144880 327274 144936
rect 327165 144878 327274 144880
rect 339493 144938 339559 144941
rect 339677 144938 339743 144941
rect 339493 144936 339743 144938
rect 339493 144880 339498 144936
rect 339554 144880 339682 144936
rect 339738 144880 339743 144936
rect 339493 144878 339743 144880
rect 327165 144875 327231 144878
rect 339493 144875 339559 144878
rect 339677 144875 339743 144878
rect 470409 144938 470475 144941
rect 470593 144938 470659 144941
rect 470409 144936 470659 144938
rect 470409 144880 470414 144936
rect 470470 144880 470598 144936
rect 470654 144880 470659 144936
rect 470409 144878 470659 144880
rect 470409 144875 470475 144878
rect 470593 144875 470659 144878
rect 324589 144802 324655 144805
rect 324454 144800 324655 144802
rect 324454 144744 324594 144800
rect 324650 144744 324655 144800
rect 324454 144742 324655 144744
rect 324589 144739 324655 144742
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 250253 135418 250319 135421
rect 266721 135418 266787 135421
rect 249934 135416 250319 135418
rect 249934 135360 250258 135416
rect 250314 135360 250319 135416
rect 249934 135358 250319 135360
rect 236269 135282 236335 135285
rect 236453 135282 236519 135285
rect 236269 135280 236519 135282
rect 236269 135224 236274 135280
rect 236330 135224 236458 135280
rect 236514 135224 236519 135280
rect 236269 135222 236519 135224
rect 236269 135219 236335 135222
rect 236453 135219 236519 135222
rect 239029 135282 239095 135285
rect 239213 135282 239279 135285
rect 239029 135280 239279 135282
rect 239029 135224 239034 135280
rect 239090 135224 239218 135280
rect 239274 135224 239279 135280
rect 239029 135222 239279 135224
rect 239029 135219 239095 135222
rect 239213 135219 239279 135222
rect 244273 135282 244339 135285
rect 244457 135282 244523 135285
rect 244273 135280 244523 135282
rect 244273 135224 244278 135280
rect 244334 135224 244462 135280
rect 244518 135224 244523 135280
rect 244273 135222 244523 135224
rect 249934 135282 249994 135358
rect 250253 135355 250319 135358
rect 266678 135416 266787 135418
rect 266678 135360 266726 135416
rect 266782 135360 266787 135416
rect 266678 135355 266787 135360
rect 266678 135285 266738 135355
rect 250069 135282 250135 135285
rect 249934 135280 250135 135282
rect 249934 135224 250074 135280
rect 250130 135224 250135 135280
rect 249934 135222 250135 135224
rect 244273 135219 244339 135222
rect 244457 135219 244523 135222
rect 250069 135219 250135 135222
rect 266629 135280 266738 135285
rect 266629 135224 266634 135280
rect 266690 135224 266738 135280
rect 266629 135222 266738 135224
rect 386413 135282 386479 135285
rect 386689 135282 386755 135285
rect 386413 135280 386755 135282
rect 386413 135224 386418 135280
rect 386474 135224 386694 135280
rect 386750 135224 386755 135280
rect 386413 135222 386755 135224
rect 266629 135219 266695 135222
rect 386413 135219 386479 135222
rect 386689 135219 386755 135222
rect 580441 134874 580507 134877
rect 583520 134874 584960 134964
rect 580441 134872 584960 134874
rect 580441 134816 580446 134872
rect 580502 134816 584960 134872
rect 580441 134814 584960 134816
rect 580441 134811 580507 134814
rect 583520 134724 584960 134814
rect 357433 125762 357499 125765
rect 357390 125760 357499 125762
rect 357390 125704 357438 125760
rect 357494 125704 357499 125760
rect 357390 125699 357499 125704
rect 262581 125626 262647 125629
rect 262765 125626 262831 125629
rect 262581 125624 262831 125626
rect 262581 125568 262586 125624
rect 262642 125568 262770 125624
rect 262826 125568 262831 125624
rect 262581 125566 262831 125568
rect 262581 125563 262647 125566
rect 262765 125563 262831 125566
rect 267733 125626 267799 125629
rect 267917 125626 267983 125629
rect 267733 125624 267983 125626
rect 267733 125568 267738 125624
rect 267794 125568 267922 125624
rect 267978 125568 267983 125624
rect 267733 125566 267983 125568
rect 267733 125563 267799 125566
rect 267917 125563 267983 125566
rect 270493 125626 270559 125629
rect 270677 125626 270743 125629
rect 270493 125624 270743 125626
rect 270493 125568 270498 125624
rect 270554 125568 270682 125624
rect 270738 125568 270743 125624
rect 270493 125566 270743 125568
rect 357390 125626 357450 125699
rect 357525 125626 357591 125629
rect 357390 125624 357591 125626
rect 357390 125568 357530 125624
rect 357586 125568 357591 125624
rect 357390 125566 357591 125568
rect 270493 125563 270559 125566
rect 270677 125563 270743 125566
rect 357525 125563 357591 125566
rect 470409 125626 470475 125629
rect 470593 125626 470659 125629
rect 470409 125624 470659 125626
rect 470409 125568 470414 125624
rect 470470 125568 470598 125624
rect 470654 125568 470659 125624
rect 470409 125566 470659 125568
rect 470409 125563 470475 125566
rect 470593 125563 470659 125566
rect 306833 124266 306899 124269
rect 307017 124266 307083 124269
rect 306833 124264 307083 124266
rect 306833 124208 306838 124264
rect 306894 124208 307022 124264
rect 307078 124208 307083 124264
rect 306833 124206 307083 124208
rect 306833 124203 306899 124206
rect 307017 124203 307083 124206
rect 580349 123178 580415 123181
rect 583520 123178 584960 123268
rect 580349 123176 584960 123178
rect 580349 123120 580354 123176
rect 580410 123120 584960 123176
rect 580349 123118 584960 123120
rect 580349 123115 580415 123118
rect 583520 123028 584960 123118
rect 285949 122770 286015 122773
rect 286225 122770 286291 122773
rect 285949 122768 286291 122770
rect 285949 122712 285954 122768
rect 286010 122712 286230 122768
rect 286286 122712 286291 122768
rect 285949 122710 286291 122712
rect 285949 122707 286015 122710
rect 286225 122707 286291 122710
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 266721 116106 266787 116109
rect 310973 116106 311039 116109
rect 323393 116106 323459 116109
rect 266678 116104 266787 116106
rect 266678 116048 266726 116104
rect 266782 116048 266787 116104
rect 266678 116043 266787 116048
rect 310838 116104 311039 116106
rect 310838 116048 310978 116104
rect 311034 116048 311039 116104
rect 310838 116046 311039 116048
rect 266678 115973 266738 116043
rect 310838 115973 310898 116046
rect 310973 116043 311039 116046
rect 323350 116104 323459 116106
rect 323350 116048 323398 116104
rect 323454 116048 323459 116104
rect 323350 116043 323459 116048
rect 323350 115973 323410 116043
rect 236269 115970 236335 115973
rect 236453 115970 236519 115973
rect 236269 115968 236519 115970
rect 236269 115912 236274 115968
rect 236330 115912 236458 115968
rect 236514 115912 236519 115968
rect 236269 115910 236519 115912
rect 236269 115907 236335 115910
rect 236453 115907 236519 115910
rect 266629 115968 266738 115973
rect 266629 115912 266634 115968
rect 266690 115912 266738 115968
rect 266629 115910 266738 115912
rect 310789 115968 310898 115973
rect 310789 115912 310794 115968
rect 310850 115912 310898 115968
rect 310789 115910 310898 115912
rect 317781 115970 317847 115973
rect 317965 115970 318031 115973
rect 317781 115968 318031 115970
rect 317781 115912 317786 115968
rect 317842 115912 317970 115968
rect 318026 115912 318031 115968
rect 317781 115910 318031 115912
rect 266629 115907 266695 115910
rect 310789 115907 310855 115910
rect 317781 115907 317847 115910
rect 317965 115907 318031 115910
rect 323301 115968 323410 115973
rect 323301 115912 323306 115968
rect 323362 115912 323410 115968
rect 323301 115910 323410 115912
rect 336733 115970 336799 115973
rect 336917 115970 336983 115973
rect 336733 115968 336983 115970
rect 336733 115912 336738 115968
rect 336794 115912 336922 115968
rect 336978 115912 336983 115968
rect 336733 115910 336983 115912
rect 323301 115907 323367 115910
rect 336733 115907 336799 115910
rect 336917 115907 336983 115910
rect 386413 115970 386479 115973
rect 386597 115970 386663 115973
rect 386413 115968 386663 115970
rect 386413 115912 386418 115968
rect 386474 115912 386602 115968
rect 386658 115912 386663 115968
rect 386413 115910 386663 115912
rect 386413 115907 386479 115910
rect 386597 115907 386663 115910
rect 580257 111482 580323 111485
rect 583520 111482 584960 111572
rect 580257 111480 584960 111482
rect 580257 111424 580262 111480
rect 580318 111424 584960 111480
rect 580257 111422 584960 111424
rect 580257 111419 580323 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 360469 106450 360535 106453
rect 360334 106448 360535 106450
rect 360334 106392 360474 106448
rect 360530 106392 360535 106448
rect 360334 106390 360535 106392
rect 360334 106317 360394 106390
rect 360469 106387 360535 106390
rect 376937 106450 377003 106453
rect 377121 106450 377187 106453
rect 376937 106448 377187 106450
rect 376937 106392 376942 106448
rect 376998 106392 377126 106448
rect 377182 106392 377187 106448
rect 376937 106390 377187 106392
rect 376937 106387 377003 106390
rect 377121 106387 377187 106390
rect 270677 106314 270743 106317
rect 270861 106314 270927 106317
rect 270677 106312 270927 106314
rect 270677 106256 270682 106312
rect 270738 106256 270866 106312
rect 270922 106256 270927 106312
rect 270677 106254 270927 106256
rect 360334 106312 360443 106317
rect 360334 106256 360382 106312
rect 360438 106256 360443 106312
rect 360334 106254 360443 106256
rect 270677 106251 270743 106254
rect 270861 106251 270927 106254
rect 360377 106251 360443 106254
rect 375557 106314 375623 106317
rect 375741 106314 375807 106317
rect 375557 106312 375807 106314
rect 375557 106256 375562 106312
rect 375618 106256 375746 106312
rect 375802 106256 375807 106312
rect 375557 106254 375807 106256
rect 375557 106251 375623 106254
rect 375741 106251 375807 106254
rect 463877 106314 463943 106317
rect 464061 106314 464127 106317
rect 463877 106312 464127 106314
rect 463877 106256 463882 106312
rect 463938 106256 464066 106312
rect 464122 106256 464127 106312
rect 463877 106254 464127 106256
rect 463877 106251 463943 106254
rect 464061 106251 464127 106254
rect 306833 103594 306899 103597
rect 307017 103594 307083 103597
rect 306833 103592 307083 103594
rect 306833 103536 306838 103592
rect 306894 103536 307022 103592
rect 307078 103536 307083 103592
rect 306833 103534 307083 103536
rect 306833 103531 306899 103534
rect 307017 103531 307083 103534
rect 329925 103594 329991 103597
rect 330109 103594 330175 103597
rect 329925 103592 330175 103594
rect 329925 103536 329930 103592
rect 329986 103536 330114 103592
rect 330170 103536 330175 103592
rect 329925 103534 330175 103536
rect 329925 103531 329991 103534
rect 330109 103531 330175 103534
rect 583520 99636 584960 99876
rect 236269 96658 236335 96661
rect 236637 96658 236703 96661
rect 236269 96656 236703 96658
rect 236269 96600 236274 96656
rect 236330 96600 236642 96656
rect 236698 96600 236703 96656
rect 236269 96598 236703 96600
rect 236269 96595 236335 96598
rect 236637 96595 236703 96598
rect 239121 96658 239187 96661
rect 239305 96658 239371 96661
rect 239121 96656 239371 96658
rect 239121 96600 239126 96656
rect 239182 96600 239310 96656
rect 239366 96600 239371 96656
rect 239121 96598 239371 96600
rect 239121 96595 239187 96598
rect 239305 96595 239371 96598
rect 360285 96658 360351 96661
rect 360561 96658 360627 96661
rect 360285 96656 360627 96658
rect 360285 96600 360290 96656
rect 360346 96600 360566 96656
rect 360622 96600 360627 96656
rect 360285 96598 360627 96600
rect 360285 96595 360351 96598
rect 360561 96595 360627 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 285622 87484 285628 87548
rect 285692 87546 285698 87548
rect 295241 87546 295307 87549
rect 285692 87544 295307 87546
rect 285692 87488 295246 87544
rect 295302 87488 295307 87544
rect 285692 87486 295307 87488
rect 285692 87484 285698 87486
rect 295241 87483 295307 87486
rect 466085 87546 466151 87549
rect 466085 87544 473370 87546
rect 466085 87488 466090 87544
rect 466146 87488 473370 87544
rect 466085 87486 473370 87488
rect 466085 87483 466151 87486
rect 315941 87410 316007 87413
rect 473310 87410 473370 87486
rect 315941 87408 317338 87410
rect 315941 87352 315946 87408
rect 316002 87352 317338 87408
rect 315941 87350 317338 87352
rect 315941 87347 316007 87350
rect 251214 87274 251220 87276
rect 246254 87214 251220 87274
rect 239990 87076 239996 87140
rect 240060 87138 240066 87140
rect 246254 87138 246314 87214
rect 251214 87212 251220 87214
rect 251284 87212 251290 87276
rect 285622 87274 285628 87276
rect 265022 87214 285628 87274
rect 240060 87104 244106 87138
rect 244230 87104 246314 87138
rect 240060 87078 246314 87104
rect 251173 87140 251239 87141
rect 251173 87136 251220 87140
rect 251284 87138 251290 87140
rect 260649 87138 260715 87141
rect 265022 87138 265082 87214
rect 285622 87212 285628 87214
rect 285692 87212 285698 87276
rect 317278 87274 317338 87350
rect 396030 87350 405658 87410
rect 473310 87350 476314 87410
rect 328453 87274 328519 87277
rect 357341 87274 357407 87277
rect 317278 87214 325802 87274
rect 251173 87080 251178 87136
rect 240060 87076 240066 87078
rect 244046 87044 244290 87078
rect 251173 87076 251220 87080
rect 251284 87078 251330 87138
rect 260649 87136 265082 87138
rect 260649 87080 260654 87136
rect 260710 87080 265082 87136
rect 260649 87078 265082 87080
rect 296621 87138 296687 87141
rect 315941 87138 316007 87141
rect 296621 87136 298018 87138
rect 296621 87080 296626 87136
rect 296682 87080 298018 87136
rect 296621 87078 298018 87080
rect 251284 87076 251290 87078
rect 251173 87075 251239 87076
rect 260649 87075 260715 87078
rect 296621 87075 296687 87078
rect 295241 87002 295307 87005
rect 296621 87002 296687 87005
rect 295241 87000 296687 87002
rect 295241 86944 295246 87000
rect 295302 86944 296626 87000
rect 296682 86944 296687 87000
rect 295241 86942 296687 86944
rect 295241 86939 295307 86942
rect 296621 86939 296687 86942
rect 297958 86866 298018 87078
rect 308814 87136 316007 87138
rect 308814 87080 315946 87136
rect 316002 87080 316007 87136
rect 308814 87078 316007 87080
rect 325742 87138 325802 87214
rect 328453 87272 340890 87274
rect 328453 87216 328458 87272
rect 328514 87216 340890 87272
rect 328453 87214 340890 87216
rect 328453 87211 328519 87214
rect 328361 87138 328427 87141
rect 325742 87136 328427 87138
rect 325742 87080 328366 87136
rect 328422 87080 328427 87136
rect 325742 87078 328427 87080
rect 308814 87002 308874 87078
rect 315941 87075 316007 87078
rect 328361 87075 328427 87078
rect 298142 86942 308874 87002
rect 340830 87002 340890 87214
rect 357341 87272 360210 87274
rect 357341 87216 357346 87272
rect 357402 87216 360210 87272
rect 357341 87214 360210 87216
rect 357341 87211 357407 87214
rect 347773 87002 347839 87005
rect 340830 87000 347839 87002
rect 340830 86944 347778 87000
rect 347834 86944 347839 87000
rect 340830 86942 347839 86944
rect 298142 86866 298202 86942
rect 347773 86939 347839 86942
rect 358721 87002 358787 87005
rect 358997 87002 359063 87005
rect 358721 87000 359063 87002
rect 358721 86944 358726 87000
rect 358782 86944 359002 87000
rect 359058 86944 359063 87000
rect 358721 86942 359063 86944
rect 360150 87002 360210 87214
rect 367142 87214 379530 87274
rect 367142 87141 367202 87214
rect 367093 87136 367202 87141
rect 367093 87080 367098 87136
rect 367154 87080 367202 87136
rect 367093 87078 367202 87080
rect 367093 87075 367159 87078
rect 367093 87002 367159 87005
rect 360150 87000 367159 87002
rect 360150 86944 367098 87000
rect 367154 86944 367159 87000
rect 360150 86942 367159 86944
rect 358721 86939 358787 86942
rect 358997 86939 359063 86942
rect 367093 86939 367159 86942
rect 375373 87002 375439 87005
rect 375649 87002 375715 87005
rect 375373 87000 375715 87002
rect 375373 86944 375378 87000
rect 375434 86944 375654 87000
rect 375710 86944 375715 87000
rect 375373 86942 375715 86944
rect 379470 87002 379530 87214
rect 396030 87138 396090 87350
rect 405598 87276 405658 87350
rect 405590 87212 405596 87276
rect 405660 87212 405666 87276
rect 454033 87274 454099 87277
rect 447182 87272 454099 87274
rect 447182 87216 454038 87272
rect 454094 87216 454099 87272
rect 447182 87214 454099 87216
rect 437197 87138 437263 87141
rect 389222 87078 396090 87138
rect 408542 87078 424978 87138
rect 389222 87002 389282 87078
rect 379470 86942 389282 87002
rect 375373 86939 375439 86942
rect 375649 86939 375715 86942
rect 405590 86940 405596 87004
rect 405660 87002 405666 87004
rect 408542 87002 408602 87078
rect 405660 86942 408602 87002
rect 424918 87002 424978 87078
rect 427862 87136 437263 87138
rect 427862 87080 437202 87136
rect 437258 87080 437263 87136
rect 427862 87078 437263 87080
rect 427862 87002 427922 87078
rect 437197 87075 437263 87078
rect 437473 87138 437539 87141
rect 437473 87136 444298 87138
rect 437473 87080 437478 87136
rect 437534 87080 444298 87136
rect 437473 87078 444298 87080
rect 437473 87075 437539 87078
rect 424918 86942 427922 87002
rect 444238 87002 444298 87078
rect 447182 87002 447242 87214
rect 454033 87211 454099 87214
rect 456977 87274 457043 87277
rect 456977 87272 463618 87274
rect 456977 87216 456982 87272
rect 457038 87216 463618 87272
rect 456977 87214 463618 87216
rect 456977 87211 457043 87214
rect 463558 87138 463618 87214
rect 466085 87138 466151 87141
rect 463558 87136 466151 87138
rect 463558 87080 466090 87136
rect 466146 87080 466151 87136
rect 463558 87078 466151 87080
rect 476254 87138 476314 87350
rect 481582 87348 481588 87412
rect 481652 87410 481658 87412
rect 491201 87410 491267 87413
rect 481652 87408 491267 87410
rect 481652 87352 491206 87408
rect 491262 87352 491267 87408
rect 481652 87350 491267 87352
rect 481652 87348 481658 87350
rect 491201 87347 491267 87350
rect 502241 87274 502307 87277
rect 502241 87272 509250 87274
rect 502241 87216 502246 87272
rect 502302 87216 509250 87272
rect 502241 87214 509250 87216
rect 502241 87211 502307 87214
rect 481582 87138 481588 87140
rect 476254 87078 481588 87138
rect 466085 87075 466151 87078
rect 481582 87076 481588 87078
rect 481652 87076 481658 87140
rect 509190 87138 509250 87214
rect 518942 87214 528570 87274
rect 509190 87078 518818 87138
rect 444238 86942 447242 87002
rect 491201 87002 491267 87005
rect 494605 87002 494671 87005
rect 491201 87000 494671 87002
rect 491201 86944 491206 87000
rect 491262 86944 494610 87000
rect 494666 86944 494671 87000
rect 491201 86942 494671 86944
rect 518758 87002 518818 87078
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 538262 87214 547890 87274
rect 528510 87078 538138 87138
rect 518758 86942 519002 87002
rect 538078 87002 538138 87078
rect 538262 87002 538322 87214
rect 547830 87138 547890 87214
rect 557582 87214 567210 87274
rect 547830 87078 557458 87138
rect 538078 86942 538322 87002
rect 557398 87002 557458 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 557398 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 405660 86940 405666 86942
rect 491201 86939 491267 86942
rect 494605 86939 494671 86942
rect 297958 86806 298202 86866
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 367001 77482 367067 77485
rect 366958 77480 367067 77482
rect 366958 77424 367006 77480
rect 367062 77424 367067 77480
rect 366958 77419 367067 77424
rect 366958 77349 367018 77419
rect 366958 77344 367067 77349
rect 366958 77288 367006 77344
rect 367062 77288 367067 77344
rect 366958 77286 367067 77288
rect 367001 77283 367067 77286
rect 386413 76530 386479 76533
rect 395838 76530 395844 76532
rect 386413 76528 395844 76530
rect 386413 76472 386418 76528
rect 386474 76472 395844 76528
rect 386413 76470 395844 76472
rect 386413 76467 386479 76470
rect 395838 76468 395844 76470
rect 395908 76468 395914 76532
rect 466085 76530 466151 76533
rect 466085 76528 473370 76530
rect 466085 76472 466090 76528
rect 466146 76472 473370 76528
rect 466085 76470 473370 76472
rect 466085 76467 466151 76470
rect 473310 76394 473370 76470
rect 482921 76394 482987 76397
rect 487797 76394 487863 76397
rect 473310 76392 482987 76394
rect 473310 76336 482926 76392
rect 482982 76336 482987 76392
rect 473310 76334 482987 76336
rect 482921 76331 482987 76334
rect 483062 76392 487863 76394
rect 483062 76336 487802 76392
rect 487858 76336 487863 76392
rect 483062 76334 487863 76336
rect 338021 76258 338087 76261
rect 376661 76258 376727 76261
rect 386413 76258 386479 76261
rect 338021 76256 340890 76258
rect 338021 76200 338026 76256
rect 338082 76200 340890 76256
rect 338021 76198 340890 76200
rect 338021 76195 338087 76198
rect 241278 76060 241284 76124
rect 241348 76122 241354 76124
rect 306281 76122 306347 76125
rect 241348 76062 254042 76122
rect 241348 76060 241354 76062
rect 253982 75986 254042 76062
rect 306281 76120 309426 76122
rect 306281 76064 306286 76120
rect 306342 76064 309426 76120
rect 306281 76062 309426 76064
rect 306281 76059 306347 76062
rect 295241 75986 295307 75989
rect 309366 75986 309426 76062
rect 328913 75986 328979 75989
rect 253982 75926 282194 75986
rect 282134 75850 282194 75926
rect 295241 75984 297834 75986
rect 295241 75928 295246 75984
rect 295302 75928 297834 75984
rect 295241 75926 297834 75928
rect 309366 75984 328979 75986
rect 309366 75928 328918 75984
rect 328974 75928 328979 75984
rect 309366 75926 328979 75928
rect 340830 75986 340890 76198
rect 376661 76256 386479 76258
rect 376661 76200 376666 76256
rect 376722 76200 386418 76256
rect 386474 76200 386479 76256
rect 376661 76198 386479 76200
rect 376661 76195 376727 76198
rect 386413 76195 386479 76198
rect 447182 76198 463618 76258
rect 369853 76122 369919 76125
rect 350582 76120 369919 76122
rect 350582 76064 369858 76120
rect 369914 76064 369919 76120
rect 350582 76062 369919 76064
rect 350582 75986 350642 76062
rect 369853 76059 369919 76062
rect 395838 76060 395844 76124
rect 395908 76122 395914 76124
rect 396073 76122 396139 76125
rect 395908 76120 396139 76122
rect 395908 76064 396078 76120
rect 396134 76064 396139 76120
rect 395908 76062 396139 76064
rect 395908 76060 395914 76062
rect 396073 76059 396139 76062
rect 399385 76122 399451 76125
rect 414013 76122 414079 76125
rect 437197 76122 437263 76125
rect 399385 76120 405658 76122
rect 399385 76064 399390 76120
rect 399446 76064 405658 76120
rect 399385 76062 405658 76064
rect 399385 76059 399451 76062
rect 340830 75926 350642 75986
rect 405598 75986 405658 76062
rect 408542 76120 414079 76122
rect 408542 76064 414018 76120
rect 414074 76064 414079 76120
rect 408542 76062 414079 76064
rect 408542 75986 408602 76062
rect 414013 76059 414079 76062
rect 427862 76120 437263 76122
rect 427862 76064 437202 76120
rect 437258 76064 437263 76120
rect 427862 76062 437263 76064
rect 405598 75926 408602 75986
rect 423489 75986 423555 75989
rect 427862 75986 427922 76062
rect 437197 76059 437263 76062
rect 437473 76122 437539 76125
rect 437473 76120 444298 76122
rect 437473 76064 437478 76120
rect 437534 76064 444298 76120
rect 437473 76062 444298 76064
rect 437473 76059 437539 76062
rect 423489 75984 427922 75986
rect 423489 75928 423494 75984
rect 423550 75928 427922 75984
rect 423489 75926 427922 75928
rect 444238 75986 444298 76062
rect 447182 75986 447242 76198
rect 463558 76122 463618 76198
rect 466085 76122 466151 76125
rect 463558 76120 466151 76122
rect 463558 76064 466090 76120
rect 466146 76064 466151 76120
rect 463558 76062 466151 76064
rect 466085 76059 466151 76062
rect 482921 76122 482987 76125
rect 483062 76122 483122 76334
rect 487797 76331 487863 76334
rect 492622 76196 492628 76260
rect 492692 76258 492698 76260
rect 583520 76258 584960 76348
rect 492692 76198 509250 76258
rect 492692 76196 492698 76198
rect 482921 76120 483122 76122
rect 482921 76064 482926 76120
rect 482982 76064 483122 76120
rect 482921 76062 483122 76064
rect 509190 76122 509250 76198
rect 518942 76198 528570 76258
rect 509190 76062 518818 76122
rect 482921 76059 482987 76062
rect 444238 75926 447242 75986
rect 487797 75986 487863 75989
rect 492622 75986 492628 75988
rect 487797 75984 492628 75986
rect 487797 75928 487802 75984
rect 487858 75928 492628 75984
rect 487797 75926 492628 75928
rect 295241 75923 295307 75926
rect 285622 75850 285628 75852
rect 282134 75790 285628 75850
rect 285622 75788 285628 75790
rect 285692 75788 285698 75852
rect 297774 75850 297834 75926
rect 328913 75923 328979 75926
rect 423489 75923 423555 75926
rect 487797 75923 487863 75926
rect 492622 75924 492628 75926
rect 492692 75924 492698 75988
rect 518758 75986 518818 76062
rect 518942 75986 519002 76198
rect 528510 76122 528570 76198
rect 538262 76198 547890 76258
rect 528510 76062 538138 76122
rect 518758 75926 519002 75986
rect 538078 75986 538138 76062
rect 538262 75986 538322 76198
rect 547830 76122 547890 76198
rect 557582 76198 567210 76258
rect 547830 76062 557458 76122
rect 538078 75926 538322 75986
rect 557398 75986 557458 76062
rect 557582 75986 557642 76198
rect 567150 76122 567210 76198
rect 583342 76198 584960 76258
rect 583342 76122 583402 76198
rect 567150 76062 576778 76122
rect 557398 75926 557642 75986
rect 576718 75986 576778 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 576718 75926 576962 75986
rect 306281 75850 306347 75853
rect 297774 75848 306347 75850
rect 297774 75792 306286 75848
rect 306342 75792 306347 75848
rect 297774 75790 306347 75792
rect 306281 75787 306347 75790
rect 285622 75516 285628 75580
rect 285692 75578 285698 75580
rect 295241 75578 295307 75581
rect 285692 75576 295307 75578
rect 285692 75520 295246 75576
rect 295302 75520 295307 75576
rect 285692 75518 295307 75520
rect 285692 75516 285698 75518
rect 295241 75515 295307 75518
rect 301221 66330 301287 66333
rect 301086 66328 301287 66330
rect 301086 66272 301226 66328
rect 301282 66272 301287 66328
rect 301086 66270 301287 66272
rect 301086 66058 301146 66270
rect 301221 66267 301287 66270
rect 301221 66058 301287 66061
rect 301086 66056 301287 66058
rect 301086 66000 301226 66056
rect 301282 66000 301287 66056
rect 301086 65998 301287 66000
rect 301221 65995 301287 65998
rect 288709 64834 288775 64837
rect 288893 64834 288959 64837
rect 288709 64832 288959 64834
rect 288709 64776 288714 64832
rect 288770 64776 288898 64832
rect 288954 64776 288959 64832
rect 288709 64774 288959 64776
rect 288709 64771 288775 64774
rect 288893 64771 288959 64774
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect 583520 64562 584960 64652
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 583342 64502 584960 64562
rect 405406 64018 405412 64020
rect 398606 63958 405412 64018
rect 327022 63820 327028 63884
rect 327092 63882 327098 63884
rect 376661 63882 376727 63885
rect 378501 63882 378567 63885
rect 327092 63822 340890 63882
rect 327092 63820 327098 63822
rect 260741 63746 260807 63749
rect 263409 63746 263475 63749
rect 260741 63744 263475 63746
rect 260741 63688 260746 63744
rect 260802 63688 263414 63744
rect 263470 63688 263475 63744
rect 260741 63686 263475 63688
rect 260741 63683 260807 63686
rect 263409 63683 263475 63686
rect 263593 63746 263659 63749
rect 273069 63746 273135 63749
rect 263593 63744 273135 63746
rect 263593 63688 263598 63744
rect 263654 63688 273074 63744
rect 273130 63688 273135 63744
rect 263593 63686 273135 63688
rect 263593 63683 263659 63686
rect 273069 63683 273135 63686
rect 273253 63746 273319 63749
rect 280102 63746 280108 63748
rect 273253 63744 280108 63746
rect 273253 63688 273258 63744
rect 273314 63688 280108 63744
rect 273253 63686 280108 63688
rect 273253 63683 273319 63686
rect 280102 63684 280108 63686
rect 280172 63684 280178 63748
rect 237230 63548 237236 63612
rect 237300 63610 237306 63612
rect 260741 63610 260807 63613
rect 327022 63610 327028 63612
rect 237300 63608 260807 63610
rect 237300 63552 260746 63608
rect 260802 63552 260807 63608
rect 237300 63550 260807 63552
rect 237300 63548 237306 63550
rect 260741 63547 260807 63550
rect 285078 63550 309058 63610
rect 280102 63412 280108 63476
rect 280172 63474 280178 63476
rect 285078 63474 285138 63550
rect 280172 63414 285138 63474
rect 308998 63474 309058 63550
rect 317278 63550 327028 63610
rect 317278 63474 317338 63550
rect 327022 63548 327028 63550
rect 327092 63548 327098 63612
rect 340830 63610 340890 63822
rect 376661 63880 378567 63882
rect 376661 63824 376666 63880
rect 376722 63824 378506 63880
rect 378562 63824 378567 63880
rect 376661 63822 378567 63824
rect 376661 63819 376727 63822
rect 378501 63819 378567 63822
rect 386321 63882 386387 63885
rect 386321 63880 389098 63882
rect 386321 63824 386326 63880
rect 386382 63824 389098 63880
rect 386321 63822 389098 63824
rect 386321 63819 386387 63822
rect 367093 63746 367159 63749
rect 350582 63744 367159 63746
rect 350582 63688 367098 63744
rect 367154 63688 367159 63744
rect 350582 63686 367159 63688
rect 350582 63610 350642 63686
rect 367093 63683 367159 63686
rect 340830 63550 350642 63610
rect 389038 63610 389098 63822
rect 398606 63746 398666 63958
rect 405406 63956 405412 63958
rect 405476 63956 405482 64020
rect 470550 63822 480178 63882
rect 417877 63746 417943 63749
rect 389222 63686 398666 63746
rect 408542 63744 417943 63746
rect 408542 63688 417882 63744
rect 417938 63688 417943 63744
rect 408542 63686 417943 63688
rect 389222 63610 389282 63686
rect 389038 63550 389282 63610
rect 405590 63548 405596 63612
rect 405660 63610 405666 63612
rect 408542 63610 408602 63686
rect 417877 63683 417943 63686
rect 418153 63746 418219 63749
rect 437197 63746 437263 63749
rect 418153 63744 424978 63746
rect 418153 63688 418158 63744
rect 418214 63688 424978 63744
rect 418153 63686 424978 63688
rect 418153 63683 418219 63686
rect 405660 63550 408602 63610
rect 424918 63610 424978 63686
rect 427862 63744 437263 63746
rect 427862 63688 437202 63744
rect 437258 63688 437263 63744
rect 427862 63686 437263 63688
rect 427862 63610 427922 63686
rect 437197 63683 437263 63686
rect 437473 63746 437539 63749
rect 456517 63746 456583 63749
rect 437473 63744 444298 63746
rect 437473 63688 437478 63744
rect 437534 63688 444298 63744
rect 437473 63686 444298 63688
rect 437473 63683 437539 63686
rect 424918 63550 427922 63610
rect 444238 63610 444298 63686
rect 447182 63744 456583 63746
rect 447182 63688 456522 63744
rect 456578 63688 456583 63744
rect 447182 63686 456583 63688
rect 447182 63610 447242 63686
rect 456517 63683 456583 63686
rect 456885 63746 456951 63749
rect 456885 63744 466378 63746
rect 456885 63688 456890 63744
rect 456946 63688 466378 63744
rect 456885 63686 466378 63688
rect 456885 63683 456951 63686
rect 444238 63550 447242 63610
rect 466318 63610 466378 63686
rect 470550 63610 470610 63822
rect 466318 63550 470610 63610
rect 480118 63610 480178 63822
rect 480302 63822 489930 63882
rect 480302 63610 480362 63822
rect 489870 63746 489930 63822
rect 499622 63822 509250 63882
rect 489870 63686 499498 63746
rect 480118 63550 480362 63610
rect 499438 63610 499498 63686
rect 499622 63610 499682 63822
rect 509190 63746 509250 63822
rect 518942 63822 528570 63882
rect 509190 63686 518818 63746
rect 499438 63550 499682 63610
rect 518758 63610 518818 63686
rect 518942 63610 519002 63822
rect 528510 63746 528570 63822
rect 538262 63822 547890 63882
rect 528510 63686 538138 63746
rect 518758 63550 519002 63610
rect 538078 63610 538138 63686
rect 538262 63610 538322 63822
rect 547830 63746 547890 63822
rect 557582 63822 567210 63882
rect 547830 63686 557458 63746
rect 538078 63550 538322 63610
rect 557398 63610 557458 63686
rect 557582 63610 557642 63822
rect 567150 63746 567210 63822
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 567150 63686 576778 63746
rect 557398 63550 557642 63610
rect 576718 63610 576778 63686
rect 576902 63686 583402 63746
rect 576902 63610 576962 63686
rect 576718 63550 576962 63610
rect 405660 63548 405666 63550
rect 308998 63414 317338 63474
rect 280172 63412 280178 63414
rect 337193 56810 337259 56813
rect 337150 56808 337259 56810
rect 337150 56752 337198 56808
rect 337254 56752 337259 56808
rect 337150 56747 337259 56752
rect 337150 56674 337210 56747
rect 337285 56674 337351 56677
rect 337150 56672 337351 56674
rect 337150 56616 337290 56672
rect 337346 56616 337351 56672
rect 337150 56614 337351 56616
rect 337285 56611 337351 56614
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 2773 50146 2839 50149
rect -960 50144 2839 50146
rect -960 50088 2778 50144
rect 2834 50088 2839 50144
rect -960 50086 2839 50088
rect -960 49996 480 50086
rect 2773 50083 2839 50086
rect 251449 48514 251515 48517
rect 251222 48512 251515 48514
rect 251222 48456 251454 48512
rect 251510 48456 251515 48512
rect 251222 48454 251515 48456
rect 232313 48378 232379 48381
rect 232270 48376 232379 48378
rect 232270 48320 232318 48376
rect 232374 48320 232379 48376
rect 232270 48315 232379 48320
rect 251222 48378 251282 48454
rect 251449 48451 251515 48454
rect 251357 48378 251423 48381
rect 251222 48376 251423 48378
rect 251222 48320 251362 48376
rect 251418 48320 251423 48376
rect 251222 48318 251423 48320
rect 251357 48315 251423 48318
rect 232270 47973 232330 48315
rect 232270 47968 232379 47973
rect 232270 47912 232318 47968
rect 232374 47912 232379 47968
rect 232270 47910 232379 47912
rect 232313 47907 232379 47910
rect 310881 45658 310947 45661
rect 311065 45658 311131 45661
rect 310881 45656 311131 45658
rect 310881 45600 310886 45656
rect 310942 45600 311070 45656
rect 311126 45600 311131 45656
rect 310881 45598 311131 45600
rect 310881 45595 310947 45598
rect 311065 45595 311131 45598
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 396030 40430 405658 40490
rect 239998 40294 251098 40354
rect 232998 40156 233004 40220
rect 233068 40218 233074 40220
rect 239998 40218 240058 40294
rect 233068 40158 240058 40218
rect 251038 40218 251098 40294
rect 251222 40294 254594 40354
rect 251222 40218 251282 40294
rect 251038 40158 251282 40218
rect 254534 40218 254594 40294
rect 327022 40292 327028 40356
rect 327092 40354 327098 40356
rect 376661 40354 376727 40357
rect 327092 40294 340890 40354
rect 327092 40292 327098 40294
rect 273069 40218 273135 40221
rect 254534 40216 273135 40218
rect 254534 40160 273074 40216
rect 273130 40160 273135 40216
rect 254534 40158 273135 40160
rect 233068 40156 233074 40158
rect 273069 40155 273135 40158
rect 273253 40218 273319 40221
rect 282729 40218 282795 40221
rect 273253 40216 282795 40218
rect 273253 40160 273258 40216
rect 273314 40160 282734 40216
rect 282790 40160 282795 40216
rect 273253 40158 282795 40160
rect 273253 40155 273319 40158
rect 282729 40155 282795 40158
rect 282913 40218 282979 40221
rect 306373 40218 306439 40221
rect 282913 40216 306439 40218
rect 282913 40160 282918 40216
rect 282974 40160 306378 40216
rect 306434 40160 306439 40216
rect 282913 40158 306439 40160
rect 282913 40155 282979 40158
rect 306373 40155 306439 40158
rect 315941 40082 316007 40085
rect 327022 40082 327028 40084
rect 315941 40080 327028 40082
rect 315941 40024 315946 40080
rect 316002 40024 327028 40080
rect 315941 40022 327028 40024
rect 315941 40019 316007 40022
rect 327022 40020 327028 40022
rect 327092 40020 327098 40084
rect 340830 40082 340890 40294
rect 376661 40352 394618 40354
rect 376661 40296 376666 40352
rect 376722 40296 394618 40352
rect 376661 40294 394618 40296
rect 376661 40291 376727 40294
rect 367093 40218 367159 40221
rect 350582 40216 367159 40218
rect 350582 40160 367098 40216
rect 367154 40160 367159 40216
rect 350582 40158 367159 40160
rect 394558 40218 394618 40294
rect 396030 40218 396090 40430
rect 405598 40356 405658 40430
rect 405590 40292 405596 40356
rect 405660 40292 405666 40356
rect 470550 40294 480178 40354
rect 417877 40218 417943 40221
rect 394558 40158 396090 40218
rect 408542 40216 417943 40218
rect 408542 40160 417882 40216
rect 417938 40160 417943 40216
rect 408542 40158 417943 40160
rect 350582 40082 350642 40158
rect 367093 40155 367159 40158
rect 340830 40022 350642 40082
rect 405590 40020 405596 40084
rect 405660 40082 405666 40084
rect 408542 40082 408602 40158
rect 417877 40155 417943 40158
rect 420361 40218 420427 40221
rect 437197 40218 437263 40221
rect 420361 40216 424978 40218
rect 420361 40160 420366 40216
rect 420422 40160 424978 40216
rect 420361 40158 424978 40160
rect 420361 40155 420427 40158
rect 405660 40022 408602 40082
rect 424918 40082 424978 40158
rect 427862 40216 437263 40218
rect 427862 40160 437202 40216
rect 437258 40160 437263 40216
rect 427862 40158 437263 40160
rect 427862 40082 427922 40158
rect 437197 40155 437263 40158
rect 437473 40218 437539 40221
rect 456517 40218 456583 40221
rect 437473 40216 444298 40218
rect 437473 40160 437478 40216
rect 437534 40160 444298 40216
rect 437473 40158 444298 40160
rect 437473 40155 437539 40158
rect 424918 40022 427922 40082
rect 444238 40082 444298 40158
rect 447182 40216 456583 40218
rect 447182 40160 456522 40216
rect 456578 40160 456583 40216
rect 447182 40158 456583 40160
rect 447182 40082 447242 40158
rect 456517 40155 456583 40158
rect 456885 40218 456951 40221
rect 456885 40216 466378 40218
rect 456885 40160 456890 40216
rect 456946 40160 466378 40216
rect 456885 40158 466378 40160
rect 456885 40155 456951 40158
rect 444238 40022 447242 40082
rect 466318 40082 466378 40158
rect 470550 40082 470610 40294
rect 466318 40022 470610 40082
rect 480118 40082 480178 40294
rect 480302 40294 489930 40354
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 405660 40020 405666 40022
rect 285949 38858 286015 38861
rect 285949 38856 286058 38858
rect 285949 38800 285954 38856
rect 286010 38800 286058 38856
rect 285949 38795 286058 38800
rect 285998 38589 286058 38795
rect 285949 38584 286058 38589
rect 285949 38528 285954 38584
rect 286010 38528 286058 38584
rect 285949 38526 286058 38528
rect 285949 38523 286015 38526
rect 386505 37362 386571 37365
rect 386689 37362 386755 37365
rect 386505 37360 386755 37362
rect 386505 37304 386510 37360
rect 386566 37304 386694 37360
rect 386750 37304 386755 37360
rect 386505 37302 386755 37304
rect 386505 37299 386571 37302
rect 386689 37299 386755 37302
rect -960 35866 480 35956
rect 3141 35866 3207 35869
rect -960 35864 3207 35866
rect -960 35808 3146 35864
rect 3202 35808 3207 35864
rect -960 35806 3207 35808
rect -960 35716 480 35806
rect 3141 35803 3207 35806
rect 287094 29548 287100 29612
rect 287164 29610 287170 29612
rect 296621 29610 296687 29613
rect 331857 29610 331923 29613
rect 287164 29608 296687 29610
rect 287164 29552 296626 29608
rect 296682 29552 296687 29608
rect 287164 29550 296687 29552
rect 287164 29548 287170 29550
rect 296621 29547 296687 29550
rect 327030 29608 331923 29610
rect 327030 29552 331862 29608
rect 331918 29552 331923 29608
rect 327030 29550 331923 29552
rect 249742 29412 249748 29476
rect 249812 29474 249818 29476
rect 249812 29414 254042 29474
rect 249812 29412 249818 29414
rect 253982 29338 254042 29414
rect 265390 29414 270418 29474
rect 265390 29338 265450 29414
rect 253982 29278 265450 29338
rect 270358 29338 270418 29414
rect 270542 29414 273914 29474
rect 270542 29338 270602 29414
rect 270358 29278 270602 29338
rect 273854 29338 273914 29414
rect 278773 29338 278839 29341
rect 273854 29336 278839 29338
rect 273854 29280 278778 29336
rect 278834 29280 278839 29336
rect 273854 29278 278839 29280
rect 278773 29275 278839 29278
rect 296621 29338 296687 29341
rect 298093 29338 298159 29341
rect 296621 29336 298159 29338
rect 296621 29280 296626 29336
rect 296682 29280 298098 29336
rect 298154 29280 298159 29336
rect 296621 29278 298159 29280
rect 296621 29275 296687 29278
rect 298093 29275 298159 29278
rect 317321 29338 317387 29341
rect 322197 29338 322263 29341
rect 327030 29338 327090 29550
rect 331857 29547 331923 29550
rect 405590 29474 405596 29476
rect 398606 29414 405596 29474
rect 317321 29336 317522 29338
rect 317321 29280 317326 29336
rect 317382 29280 317522 29336
rect 317321 29278 317522 29280
rect 317321 29275 317387 29278
rect 235758 29140 235764 29204
rect 235828 29202 235834 29204
rect 240133 29202 240199 29205
rect 235828 29200 240199 29202
rect 235828 29144 240138 29200
rect 240194 29144 240199 29200
rect 235828 29142 240199 29144
rect 235828 29140 235834 29142
rect 240133 29139 240199 29142
rect 281257 29202 281323 29205
rect 287094 29202 287100 29204
rect 281257 29200 287100 29202
rect 281257 29144 281262 29200
rect 281318 29144 287100 29200
rect 281257 29142 287100 29144
rect 281257 29139 281323 29142
rect 287094 29140 287100 29142
rect 287164 29140 287170 29204
rect 249701 29066 249767 29069
rect 317462 29066 317522 29278
rect 322197 29336 327090 29338
rect 322197 29280 322202 29336
rect 322258 29280 327090 29336
rect 322197 29278 327090 29280
rect 331857 29338 331923 29341
rect 357341 29338 357407 29341
rect 376661 29338 376727 29341
rect 331857 29336 340890 29338
rect 331857 29280 331862 29336
rect 331918 29280 340890 29336
rect 331857 29278 340890 29280
rect 322197 29275 322263 29278
rect 331857 29275 331923 29278
rect 322197 29066 322263 29069
rect 249620 29064 249810 29066
rect 249620 29008 249706 29064
rect 249762 29008 249810 29064
rect 249620 29006 249810 29008
rect 317462 29064 322263 29066
rect 317462 29008 322202 29064
rect 322258 29008 322263 29064
rect 317462 29006 322263 29008
rect 340830 29066 340890 29278
rect 357341 29336 360210 29338
rect 357341 29280 357346 29336
rect 357402 29280 360210 29336
rect 357341 29278 360210 29280
rect 357341 29275 357407 29278
rect 347773 29066 347839 29069
rect 340830 29064 347839 29066
rect 340830 29008 347778 29064
rect 347834 29008 347839 29064
rect 340830 29006 347839 29008
rect 360150 29066 360210 29278
rect 376661 29336 379530 29338
rect 376661 29280 376666 29336
rect 376722 29280 379530 29336
rect 376661 29278 379530 29280
rect 376661 29275 376727 29278
rect 367093 29066 367159 29069
rect 360150 29064 367159 29066
rect 360150 29008 367098 29064
rect 367154 29008 367159 29064
rect 360150 29006 367159 29008
rect 379470 29066 379530 29278
rect 398606 29202 398666 29414
rect 405590 29412 405596 29414
rect 405660 29412 405666 29476
rect 481582 29412 481588 29476
rect 481652 29474 481658 29476
rect 491201 29474 491267 29477
rect 481652 29472 491267 29474
rect 481652 29416 491206 29472
rect 491262 29416 491267 29472
rect 481652 29414 491267 29416
rect 481652 29412 481658 29414
rect 491201 29411 491267 29414
rect 476021 29338 476087 29341
rect 466502 29336 476087 29338
rect 466502 29280 476026 29336
rect 476082 29280 476087 29336
rect 466502 29278 476087 29280
rect 437197 29202 437263 29205
rect 389222 29142 398666 29202
rect 408542 29142 424978 29202
rect 389222 29066 389282 29142
rect 379470 29006 389282 29066
rect 249701 29003 249810 29006
rect 322197 29003 322263 29006
rect 347773 29003 347839 29006
rect 367093 29003 367159 29006
rect 405590 29004 405596 29068
rect 405660 29066 405666 29068
rect 408542 29066 408602 29142
rect 405660 29006 408602 29066
rect 424918 29066 424978 29142
rect 427862 29200 437263 29202
rect 427862 29144 437202 29200
rect 437258 29144 437263 29200
rect 427862 29142 437263 29144
rect 427862 29066 427922 29142
rect 437197 29139 437263 29142
rect 437473 29202 437539 29205
rect 456517 29202 456583 29205
rect 437473 29200 444298 29202
rect 437473 29144 437478 29200
rect 437534 29144 444298 29200
rect 437473 29142 444298 29144
rect 437473 29139 437539 29142
rect 424918 29006 427922 29066
rect 444238 29066 444298 29142
rect 447182 29200 456583 29202
rect 447182 29144 456522 29200
rect 456578 29144 456583 29200
rect 447182 29142 456583 29144
rect 447182 29066 447242 29142
rect 456517 29139 456583 29142
rect 456793 29202 456859 29205
rect 456793 29200 463618 29202
rect 456793 29144 456798 29200
rect 456854 29144 463618 29200
rect 456793 29142 463618 29144
rect 456793 29139 456859 29142
rect 444238 29006 447242 29066
rect 463558 29066 463618 29142
rect 466502 29066 466562 29278
rect 476021 29275 476087 29278
rect 502241 29338 502307 29341
rect 583520 29338 584960 29428
rect 502241 29336 509250 29338
rect 502241 29280 502246 29336
rect 502302 29280 509250 29336
rect 502241 29278 509250 29280
rect 502241 29275 502307 29278
rect 476205 29202 476271 29205
rect 481582 29202 481588 29204
rect 476205 29200 481588 29202
rect 476205 29144 476210 29200
rect 476266 29144 481588 29200
rect 476205 29142 481588 29144
rect 476205 29139 476271 29142
rect 481582 29140 481588 29142
rect 481652 29140 481658 29204
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 463558 29006 466562 29066
rect 491201 29066 491267 29069
rect 492765 29066 492831 29069
rect 491201 29064 492831 29066
rect 491201 29008 491206 29064
rect 491262 29008 492770 29064
rect 492826 29008 492831 29064
rect 491201 29006 492831 29008
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 405660 29004 405666 29006
rect 491201 29003 491267 29006
rect 492765 29003 492831 29006
rect 249750 28932 249810 29003
rect 249742 28868 249748 28932
rect 249812 28868 249818 28932
rect 298093 28930 298159 28933
rect 306373 28930 306439 28933
rect 298093 28928 306439 28930
rect 298093 28872 298098 28928
rect 298154 28872 306378 28928
rect 306434 28872 306439 28928
rect 298093 28870 306439 28872
rect 298093 28867 298159 28870
rect 306373 28867 306439 28870
rect 315941 28930 316007 28933
rect 317321 28930 317387 28933
rect 330109 28930 330175 28933
rect 315941 28928 317387 28930
rect 315941 28872 315946 28928
rect 316002 28872 317326 28928
rect 317382 28872 317387 28928
rect 315941 28870 317387 28872
rect 315941 28867 316007 28870
rect 317321 28867 317387 28870
rect 329974 28928 330175 28930
rect 329974 28872 330114 28928
rect 330170 28872 330175 28928
rect 329974 28870 330175 28872
rect 329974 28794 330034 28870
rect 330109 28867 330175 28870
rect 330201 28794 330267 28797
rect 329974 28792 330267 28794
rect 329974 28736 330206 28792
rect 330262 28736 330267 28792
rect 329974 28734 330267 28736
rect 330201 28731 330267 28734
rect 251173 27706 251239 27709
rect 251357 27706 251423 27709
rect 251173 27704 251423 27706
rect 251173 27648 251178 27704
rect 251234 27648 251362 27704
rect 251418 27648 251423 27704
rect 251173 27646 251423 27648
rect 251173 27643 251239 27646
rect 251357 27643 251423 27646
rect 357617 27706 357683 27709
rect 357801 27706 357867 27709
rect 357617 27704 357867 27706
rect 357617 27648 357622 27704
rect 357678 27648 357806 27704
rect 357862 27648 357867 27704
rect 357617 27646 357867 27648
rect 357617 27643 357683 27646
rect 357801 27643 357867 27646
rect 465574 21994 465580 21996
rect 614 21934 465580 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 465574 21932 465580 21934
rect 465644 21932 465650 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 376702 17172 376708 17236
rect 376772 17234 376778 17236
rect 386321 17234 386387 17237
rect 376772 17232 386387 17234
rect 376772 17176 386326 17232
rect 386382 17176 386387 17232
rect 376772 17174 386387 17176
rect 376772 17172 376778 17174
rect 386321 17171 386387 17174
rect 249742 17036 249748 17100
rect 249812 17098 249818 17100
rect 259361 17098 259427 17101
rect 336641 17098 336707 17101
rect 396022 17098 396028 17100
rect 249812 17096 259427 17098
rect 249812 17040 259366 17096
rect 259422 17040 259427 17096
rect 249812 17038 259427 17040
rect 249812 17036 249818 17038
rect 259361 17035 259427 17038
rect 327030 17096 336707 17098
rect 327030 17040 336646 17096
rect 336702 17040 336707 17096
rect 327030 17038 336707 17040
rect 249742 16826 249748 16828
rect 239998 16766 249748 16826
rect 231710 16628 231716 16692
rect 231780 16690 231786 16692
rect 239998 16690 240058 16766
rect 249742 16764 249748 16766
rect 249812 16764 249818 16828
rect 260966 16764 260972 16828
rect 261036 16826 261042 16828
rect 298001 16826 298067 16829
rect 261036 16766 273178 16826
rect 261036 16764 261042 16766
rect 231780 16630 240058 16690
rect 259361 16690 259427 16693
rect 260782 16690 260788 16692
rect 259361 16688 260788 16690
rect 259361 16632 259366 16688
rect 259422 16632 260788 16688
rect 259361 16630 260788 16632
rect 231780 16628 231786 16630
rect 259361 16627 259427 16630
rect 260782 16628 260788 16630
rect 260852 16628 260858 16692
rect 273118 16690 273178 16766
rect 295382 16824 298067 16826
rect 295382 16768 298006 16824
rect 298062 16768 298067 16824
rect 295382 16766 298067 16768
rect 290549 16690 290615 16693
rect 295382 16690 295442 16766
rect 298001 16763 298067 16766
rect 325601 16826 325667 16829
rect 327030 16826 327090 17038
rect 336641 17035 336707 17038
rect 389222 17038 396028 17098
rect 347773 16962 347839 16965
rect 325601 16824 327090 16826
rect 325601 16768 325606 16824
rect 325662 16768 327090 16824
rect 325601 16766 327090 16768
rect 340830 16960 347839 16962
rect 340830 16904 347778 16960
rect 347834 16904 347839 16960
rect 340830 16902 347839 16904
rect 325601 16763 325667 16766
rect 273118 16630 273362 16690
rect 273302 16554 273362 16630
rect 290549 16688 295442 16690
rect 290549 16632 290554 16688
rect 290610 16632 295442 16688
rect 290549 16630 295442 16632
rect 298093 16690 298159 16693
rect 304758 16690 304764 16692
rect 298093 16688 304764 16690
rect 298093 16632 298098 16688
rect 298154 16632 304764 16688
rect 298093 16630 304764 16632
rect 290549 16627 290615 16630
rect 298093 16627 298159 16630
rect 304758 16628 304764 16630
rect 304828 16628 304834 16692
rect 320817 16690 320883 16693
rect 312126 16688 320883 16690
rect 312126 16632 320822 16688
rect 320878 16632 320883 16688
rect 312126 16630 320883 16632
rect 278773 16554 278839 16557
rect 273302 16552 278839 16554
rect 273302 16496 278778 16552
rect 278834 16496 278839 16552
rect 273302 16494 278839 16496
rect 278773 16491 278839 16494
rect 304942 16492 304948 16556
rect 305012 16554 305018 16556
rect 312126 16554 312186 16630
rect 320817 16627 320883 16630
rect 336641 16690 336707 16693
rect 340830 16690 340890 16902
rect 347773 16899 347839 16902
rect 357382 16900 357388 16964
rect 357452 16962 357458 16964
rect 367001 16962 367067 16965
rect 357452 16960 367067 16962
rect 357452 16904 367006 16960
rect 367062 16904 367067 16960
rect 357452 16902 367067 16904
rect 357452 16900 357458 16902
rect 367001 16899 367067 16902
rect 376661 16964 376727 16965
rect 376661 16960 376708 16964
rect 376772 16962 376778 16964
rect 376661 16904 376666 16960
rect 376661 16900 376708 16904
rect 376772 16902 376854 16962
rect 376772 16900 376778 16902
rect 376661 16899 376727 16900
rect 367001 16826 367067 16829
rect 369669 16826 369735 16829
rect 367001 16824 369735 16826
rect 367001 16768 367006 16824
rect 367062 16768 369674 16824
rect 369730 16768 369735 16824
rect 367001 16766 369735 16768
rect 367001 16763 367067 16766
rect 369669 16763 369735 16766
rect 386321 16826 386387 16829
rect 389222 16826 389282 17038
rect 396022 17036 396028 17038
rect 396092 17036 396098 17100
rect 487797 17098 487863 17101
rect 483062 17096 487863 17098
rect 483062 17040 487802 17096
rect 487858 17040 487863 17096
rect 483062 17038 487863 17040
rect 456517 16962 456583 16965
rect 447182 16960 456583 16962
rect 447182 16904 456522 16960
rect 456578 16904 456583 16960
rect 447182 16902 456583 16904
rect 437197 16826 437263 16829
rect 386321 16824 389282 16826
rect 386321 16768 386326 16824
rect 386382 16768 389282 16824
rect 386321 16766 389282 16768
rect 408542 16766 424978 16826
rect 386321 16763 386387 16766
rect 336641 16688 340890 16690
rect 336641 16632 336646 16688
rect 336702 16632 340890 16688
rect 336641 16630 340890 16632
rect 352649 16690 352715 16693
rect 357382 16690 357388 16692
rect 352649 16688 357388 16690
rect 352649 16632 352654 16688
rect 352710 16632 357388 16688
rect 352649 16630 357388 16632
rect 336641 16627 336707 16630
rect 352649 16627 352715 16630
rect 357382 16628 357388 16630
rect 357452 16628 357458 16692
rect 396022 16628 396028 16692
rect 396092 16690 396098 16692
rect 398741 16690 398807 16693
rect 396092 16688 398807 16690
rect 396092 16632 398746 16688
rect 398802 16632 398807 16688
rect 396092 16630 398807 16632
rect 396092 16628 396098 16630
rect 398741 16627 398807 16630
rect 398925 16690 398991 16693
rect 408542 16690 408602 16766
rect 398925 16688 408602 16690
rect 398925 16632 398930 16688
rect 398986 16632 408602 16688
rect 398925 16630 408602 16632
rect 424918 16690 424978 16766
rect 427862 16824 437263 16826
rect 427862 16768 437202 16824
rect 437258 16768 437263 16824
rect 427862 16766 437263 16768
rect 427862 16690 427922 16766
rect 437197 16763 437263 16766
rect 437473 16826 437539 16829
rect 437473 16824 444298 16826
rect 437473 16768 437478 16824
rect 437534 16768 444298 16824
rect 437473 16766 444298 16768
rect 437473 16763 437539 16766
rect 424918 16630 427922 16690
rect 444238 16690 444298 16766
rect 447182 16690 447242 16902
rect 456517 16899 456583 16902
rect 457437 16826 457503 16829
rect 475561 16826 475627 16829
rect 457437 16824 475627 16826
rect 457437 16768 457442 16824
rect 457498 16768 475566 16824
rect 475622 16768 475627 16824
rect 457437 16766 475627 16768
rect 457437 16763 457503 16766
rect 475561 16763 475627 16766
rect 482921 16826 482987 16829
rect 483062 16826 483122 17038
rect 487797 17035 487863 17038
rect 492622 16900 492628 16964
rect 492692 16962 492698 16964
rect 492692 16902 509250 16962
rect 492692 16900 492698 16902
rect 482921 16824 483122 16826
rect 482921 16768 482926 16824
rect 482982 16768 483122 16824
rect 482921 16766 483122 16768
rect 509190 16826 509250 16902
rect 518942 16902 528570 16962
rect 509190 16766 518818 16826
rect 482921 16763 482987 16766
rect 444238 16630 447242 16690
rect 487797 16690 487863 16693
rect 492622 16690 492628 16692
rect 487797 16688 492628 16690
rect 487797 16632 487802 16688
rect 487858 16632 492628 16688
rect 487797 16630 492628 16632
rect 398925 16627 398991 16630
rect 487797 16627 487863 16630
rect 492622 16628 492628 16630
rect 492692 16628 492698 16692
rect 518758 16690 518818 16766
rect 518942 16690 519002 16902
rect 528510 16826 528570 16902
rect 538262 16902 547890 16962
rect 528510 16766 538138 16826
rect 518758 16630 519002 16690
rect 538078 16690 538138 16766
rect 538262 16690 538322 16902
rect 547830 16826 547890 16902
rect 557582 16902 567210 16962
rect 547830 16766 557458 16826
rect 538078 16630 538322 16690
rect 557398 16690 557458 16766
rect 557582 16690 557642 16902
rect 567150 16826 567210 16902
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 567150 16766 576778 16826
rect 557398 16630 557642 16690
rect 576718 16690 576778 16766
rect 576902 16766 583402 16826
rect 576902 16690 576962 16766
rect 576718 16630 576962 16690
rect 305012 16494 312186 16554
rect 305012 16492 305018 16494
rect 3141 11658 3207 11661
rect 466494 11658 466500 11660
rect 3141 11656 466500 11658
rect 3141 11600 3146 11656
rect 3202 11600 466500 11656
rect 3141 11598 466500 11600
rect 3141 11595 3207 11598
rect 466494 11596 466500 11598
rect 466564 11596 466570 11660
rect 376753 9618 376819 9621
rect 377029 9618 377095 9621
rect 376753 9616 377095 9618
rect 376753 9560 376758 9616
rect 376814 9560 377034 9616
rect 377090 9560 377095 9616
rect 376753 9558 377095 9560
rect 376753 9555 376819 9558
rect 377029 9555 377095 9558
rect 132585 8938 132651 8941
rect 284477 8938 284543 8941
rect 132585 8936 284543 8938
rect 132585 8880 132590 8936
rect 132646 8880 284482 8936
rect 284538 8880 284543 8936
rect 132585 8878 284543 8880
rect 132585 8875 132651 8878
rect 284477 8875 284543 8878
rect 128997 7578 129063 7581
rect 283097 7578 283163 7581
rect 128997 7576 283163 7578
rect 128997 7520 129002 7576
rect 129058 7520 283102 7576
rect 283158 7520 283163 7576
rect 128997 7518 283163 7520
rect 128997 7515 129063 7518
rect 283097 7515 283163 7518
rect -960 7170 480 7260
rect 3141 7170 3207 7173
rect -960 7168 3207 7170
rect -960 7112 3146 7168
rect 3202 7112 3207 7168
rect -960 7110 3207 7112
rect -960 7020 480 7110
rect 3141 7107 3207 7110
rect 51625 6218 51691 6221
rect 249977 6218 250043 6221
rect 51625 6216 250043 6218
rect 51625 6160 51630 6216
rect 51686 6160 249982 6216
rect 250038 6160 250043 6216
rect 51625 6158 250043 6160
rect 51625 6155 51691 6158
rect 249977 6155 250043 6158
rect 583520 5796 584960 6036
rect 312077 4994 312143 4997
rect 315941 4994 316007 4997
rect 312077 4992 316007 4994
rect 312077 4936 312082 4992
rect 312138 4936 315946 4992
rect 316002 4936 316007 4992
rect 312077 4934 316007 4936
rect 312077 4931 312143 4934
rect 315941 4931 316007 4934
rect 208669 4858 208735 4861
rect 314653 4858 314719 4861
rect 208669 4856 314719 4858
rect 208669 4800 208674 4856
rect 208730 4800 314658 4856
rect 314714 4800 314719 4856
rect 208669 4798 314719 4800
rect 208669 4795 208735 4798
rect 314653 4795 314719 4798
rect 467741 4858 467807 4861
rect 576209 4858 576275 4861
rect 467741 4856 576275 4858
rect 467741 4800 467746 4856
rect 467802 4800 576214 4856
rect 576270 4800 576275 4856
rect 467741 4798 576275 4800
rect 467741 4795 467807 4798
rect 576209 4795 576275 4798
rect 420729 3770 420795 3773
rect 434529 3770 434595 3773
rect 420729 3768 434595 3770
rect 420729 3712 420734 3768
rect 420790 3712 434534 3768
rect 434590 3712 434595 3768
rect 420729 3710 434595 3712
rect 420729 3707 420795 3710
rect 434529 3707 434595 3710
rect 6453 3362 6519 3365
rect 232037 3362 232103 3365
rect 6453 3360 232103 3362
rect 6453 3304 6458 3360
rect 6514 3304 232042 3360
rect 232098 3304 232103 3360
rect 6453 3302 232103 3304
rect 6453 3299 6519 3302
rect 232037 3299 232103 3302
rect 307385 3362 307451 3365
rect 356237 3362 356303 3365
rect 307385 3360 356303 3362
rect 307385 3304 307390 3360
rect 307446 3304 356242 3360
rect 356298 3304 356303 3360
rect 307385 3302 356303 3304
rect 307385 3299 307451 3302
rect 356237 3299 356303 3302
rect 468753 3362 468819 3365
rect 580993 3362 581059 3365
rect 468753 3360 581059 3362
rect 468753 3304 468758 3360
rect 468814 3304 580998 3360
rect 581054 3304 581059 3360
rect 468753 3302 581059 3304
rect 468753 3299 468819 3302
rect 580993 3299 581059 3302
<< via3 >>
rect 465948 583340 466012 583404
rect 465764 583204 465828 583268
rect 239444 583068 239508 583132
rect 239260 582932 239324 582996
rect 465580 579668 465644 579732
rect 231716 579260 231780 579324
rect 233004 579320 233068 579324
rect 233004 579264 233018 579320
rect 233018 579264 233068 579320
rect 233004 579260 233068 579264
rect 235764 579260 235828 579324
rect 237236 579320 237300 579324
rect 237236 579264 237250 579320
rect 237250 579264 237300 579320
rect 237236 579260 237300 579264
rect 239996 579260 240060 579324
rect 241284 579260 241348 579324
rect 249564 579320 249628 579324
rect 249564 579264 249578 579320
rect 249578 579264 249628 579320
rect 249564 579260 249628 579264
rect 466500 579320 466564 579324
rect 466500 579264 466514 579320
rect 466514 579264 466564 579320
rect 466500 579260 466564 579264
rect 465948 533020 466012 533084
rect 465764 486100 465828 486164
rect 239444 337996 239508 338060
rect 249380 334188 249444 334252
rect 249380 328442 249444 328506
rect 249380 322220 249444 322284
rect 249012 317460 249076 317524
rect 249012 309164 249076 309228
rect 249196 308892 249260 308956
rect 249196 302228 249260 302292
rect 249196 302092 249260 302156
rect 341380 299372 341444 299436
rect 249196 298072 249260 298076
rect 249196 298016 249246 298072
rect 249246 298016 249260 298072
rect 249196 298012 249260 298016
rect 239260 295156 239324 295220
rect 341380 289852 341444 289916
rect 249380 288492 249444 288556
rect 249380 288356 249444 288420
rect 341380 280060 341444 280124
rect 249196 279032 249260 279036
rect 249196 278976 249246 279032
rect 249246 278976 249260 279032
rect 249196 278972 249260 278976
rect 249196 277340 249260 277404
rect 336964 273940 337028 274004
rect 341380 270540 341444 270604
rect 236316 270464 236380 270468
rect 236316 270408 236330 270464
rect 236330 270408 236380 270464
rect 236316 270404 236380 270408
rect 249380 267880 249444 267884
rect 249380 267824 249430 267880
rect 249430 267824 249444 267880
rect 249380 267820 249444 267824
rect 249380 263740 249444 263804
rect 249196 263468 249260 263532
rect 236316 260884 236380 260948
rect 341380 260748 341444 260812
rect 336964 260672 337028 260676
rect 336964 260616 336978 260672
rect 336978 260616 337028 260672
rect 336964 260612 337028 260616
rect 341380 251228 341444 251292
rect 249380 241844 249444 241908
rect 249196 241708 249260 241772
rect 249196 241436 249260 241500
rect 249380 240892 249444 240956
rect 249380 224980 249444 225044
rect 249564 224708 249628 224772
rect 366956 222184 367020 222188
rect 366956 222128 367006 222184
rect 367006 222128 367020 222184
rect 366956 222124 367020 222128
rect 236316 221988 236380 222052
rect 358860 220764 358924 220828
rect 249196 217364 249260 217428
rect 249564 217364 249628 217428
rect 236316 212664 236380 212668
rect 236316 212608 236330 212664
rect 236330 212608 236380 212664
rect 236316 212604 236380 212608
rect 366956 212664 367020 212668
rect 366956 212608 367006 212664
rect 367006 212608 367020 212664
rect 366956 212604 367020 212608
rect 249196 212528 249260 212532
rect 249196 212472 249246 212528
rect 249246 212472 249260 212528
rect 249196 212468 249260 212472
rect 358860 211108 358924 211172
rect 249564 205396 249628 205460
rect 236316 202812 236380 202876
rect 249564 202872 249628 202876
rect 249564 202816 249614 202872
rect 249614 202816 249628 202872
rect 249564 202812 249628 202816
rect 249380 196556 249444 196620
rect 236316 193352 236380 193356
rect 236316 193296 236330 193352
rect 236330 193296 236380 193352
rect 236316 193292 236380 193296
rect 249380 191762 249444 191826
rect 249196 182200 249260 182204
rect 249196 182144 249246 182200
rect 249246 182144 249260 182200
rect 249196 182140 249260 182144
rect 249196 180644 249260 180708
rect 249748 173844 249812 173908
rect 249380 164188 249444 164252
rect 249748 164188 249812 164252
rect 276060 157932 276124 157996
rect 395844 157932 395908 157996
rect 276060 157660 276124 157724
rect 249380 157388 249444 157452
rect 314700 157388 314764 157452
rect 395844 157524 395908 157588
rect 314700 157116 314764 157180
rect 285628 87484 285692 87548
rect 239996 87076 240060 87140
rect 251220 87212 251284 87276
rect 251220 87136 251284 87140
rect 285628 87212 285692 87276
rect 251220 87080 251234 87136
rect 251234 87080 251284 87136
rect 251220 87076 251284 87080
rect 405596 87212 405660 87276
rect 405596 86940 405660 87004
rect 481588 87348 481652 87412
rect 481588 87076 481652 87140
rect 395844 76468 395908 76532
rect 241284 76060 241348 76124
rect 395844 76060 395908 76124
rect 492628 76196 492692 76260
rect 285628 75788 285692 75852
rect 492628 75924 492692 75988
rect 285628 75516 285692 75580
rect 327028 63820 327092 63884
rect 280108 63684 280172 63748
rect 237236 63548 237300 63612
rect 280108 63412 280172 63476
rect 327028 63548 327092 63612
rect 405412 63956 405476 64020
rect 405596 63548 405660 63612
rect 233004 40156 233068 40220
rect 327028 40292 327092 40356
rect 327028 40020 327092 40084
rect 405596 40292 405660 40356
rect 405596 40020 405660 40084
rect 287100 29548 287164 29612
rect 249748 29412 249812 29476
rect 235764 29140 235828 29204
rect 287100 29140 287164 29204
rect 405596 29412 405660 29476
rect 481588 29412 481652 29476
rect 405596 29004 405660 29068
rect 481588 29140 481652 29204
rect 249748 28868 249812 28932
rect 465580 21932 465644 21996
rect 376708 17172 376772 17236
rect 249748 17036 249812 17100
rect 231716 16628 231780 16692
rect 249748 16764 249812 16828
rect 260972 16764 261036 16828
rect 260788 16628 260852 16692
rect 304764 16628 304828 16692
rect 304948 16492 305012 16556
rect 357388 16900 357452 16964
rect 376708 16960 376772 16964
rect 376708 16904 376722 16960
rect 376722 16904 376772 16960
rect 376708 16900 376772 16904
rect 396028 17036 396092 17100
rect 357388 16628 357452 16692
rect 396028 16628 396092 16692
rect 492628 16900 492692 16964
rect 492628 16628 492692 16692
rect 466500 11596 466564 11660
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 231715 579324 231781 579325
rect 231715 579260 231716 579324
rect 231780 579260 231781 579324
rect 231715 579259 231781 579260
rect 233003 579324 233069 579325
rect 233003 579260 233004 579324
rect 233068 579260 233069 579324
rect 233003 579259 233069 579260
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 16693 231778 579259
rect 233006 40221 233066 579259
rect 234804 560454 235404 595898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 235763 579324 235829 579325
rect 235763 579260 235764 579324
rect 235828 579260 235829 579324
rect 235763 579259 235829 579260
rect 237235 579324 237301 579325
rect 237235 579260 237236 579324
rect 237300 579260 237301 579324
rect 237235 579259 237301 579260
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 233003 40220 233069 40221
rect 233003 40156 233004 40220
rect 233068 40156 233069 40220
rect 233003 40155 233069 40156
rect 234804 20454 235404 55898
rect 235766 29205 235826 579259
rect 236315 270468 236381 270469
rect 236315 270404 236316 270468
rect 236380 270404 236381 270468
rect 236315 270403 236381 270404
rect 236318 260949 236378 270403
rect 236315 260948 236381 260949
rect 236315 260884 236316 260948
rect 236380 260884 236381 260948
rect 236315 260883 236381 260884
rect 236315 222052 236381 222053
rect 236315 221988 236316 222052
rect 236380 221988 236381 222052
rect 236315 221987 236381 221988
rect 236318 212669 236378 221987
rect 236315 212668 236381 212669
rect 236315 212604 236316 212668
rect 236380 212604 236381 212668
rect 236315 212603 236381 212604
rect 236315 202876 236381 202877
rect 236315 202812 236316 202876
rect 236380 202812 236381 202876
rect 236315 202811 236381 202812
rect 236318 193357 236378 202811
rect 236315 193356 236381 193357
rect 236315 193292 236316 193356
rect 236380 193292 236381 193356
rect 236315 193291 236381 193292
rect 237238 63613 237298 579259
rect 238404 564054 239004 599498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 239443 583132 239509 583133
rect 239443 583068 239444 583132
rect 239508 583068 239509 583132
rect 239443 583067 239509 583068
rect 239259 582996 239325 582997
rect 239259 582932 239260 582996
rect 239324 582932 239325 582996
rect 239259 582931 239325 582932
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238158 422058 238218 428622
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 239262 295221 239322 582931
rect 239446 338061 239506 583067
rect 239995 579324 240061 579325
rect 239995 579260 239996 579324
rect 240060 579260 240061 579324
rect 239995 579259 240061 579260
rect 241283 579324 241349 579325
rect 241283 579260 241284 579324
rect 241348 579260 241349 579324
rect 241283 579259 241349 579260
rect 239443 338060 239509 338061
rect 239443 337996 239444 338060
rect 239508 337996 239509 338060
rect 239443 337995 239509 337996
rect 239259 295220 239325 295221
rect 239259 295156 239260 295220
rect 239324 295156 239325 295220
rect 239259 295155 239325 295156
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 237235 63612 237301 63613
rect 237235 63548 237236 63612
rect 237300 63548 237301 63612
rect 237235 63547 237301 63548
rect 238404 60054 239004 95498
rect 239998 87141 240058 579259
rect 240918 442458 240978 451062
rect 241286 429538 241346 579259
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 240550 424690 240610 429302
rect 240550 424630 240978 424690
rect 240918 424010 240978 424630
rect 240918 423950 241346 424010
rect 241286 423330 241346 423950
rect 240918 423270 241346 423330
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 240550 421290 240610 421822
rect 240550 421230 240794 421290
rect 240734 407098 240794 421230
rect 240918 418570 240978 423270
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 240918 418510 241346 418570
rect 240918 394858 240978 403462
rect 240918 385338 240978 393942
rect 240918 375818 240978 382382
rect 240918 368338 240978 374902
rect 240918 356778 240978 364702
rect 240734 349298 240794 355862
rect 239995 87140 240061 87141
rect 239995 87076 239996 87140
rect 240060 87076 240061 87140
rect 239995 87075 240061 87076
rect 241286 76125 241346 418510
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 241283 76124 241349 76125
rect 241283 76060 241284 76124
rect 241348 76060 241349 76124
rect 241283 76059 241349 76060
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 235763 29204 235829 29205
rect 235763 29140 235764 29204
rect 235828 29140 235829 29204
rect 235763 29139 235829 29140
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 231715 16692 231781 16693
rect 231715 16628 231716 16692
rect 231780 16628 231781 16692
rect 231715 16627 231781 16628
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 249563 579324 249629 579325
rect 249563 579260 249564 579324
rect 249628 579260 249629 579324
rect 249563 579259 249629 579260
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 249566 457330 249626 579259
rect 249382 457270 249626 457330
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 249382 451978 249442 457270
rect 249566 433530 249626 442222
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 249566 433470 249846 433530
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 249566 404970 249626 406862
rect 249382 404910 249626 404970
rect 249382 403610 249442 404910
rect 249382 403550 249626 403610
rect 249566 403018 249626 403550
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 249566 385930 249626 386462
rect 249382 385870 249626 385930
rect 249382 382618 249442 385870
rect 249382 364938 249442 366742
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 249382 334253 249442 350422
rect 249379 334252 249445 334253
rect 249379 334188 249380 334252
rect 249444 334188 249445 334252
rect 249379 334187 249445 334188
rect 249379 328506 249445 328507
rect 249379 328442 249380 328506
rect 249444 328442 249445 328506
rect 249379 328441 249445 328442
rect 249382 322285 249442 328441
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 249379 322284 249445 322285
rect 249379 322220 249380 322284
rect 249444 322220 249445 322284
rect 249379 322219 249445 322220
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 249011 317524 249077 317525
rect 249011 317460 249012 317524
rect 249076 317460 249077 317524
rect 249011 317459 249077 317460
rect 249014 309229 249074 317459
rect 249011 309228 249077 309229
rect 249011 309164 249012 309228
rect 249076 309164 249077 309228
rect 249011 309163 249077 309164
rect 249195 308956 249261 308957
rect 249195 308892 249196 308956
rect 249260 308892 249261 308956
rect 249195 308891 249261 308892
rect 249198 302293 249258 308891
rect 249195 302292 249261 302293
rect 249195 302228 249196 302292
rect 249260 302228 249261 302292
rect 249195 302227 249261 302228
rect 249195 302156 249261 302157
rect 249195 302092 249196 302156
rect 249260 302092 249261 302156
rect 249195 302091 249261 302092
rect 249198 298077 249258 302091
rect 249195 298076 249261 298077
rect 249195 298012 249196 298076
rect 249260 298012 249261 298076
rect 249195 298011 249261 298012
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 249379 288556 249445 288557
rect 249379 288492 249380 288556
rect 249444 288492 249445 288556
rect 249379 288491 249445 288492
rect 249382 288421 249442 288491
rect 249379 288420 249445 288421
rect 249379 288356 249380 288420
rect 249444 288356 249445 288420
rect 249379 288355 249445 288356
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 249195 279036 249261 279037
rect 249195 278972 249196 279036
rect 249260 278972 249261 279036
rect 249195 278971 249261 278972
rect 249198 277405 249258 278971
rect 249195 277404 249261 277405
rect 249195 277340 249196 277404
rect 249260 277340 249261 277404
rect 249195 277339 249261 277340
rect 249379 267884 249445 267885
rect 249379 267820 249380 267884
rect 249444 267820 249445 267884
rect 249379 267819 249445 267820
rect 249382 263805 249442 267819
rect 249379 263804 249445 263805
rect 249379 263740 249380 263804
rect 249444 263740 249445 263804
rect 249379 263739 249445 263740
rect 249195 263532 249261 263533
rect 249195 263468 249196 263532
rect 249260 263468 249261 263532
rect 249195 263467 249261 263468
rect 249198 259538 249258 263467
rect 249566 253330 249626 259302
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 249382 253270 249626 253330
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 249382 241909 249442 253270
rect 249379 241908 249445 241909
rect 249379 241844 249380 241908
rect 249444 241844 249445 241908
rect 249379 241843 249445 241844
rect 249195 241772 249261 241773
rect 249195 241708 249196 241772
rect 249260 241708 249261 241772
rect 249195 241707 249261 241708
rect 249198 241501 249258 241707
rect 249195 241500 249261 241501
rect 249195 241436 249196 241500
rect 249260 241436 249261 241500
rect 249195 241435 249261 241436
rect 249379 240956 249445 240957
rect 249379 240892 249380 240956
rect 249444 240892 249445 240956
rect 249379 240891 249445 240892
rect 249382 225045 249442 240891
rect 249379 225044 249445 225045
rect 249379 224980 249380 225044
rect 249444 224980 249445 225044
rect 249379 224979 249445 224980
rect 249563 224772 249629 224773
rect 249563 224708 249564 224772
rect 249628 224708 249629 224772
rect 249563 224707 249629 224708
rect 249566 217429 249626 224707
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 249195 217428 249261 217429
rect 249195 217364 249196 217428
rect 249260 217364 249261 217428
rect 249195 217363 249261 217364
rect 249563 217428 249629 217429
rect 249563 217364 249564 217428
rect 249628 217364 249629 217428
rect 249563 217363 249629 217364
rect 249198 212533 249258 217363
rect 249195 212532 249261 212533
rect 249195 212468 249196 212532
rect 249260 212468 249261 212532
rect 249195 212467 249261 212468
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 249563 205460 249629 205461
rect 249563 205396 249564 205460
rect 249628 205396 249629 205460
rect 249563 205395 249629 205396
rect 249566 202877 249626 205395
rect 249563 202876 249629 202877
rect 249563 202812 249564 202876
rect 249628 202812 249629 202876
rect 249563 202811 249629 202812
rect 249379 196620 249445 196621
rect 249379 196556 249380 196620
rect 249444 196556 249445 196620
rect 249379 196555 249445 196556
rect 249382 191827 249442 196555
rect 249379 191826 249445 191827
rect 249379 191762 249380 191826
rect 249444 191762 249445 191826
rect 249379 191761 249445 191762
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 249195 182204 249261 182205
rect 249195 182140 249196 182204
rect 249260 182140 249261 182204
rect 249195 182139 249261 182140
rect 249198 180709 249258 182139
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 249195 180708 249261 180709
rect 249195 180644 249196 180708
rect 249260 180644 249261 180708
rect 249195 180643 249261 180644
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 249747 173908 249813 173909
rect 249747 173844 249748 173908
rect 249812 173844 249813 173908
rect 249747 173843 249813 173844
rect 249750 164253 249810 173843
rect 249379 164252 249445 164253
rect 249379 164188 249380 164252
rect 249444 164188 249445 164252
rect 249379 164187 249445 164188
rect 249747 164252 249813 164253
rect 249747 164188 249748 164252
rect 249812 164188 249813 164252
rect 249747 164187 249813 164188
rect 249382 157453 249442 164187
rect 249379 157452 249445 157453
rect 249379 157388 249380 157452
rect 249444 157388 249445 157452
rect 249379 157387 249445 157388
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 251219 87276 251285 87277
rect 251219 87212 251220 87276
rect 251284 87212 251285 87276
rect 251219 87211 251285 87212
rect 251222 87141 251282 87211
rect 251219 87140 251285 87141
rect 251219 87076 251220 87140
rect 251284 87076 251285 87140
rect 251219 87075 251285 87076
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 249747 29476 249813 29477
rect 249747 29412 249748 29476
rect 249812 29412 249813 29476
rect 249747 29411 249813 29412
rect 249750 28933 249810 29411
rect 249747 28932 249813 28933
rect 249747 28868 249748 28932
rect 249812 28868 249813 28932
rect 249747 28867 249813 28868
rect 249747 17100 249813 17101
rect 249747 17036 249748 17100
rect 249812 17036 249813 17100
rect 249747 17035 249813 17036
rect 249750 16829 249810 17035
rect 249747 16828 249813 16829
rect 249747 16764 249748 16828
rect 249812 16764 249813 16828
rect 249747 16763 249813 16764
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 260971 16828 261037 16829
rect 260971 16764 260972 16828
rect 261036 16764 261037 16828
rect 260971 16763 261037 16764
rect 260787 16692 260853 16693
rect 260787 16628 260788 16692
rect 260852 16690 260853 16692
rect 260974 16690 261034 16763
rect 260852 16630 261034 16690
rect 260852 16628 260853 16630
rect 260787 16627 260853 16628
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 276059 157996 276125 157997
rect 276059 157932 276060 157996
rect 276124 157932 276125 157996
rect 276059 157931 276125 157932
rect 276062 157725 276122 157931
rect 276059 157724 276125 157725
rect 276059 157660 276060 157724
rect 276124 157660 276125 157724
rect 276059 157659 276125 157660
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 285627 87548 285693 87549
rect 285627 87484 285628 87548
rect 285692 87484 285693 87548
rect 285627 87483 285693 87484
rect 285630 87277 285690 87483
rect 285627 87276 285693 87277
rect 285627 87212 285628 87276
rect 285692 87212 285693 87276
rect 285627 87211 285693 87212
rect 285627 75852 285693 75853
rect 285627 75788 285628 75852
rect 285692 75788 285693 75852
rect 285627 75787 285693 75788
rect 285630 75581 285690 75787
rect 285627 75580 285693 75581
rect 285627 75516 285628 75580
rect 285692 75516 285693 75580
rect 285627 75515 285693 75516
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 280107 63748 280173 63749
rect 280107 63684 280108 63748
rect 280172 63684 280173 63748
rect 280107 63683 280173 63684
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 280110 63477 280170 63683
rect 278004 63334 278604 63418
rect 280107 63476 280173 63477
rect 280107 63412 280108 63476
rect 280172 63412 280173 63476
rect 280107 63411 280173 63412
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 287099 29612 287165 29613
rect 287099 29548 287100 29612
rect 287164 29548 287165 29612
rect 287099 29547 287165 29548
rect 287102 29205 287162 29547
rect 287099 29204 287165 29205
rect 287099 29140 287100 29204
rect 287164 29140 287165 29204
rect 287099 29139 287165 29140
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 304763 16692 304829 16693
rect 304763 16628 304764 16692
rect 304828 16690 304829 16692
rect 304828 16630 305010 16690
rect 304828 16628 304829 16630
rect 304763 16627 304829 16628
rect 304950 16557 305010 16630
rect 304947 16556 305013 16557
rect 304947 16492 304948 16556
rect 305012 16492 305013 16556
rect 304947 16491 305013 16492
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 314699 157452 314765 157453
rect 314699 157388 314700 157452
rect 314764 157388 314765 157452
rect 314699 157387 314765 157388
rect 314702 157181 314762 157387
rect 314699 157180 314765 157181
rect 314699 157116 314700 157180
rect 314764 157116 314765 157180
rect 314699 157115 314765 157116
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 327027 63884 327093 63885
rect 327027 63820 327028 63884
rect 327092 63820 327093 63884
rect 327027 63819 327093 63820
rect 327030 63613 327090 63819
rect 327027 63612 327093 63613
rect 327027 63548 327028 63612
rect 327092 63548 327093 63612
rect 327027 63547 327093 63548
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 327027 40356 327093 40357
rect 327027 40292 327028 40356
rect 327092 40292 327093 40356
rect 327027 40291 327093 40292
rect 327030 40085 327090 40291
rect 327027 40084 327093 40085
rect 327027 40020 327028 40084
rect 327092 40020 327093 40084
rect 327027 40019 327093 40020
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 341379 299436 341445 299437
rect 341379 299372 341380 299436
rect 341444 299372 341445 299436
rect 341379 299371 341445 299372
rect 341382 289917 341442 299371
rect 341379 289916 341445 289917
rect 341379 289852 341380 289916
rect 341444 289852 341445 289916
rect 341379 289851 341445 289852
rect 341379 280124 341445 280125
rect 341379 280060 341380 280124
rect 341444 280060 341445 280124
rect 341379 280059 341445 280060
rect 336963 274004 337029 274005
rect 336963 273940 336964 274004
rect 337028 273940 337029 274004
rect 336963 273939 337029 273940
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 336966 260677 337026 273939
rect 341382 270605 341442 280059
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 341379 270604 341445 270605
rect 341379 270540 341380 270604
rect 341444 270540 341445 270604
rect 341379 270539 341445 270540
rect 341379 260812 341445 260813
rect 341379 260748 341380 260812
rect 341444 260748 341445 260812
rect 341379 260747 341445 260748
rect 336963 260676 337029 260677
rect 336963 260612 336964 260676
rect 337028 260612 337029 260676
rect 336963 260611 337029 260612
rect 341382 251293 341442 260747
rect 341379 251292 341445 251293
rect 341379 251228 341380 251292
rect 341444 251228 341445 251292
rect 341379 251227 341445 251228
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 358859 220828 358925 220829
rect 358859 220764 358860 220828
rect 358924 220764 358925 220828
rect 358859 220763 358925 220764
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 358862 211173 358922 220763
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 358859 211172 358925 211173
rect 358859 211108 358860 211172
rect 358924 211108 358925 211172
rect 358859 211107 358925 211108
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 357387 16964 357453 16965
rect 357387 16900 357388 16964
rect 357452 16900 357453 16964
rect 357387 16899 357453 16900
rect 357390 16693 357450 16899
rect 357387 16692 357453 16693
rect 357387 16628 357388 16692
rect 357452 16628 357453 16692
rect 357387 16627 357453 16628
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 366955 222188 367021 222189
rect 366955 222124 366956 222188
rect 367020 222124 367021 222188
rect 366955 222123 367021 222124
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 366958 212669 367018 222123
rect 366955 212668 367021 212669
rect 366955 212604 366956 212668
rect 367020 212604 367021 212668
rect 366955 212603 367021 212604
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 376707 17236 376773 17237
rect 376707 17172 376708 17236
rect 376772 17172 376773 17236
rect 376707 17171 376773 17172
rect 376710 16965 376770 17171
rect 376707 16964 376773 16965
rect 376707 16900 376708 16964
rect 376772 16900 376773 16964
rect 376707 16899 376773 16900
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 395843 157996 395909 157997
rect 395843 157932 395844 157996
rect 395908 157932 395909 157996
rect 395843 157931 395909 157932
rect 395846 157589 395906 157931
rect 395843 157588 395909 157589
rect 395843 157524 395844 157588
rect 395908 157524 395909 157588
rect 395843 157523 395909 157524
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 395843 76532 395909 76533
rect 395843 76468 395844 76532
rect 395908 76468 395909 76532
rect 395843 76467 395909 76468
rect 395846 76125 395906 76467
rect 395843 76124 395909 76125
rect 395843 76060 395844 76124
rect 395908 76060 395909 76124
rect 395843 76059 395909 76060
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396027 17100 396093 17101
rect 396027 17036 396028 17100
rect 396092 17036 396093 17100
rect 396027 17035 396093 17036
rect 396030 16693 396090 17035
rect 396027 16692 396093 16693
rect 396027 16628 396028 16692
rect 396092 16628 396093 16692
rect 396027 16627 396093 16628
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 405595 87276 405661 87277
rect 405595 87212 405596 87276
rect 405660 87212 405661 87276
rect 405595 87211 405661 87212
rect 405598 87005 405658 87211
rect 405595 87004 405661 87005
rect 405595 86940 405596 87004
rect 405660 86940 405661 87004
rect 405595 86939 405661 86940
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 405411 64020 405477 64021
rect 405411 63956 405412 64020
rect 405476 63956 405477 64020
rect 405411 63955 405477 63956
rect 405414 63610 405474 63955
rect 405595 63612 405661 63613
rect 405595 63610 405596 63612
rect 405414 63550 405596 63610
rect 405595 63548 405596 63550
rect 405660 63548 405661 63612
rect 405595 63547 405661 63548
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 405595 40356 405661 40357
rect 405595 40292 405596 40356
rect 405660 40292 405661 40356
rect 405595 40291 405661 40292
rect 405598 40085 405658 40291
rect 405595 40084 405661 40085
rect 405595 40020 405596 40084
rect 405660 40020 405661 40084
rect 405595 40019 405661 40020
rect 405595 29476 405661 29477
rect 405595 29412 405596 29476
rect 405660 29412 405661 29476
rect 405595 29411 405661 29412
rect 405598 29069 405658 29411
rect 405595 29068 405661 29069
rect 405595 29004 405596 29068
rect 405660 29004 405661 29068
rect 405595 29003 405661 29004
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 465947 583404 466013 583405
rect 465947 583340 465948 583404
rect 466012 583340 466013 583404
rect 465947 583339 466013 583340
rect 465763 583268 465829 583269
rect 465763 583204 465764 583268
rect 465828 583204 465829 583268
rect 465763 583203 465829 583204
rect 465579 579732 465645 579733
rect 465579 579668 465580 579732
rect 465644 579668 465645 579732
rect 465579 579667 465645 579668
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 465582 21997 465642 579667
rect 465766 486165 465826 583203
rect 465950 533085 466010 583339
rect 466499 579324 466565 579325
rect 466499 579260 466500 579324
rect 466564 579260 466565 579324
rect 466499 579259 466565 579260
rect 465947 533084 466013 533085
rect 465947 533020 465948 533084
rect 466012 533020 466013 533084
rect 465947 533019 466013 533020
rect 465763 486164 465829 486165
rect 465763 486100 465764 486164
rect 465828 486100 465829 486164
rect 465763 486099 465829 486100
rect 465579 21996 465645 21997
rect 465579 21932 465580 21996
rect 465644 21932 465645 21996
rect 465579 21931 465645 21932
rect 466502 11661 466562 579259
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 466499 11660 466565 11661
rect 466499 11596 466500 11660
rect 466564 11596 466565 11660
rect 466499 11595 466565 11596
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 481587 87412 481653 87413
rect 481587 87348 481588 87412
rect 481652 87348 481653 87412
rect 481587 87347 481653 87348
rect 481590 87141 481650 87347
rect 481587 87140 481653 87141
rect 481587 87076 481588 87140
rect 481652 87076 481653 87140
rect 481587 87075 481653 87076
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 481587 29476 481653 29477
rect 481587 29412 481588 29476
rect 481652 29412 481653 29476
rect 481587 29411 481653 29412
rect 481590 29205 481650 29411
rect 481587 29204 481653 29205
rect 481587 29140 481588 29204
rect 481652 29140 481653 29204
rect 481587 29139 481653 29140
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 492627 76260 492693 76261
rect 492627 76196 492628 76260
rect 492692 76196 492693 76260
rect 492627 76195 492693 76196
rect 492630 75989 492690 76195
rect 492627 75988 492693 75989
rect 492627 75924 492628 75988
rect 492692 75924 492693 75988
rect 492627 75923 492693 75924
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 492627 16964 492693 16965
rect 492627 16900 492628 16964
rect 492692 16900 492693 16964
rect 492627 16899 492693 16900
rect 492630 16693 492690 16899
rect 492627 16692 492693 16693
rect 492627 16628 492628 16692
rect 492692 16628 492693 16692
rect 492627 16627 492693 16628
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238070 428622 238306 428858
rect 238070 421822 238306 422058
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 240830 451062 241066 451298
rect 240830 442222 241066 442458
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 240462 429302 240698 429538
rect 241198 429302 241434 429538
rect 242186 423418 242422 423654
rect 240462 421822 240698 422058
rect 242186 423098 242422 423334
rect 240646 406862 240882 407098
rect 240830 403462 241066 403698
rect 240830 394622 241066 394858
rect 240830 393942 241066 394178
rect 240830 385102 241066 385338
rect 240830 382382 241066 382618
rect 240830 375582 241066 375818
rect 240830 374902 241066 375138
rect 240830 368102 241066 368338
rect 240830 364702 241066 364938
rect 240830 356542 241066 356778
rect 240646 355862 240882 356098
rect 240646 349062 240882 349298
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 249294 451742 249530 451978
rect 249478 442222 249714 442458
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 249846 433382 250082 433618
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 249478 406862 249714 407098
rect 249478 402782 249714 403018
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 249478 386462 249714 386698
rect 249294 382382 249530 382618
rect 249294 366742 249530 366978
rect 249294 364702 249530 364938
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 249294 350422 249530 350658
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 249110 259302 249346 259538
rect 249478 259302 249714 259538
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 353786 211018 354022 211254
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451978 270986 452134
rect 235222 451898 249294 451978
rect -2916 451876 249294 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 249068 451742 249294 451876
rect 249530 451898 270986 451978
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect 249530 451876 586840 451898
rect 249530 451742 249572 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect 249068 451700 249572 451742
rect 249068 451340 249388 451700
rect 240788 451298 249388 451340
rect 240788 451062 240830 451298
rect 241066 451062 249388 451298
rect 240788 451020 249388 451062
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect 240788 442458 249756 442500
rect 240788 442222 240830 442458
rect 241066 442222 249478 442458
rect 249714 442222 249756 442458
rect 240788 442180 249756 442222
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect 249804 433618 250124 433660
rect 249804 433382 249846 433618
rect 250082 433382 250124 433618
rect 240420 429538 241476 429580
rect 240420 429302 240462 429538
rect 240698 429302 241198 429538
rect 241434 429302 241476 429538
rect 240420 429260 241476 429302
rect 249804 428900 250124 433382
rect 238028 428858 250124 428900
rect 238028 428622 238070 428858
rect 238306 428622 250124 428858
rect 238028 428580 250124 428622
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect 238028 422058 240740 422100
rect 238028 421822 238070 422058
rect 238306 421822 240462 422058
rect 240698 421822 240740 422058
rect 238028 421780 240740 421822
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect 240604 407098 249756 407140
rect 240604 406862 240646 407098
rect 240882 406862 249478 407098
rect 249714 406862 249756 407098
rect 240604 406820 249756 406862
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect 240788 403698 247548 403740
rect 240788 403462 240830 403698
rect 241066 403462 247548 403698
rect 240788 403420 247548 403462
rect 247228 403060 247548 403420
rect 247228 403018 249756 403060
rect 247228 402782 249478 403018
rect 249714 402782 249756 403018
rect 247228 402740 249756 402782
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect 240788 394858 245524 394900
rect 240788 394622 240830 394858
rect 241066 394622 245524 394858
rect 240788 394580 245524 394622
rect 245204 394220 245524 394580
rect 240788 394178 245524 394220
rect 240788 393942 240830 394178
rect 241066 393942 245524 394178
rect 240788 393900 245524 393942
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect 249436 386698 249756 386740
rect 249436 386462 249478 386698
rect 249714 386462 249756 386698
rect 249436 385380 249756 386462
rect 240788 385338 249756 385380
rect 240788 385102 240830 385338
rect 241066 385102 249756 385338
rect 240788 385060 249756 385102
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect 240788 382618 249572 382660
rect 240788 382382 240830 382618
rect 241066 382382 249294 382618
rect 249530 382382 249572 382618
rect 240788 382340 249572 382382
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect 240788 375818 241660 375860
rect 240788 375582 240830 375818
rect 241066 375582 241660 375818
rect 240788 375540 241660 375582
rect 241340 375180 241660 375540
rect 240788 375138 241660 375180
rect 240788 374902 240830 375138
rect 241066 374902 241660 375138
rect 240788 374860 241660 374902
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect 240788 368338 249572 368380
rect 240788 368102 240830 368338
rect 241066 368102 249572 368338
rect 240788 368060 249572 368102
rect 249252 366978 249572 368060
rect 249252 366742 249294 366978
rect 249530 366742 249572 366978
rect 249252 366700 249572 366742
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect 240788 364938 249572 364980
rect 240788 364702 240830 364938
rect 241066 364702 249294 364938
rect 249530 364702 249572 364938
rect 240788 364660 249572 364702
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect 240788 356778 244420 356820
rect 240788 356542 240830 356778
rect 241066 356542 244420 356778
rect 240788 356500 244420 356542
rect 244100 356140 244420 356500
rect 240604 356098 244420 356140
rect 240604 355862 240646 356098
rect 240882 355862 244420 356098
rect 240604 355820 244420 355862
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect 249252 350658 249940 350700
rect 249252 350422 249294 350658
rect 249530 350422 249940 350658
rect 249252 350380 249940 350422
rect 249620 349340 249940 350380
rect 240604 349298 249940 349340
rect 240604 349062 240646 349298
rect 240882 349062 249940 349298
rect 240604 349020 249940 349062
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect 249068 259538 249756 259580
rect 249068 259302 249110 259538
rect 249346 259302 249478 259538
rect 249714 259302 249756 259538
rect 249068 259260 249756 259302
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1608061857
transform 1 0 230000 0 1 340000
box 0 0 239540 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
