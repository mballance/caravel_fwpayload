VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 3700.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3203.520 2700.000 3204.120 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 346.470 3697.600 346.750 3700.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 269.650 3697.600 269.930 3700.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3336.120 2700.000 3336.720 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2691.550 0.000 2691.830 2.400 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3402.080 2700.000 3402.680 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 192.370 3697.600 192.650 3700.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3468.040 2700.000 3468.640 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 2.400 486.840 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 2.400 421.560 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 2.400 356.960 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 501.030 3697.600 501.310 3700.000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 2.400 291.680 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 2.400 227.080 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3534.000 2700.000 3534.600 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 3697.600 115.370 3700.000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2697.070 0.000 2697.350 2.400 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 2.400 161.800 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 2.400 97.200 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 3697.600 38.550 3700.000 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 2.400 32.600 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3599.960 2700.000 3600.560 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 2.400 681.320 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3665.920 2700.000 3666.520 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 2.400 616.720 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 423.750 3697.600 424.030 3700.000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2674.990 0.000 2675.270 2.400 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2680.510 0.000 2680.790 2.400 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3269.480 2700.000 3270.080 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 2.400 551.440 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2686.030 0.000 2686.310 2.400 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 32.680 2700.000 33.280 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2146.800 2700.000 2147.400 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2344.680 2700.000 2345.280 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2543.240 2700.000 2543.840 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2741.120 2700.000 2741.720 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3005.640 2700.000 3006.240 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.190 3697.600 2661.470 3700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2352.530 3697.600 2352.810 3700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2121.150 3697.600 2121.430 3700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1889.770 3697.600 1890.050 3700.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1658.390 3697.600 1658.670 3700.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 230.560 2700.000 231.160 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1426.550 3697.600 1426.830 3700.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 3697.600 1195.450 3700.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 963.790 3697.600 964.070 3700.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 732.410 3697.600 732.690 3700.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3666.600 2.400 3667.200 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3342.240 2.400 3342.840 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3147.080 2.400 3147.680 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2952.600 2.400 2953.200 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2758.120 2.400 2758.720 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2562.960 2.400 2563.560 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 428.440 2700.000 429.040 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2368.480 2.400 2369.080 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2174.000 2.400 2174.600 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1848.960 2.400 1849.560 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1654.480 2.400 1655.080 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1460.000 2.400 1460.600 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 2.400 1265.440 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1070.360 2.400 1070.960 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.200 2.400 875.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 627.000 2700.000 627.600 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 824.880 2700.000 825.480 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1023.440 2700.000 1024.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1221.320 2700.000 1221.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1551.800 2700.000 1552.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1750.360 2700.000 1750.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1948.240 2700.000 1948.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 164.600 2700.000 165.200 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2278.720 2700.000 2279.320 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2476.600 2700.000 2477.200 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2675.160 2700.000 2675.760 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2873.040 2700.000 2873.640 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3137.560 2700.000 3138.160 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2506.630 3697.600 2506.910 3700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2198.430 3697.600 2198.710 3700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1966.590 3697.600 1966.870 3700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1735.210 3697.600 1735.490 3700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1503.830 3697.600 1504.110 3700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 362.480 2700.000 363.080 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1272.450 3697.600 1272.730 3700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1041.070 3697.600 1041.350 3700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 809.690 3697.600 809.970 3700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 578.310 3697.600 578.590 3700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3536.720 2.400 3537.320 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3212.360 2.400 3212.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3017.200 2.400 3017.800 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2822.720 2.400 2823.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2628.240 2.400 2628.840 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2433.080 2.400 2433.680 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 561.040 2700.000 561.640 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2238.600 2.400 2239.200 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2044.120 2.400 2044.720 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1719.080 2.400 1719.680 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1524.600 2.400 1525.200 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1330.120 2.400 1330.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 2.400 1135.560 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 940.480 2.400 941.080 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.000 2.400 746.600 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 758.920 2700.000 759.520 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 957.480 2700.000 958.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1155.360 2700.000 1155.960 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1353.920 2700.000 1354.520 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1684.400 2700.000 1685.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1882.280 2700.000 1882.880 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2080.160 2700.000 2080.760 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 98.640 2700.000 99.240 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2212.760 2700.000 2213.360 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2410.640 2700.000 2411.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2609.200 2700.000 2609.800 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2807.080 2700.000 2807.680 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3071.600 2700.000 3072.200 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.910 3697.600 2584.190 3700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2275.250 3697.600 2275.530 3700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2043.870 3697.600 2044.150 3700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1812.490 3697.600 1812.770 3700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1581.110 3697.600 1581.390 3700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 296.520 2700.000 297.120 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1349.730 3697.600 1350.010 3700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1118.350 3697.600 1118.630 3700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.510 3697.600 886.790 3700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 655.130 3697.600 655.410 3700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3602.000 2.400 3602.600 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3276.960 2.400 3277.560 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3082.480 2.400 3083.080 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2888.000 2.400 2888.600 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2692.840 2.400 2693.440 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2498.360 2.400 2498.960 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 495.080 2700.000 495.680 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2303.200 2.400 2303.800 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2108.720 2.400 2109.320 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1784.360 2.400 1784.960 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1589.200 2.400 1589.800 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.720 2.400 1395.320 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 2.400 1200.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.080 2.400 1005.680 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 2.400 811.200 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 692.960 2700.000 693.560 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 891.520 2700.000 892.120 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1089.400 2700.000 1090.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1287.960 2700.000 1288.560 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1617.760 2700.000 1618.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1816.320 2700.000 1816.920 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2014.200 2700.000 2014.800 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2212.230 0.000 2212.510 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2228.790 0.000 2229.070 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2244.890 0.000 2245.170 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2261.450 0.000 2261.730 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2277.550 0.000 2277.830 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2294.110 0.000 2294.390 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.210 0.000 2310.490 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2326.770 0.000 2327.050 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2342.870 0.000 2343.150 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2359.430 0.000 2359.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.530 0.000 2375.810 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2392.090 0.000 2392.370 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2408.190 0.000 2408.470 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2424.750 0.000 2425.030 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2440.850 0.000 2441.130 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2457.410 0.000 2457.690 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.510 0.000 2473.790 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2490.070 0.000 2490.350 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.170 0.000 2506.450 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2522.730 0.000 2523.010 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2538.830 0.000 2539.110 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2555.390 0.000 2555.670 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.490 0.000 2571.770 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2588.050 0.000 2588.330 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2604.150 0.000 2604.430 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2620.710 0.000 2620.990 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2636.810 0.000 2637.090 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2653.370 0.000 2653.650 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 791.750 0.000 792.030 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.070 0.000 857.350 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 905.830 0.000 906.110 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.390 0.000 922.670 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.150 0.000 971.430 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.810 0.000 1004.090 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.470 0.000 1036.750 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1085.690 0.000 1085.970 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1101.790 0.000 1102.070 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1118.350 0.000 1118.630 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1151.010 0.000 1151.290 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1167.110 0.000 1167.390 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1199.770 0.000 1200.050 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1216.330 0.000 1216.610 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1232.430 0.000 1232.710 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1248.990 0.000 1249.270 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1265.090 0.000 1265.370 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1297.750 0.000 1298.030 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1314.310 0.000 1314.590 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1330.410 0.000 1330.690 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.970 0.000 1347.250 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1363.070 0.000 1363.350 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1379.630 0.000 1379.910 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.290 0.000 1412.570 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1428.390 0.000 1428.670 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.950 0.000 1445.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1461.050 0.000 1461.330 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1477.610 0.000 1477.890 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1493.710 0.000 1493.990 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.930 0.000 1543.210 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1559.030 0.000 1559.310 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1575.590 0.000 1575.870 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1591.690 0.000 1591.970 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.250 0.000 1608.530 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1624.350 0.000 1624.630 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1640.910 0.000 1641.190 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1657.010 0.000 1657.290 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1673.570 0.000 1673.850 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1689.670 0.000 1689.950 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1706.230 0.000 1706.510 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1722.330 0.000 1722.610 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1738.890 0.000 1739.170 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1771.550 0.000 1771.830 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1787.650 0.000 1787.930 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.210 0.000 1804.490 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1820.310 0.000 1820.590 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1836.870 0.000 1837.150 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1852.970 0.000 1853.250 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1869.530 0.000 1869.810 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1885.630 0.000 1885.910 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1902.190 0.000 1902.470 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1918.290 0.000 1918.570 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1934.850 0.000 1935.130 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1950.950 0.000 1951.230 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1967.510 0.000 1967.790 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.610 0.000 1983.890 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.170 0.000 2000.450 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2016.270 0.000 2016.550 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2032.830 0.000 2033.110 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.870 0.000 710.150 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2048.930 0.000 2049.210 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2065.490 0.000 2065.770 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2081.590 0.000 2081.870 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2098.150 0.000 2098.430 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2114.250 0.000 2114.530 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2130.810 0.000 2131.090 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2146.910 0.000 2147.190 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2163.470 0.000 2163.750 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2179.570 0.000 2179.850 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.130 0.000 2196.410 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2217.750 0.000 2218.030 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2234.310 0.000 2234.590 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2250.410 0.000 2250.690 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2266.970 0.000 2267.250 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2283.070 0.000 2283.350 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2299.630 0.000 2299.910 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2315.730 0.000 2316.010 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2332.290 0.000 2332.570 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2348.390 0.000 2348.670 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2364.950 0.000 2365.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2381.050 0.000 2381.330 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2397.610 0.000 2397.890 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2413.710 0.000 2413.990 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2430.270 0.000 2430.550 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2446.370 0.000 2446.650 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2462.930 0.000 2463.210 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2479.030 0.000 2479.310 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2495.590 0.000 2495.870 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2511.690 0.000 2511.970 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2528.250 0.000 2528.530 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2544.350 0.000 2544.630 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2560.910 0.000 2561.190 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2577.010 0.000 2577.290 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2593.570 0.000 2593.850 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2609.670 0.000 2609.950 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2626.230 0.000 2626.510 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2642.330 0.000 2642.610 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2658.890 0.000 2659.170 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 780.710 0.000 780.990 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.370 0.000 813.650 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 862.130 0.000 862.410 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 911.350 0.000 911.630 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1025.430 0.000 1025.710 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1041.990 0.000 1042.270 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1074.650 0.000 1074.930 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1107.310 0.000 1107.590 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1123.410 0.000 1123.690 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1172.630 0.000 1172.910 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1188.730 0.000 1189.010 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1205.290 0.000 1205.570 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1221.390 0.000 1221.670 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1237.950 0.000 1238.230 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1254.050 0.000 1254.330 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1270.610 0.000 1270.890 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1286.710 0.000 1286.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1303.270 0.000 1303.550 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1319.370 0.000 1319.650 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1401.250 0.000 1401.530 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1417.810 0.000 1418.090 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1433.910 0.000 1434.190 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1450.470 0.000 1450.750 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1466.570 0.000 1466.850 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1483.130 0.000 1483.410 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1499.230 0.000 1499.510 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1515.790 0.000 1516.070 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1531.890 0.000 1532.170 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.450 0.000 1548.730 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1564.550 0.000 1564.830 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1581.110 0.000 1581.390 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1597.210 0.000 1597.490 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1613.770 0.000 1614.050 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1629.870 0.000 1630.150 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1646.430 0.000 1646.710 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.530 0.000 1662.810 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1679.090 0.000 1679.370 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1695.190 0.000 1695.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1711.750 0.000 1712.030 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.850 0.000 1728.130 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1744.410 0.000 1744.690 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1760.510 0.000 1760.790 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1777.070 0.000 1777.350 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1793.170 0.000 1793.450 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1809.730 0.000 1810.010 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1825.830 0.000 1826.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1842.390 0.000 1842.670 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1858.490 0.000 1858.770 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1875.050 0.000 1875.330 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1891.150 0.000 1891.430 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1907.710 0.000 1907.990 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.810 0.000 1924.090 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1940.370 0.000 1940.650 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1956.470 0.000 1956.750 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1973.030 0.000 1973.310 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1989.130 0.000 1989.410 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2005.690 0.000 2005.970 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2021.790 0.000 2022.070 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2038.350 0.000 2038.630 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2054.450 0.000 2054.730 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2071.010 0.000 2071.290 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2087.110 0.000 2087.390 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2103.670 0.000 2103.950 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.770 0.000 2120.050 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2136.330 0.000 2136.610 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2152.430 0.000 2152.710 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2168.990 0.000 2169.270 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2185.090 0.000 2185.370 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2201.650 0.000 2201.930 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2223.270 0.000 2223.550 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2239.830 0.000 2240.110 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2255.930 0.000 2256.210 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2272.490 0.000 2272.770 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2288.590 0.000 2288.870 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2305.150 0.000 2305.430 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2321.250 0.000 2321.530 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2337.810 0.000 2338.090 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2353.910 0.000 2354.190 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2370.470 0.000 2370.750 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2386.570 0.000 2386.850 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2403.130 0.000 2403.410 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2419.230 0.000 2419.510 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2435.790 0.000 2436.070 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2451.890 0.000 2452.170 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2468.450 0.000 2468.730 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2484.550 0.000 2484.830 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2501.110 0.000 2501.390 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.210 0.000 2517.490 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2533.770 0.000 2534.050 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2549.870 0.000 2550.150 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2566.430 0.000 2566.710 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2582.530 0.000 2582.810 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2599.090 0.000 2599.370 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2615.190 0.000 2615.470 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.750 0.000 2632.030 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2647.850 0.000 2648.130 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2664.410 0.000 2664.690 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 818.890 0.000 819.170 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.550 0.000 851.830 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.310 0.000 900.590 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 916.870 0.000 917.150 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.970 0.000 933.250 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.530 0.000 949.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.850 0.000 1015.130 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1047.510 0.000 1047.790 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.610 0.000 1063.890 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.170 0.000 1080.450 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.270 0.000 1096.550 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1112.830 0.000 1113.110 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.490 0.000 1145.770 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.590 0.000 1161.870 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1226.910 0.000 1227.190 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.470 0.000 1243.750 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.570 0.000 1259.850 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1276.130 0.000 1276.410 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1292.230 0.000 1292.510 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1308.790 0.000 1309.070 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1324.890 0.000 1325.170 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.450 0.000 1341.730 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1390.210 0.000 1390.490 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1406.770 0.000 1407.050 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1472.090 0.000 1472.370 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1488.190 0.000 1488.470 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1504.750 0.000 1505.030 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1520.850 0.000 1521.130 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1537.410 0.000 1537.690 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1553.510 0.000 1553.790 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1570.070 0.000 1570.350 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1586.170 0.000 1586.450 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1602.730 0.000 1603.010 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1618.830 0.000 1619.110 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1635.390 0.000 1635.670 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1651.490 0.000 1651.770 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1668.050 0.000 1668.330 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1684.150 0.000 1684.430 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1700.710 0.000 1700.990 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1716.810 0.000 1717.090 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.370 0.000 1733.650 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1749.470 0.000 1749.750 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1766.030 0.000 1766.310 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1782.130 0.000 1782.410 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1798.690 0.000 1798.970 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1814.790 0.000 1815.070 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1831.350 0.000 1831.630 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1847.450 0.000 1847.730 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1864.010 0.000 1864.290 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1880.110 0.000 1880.390 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1896.670 0.000 1896.950 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1912.770 0.000 1913.050 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.330 0.000 1929.610 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1945.430 0.000 1945.710 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1961.990 0.000 1962.270 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1978.090 0.000 1978.370 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1994.650 0.000 1994.930 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2010.750 0.000 2011.030 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2027.310 0.000 2027.590 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2043.870 0.000 2044.150 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2059.970 0.000 2060.250 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2076.530 0.000 2076.810 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2092.630 0.000 2092.910 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2109.190 0.000 2109.470 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.290 0.000 2125.570 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2141.850 0.000 2142.130 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2157.950 0.000 2158.230 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2174.510 0.000 2174.790 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2190.610 0.000 2190.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2207.170 0.000 2207.450 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2669.470 0.000 2669.750 2.400 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2939.680 2700.000 2940.280 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3472.120 2.400 3472.720 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1485.840 2700.000 1486.440 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1978.840 2.400 1979.440 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2429.810 3697.600 2430.090 3700.000 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3406.840 2.400 3407.440 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1419.880 2700.000 1420.480 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1914.240 2.400 1914.840 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 2.400 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2694.220 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 2694.220 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2694.220 3688.405 ;
      LAYER met1 ;
        RECT 2.370 2.420 2694.220 3688.560 ;
      LAYER met2 ;
        RECT 2.400 3697.320 37.990 3698.250 ;
        RECT 38.830 3697.320 114.810 3698.250 ;
        RECT 115.650 3697.320 192.090 3698.250 ;
        RECT 192.930 3697.320 269.370 3698.250 ;
        RECT 270.210 3697.320 346.190 3698.250 ;
        RECT 347.030 3697.320 423.470 3698.250 ;
        RECT 424.310 3697.320 500.750 3698.250 ;
        RECT 501.590 3697.320 578.030 3698.250 ;
        RECT 578.870 3697.320 654.850 3698.250 ;
        RECT 655.690 3697.320 732.130 3698.250 ;
        RECT 732.970 3697.320 809.410 3698.250 ;
        RECT 810.250 3697.320 886.230 3698.250 ;
        RECT 887.070 3697.320 963.510 3698.250 ;
        RECT 964.350 3697.320 1040.790 3698.250 ;
        RECT 1041.630 3697.320 1118.070 3698.250 ;
        RECT 1118.910 3697.320 1194.890 3698.250 ;
        RECT 1195.730 3697.320 1272.170 3698.250 ;
        RECT 1273.010 3697.320 1349.450 3698.250 ;
        RECT 1350.290 3697.320 1426.270 3698.250 ;
        RECT 1427.110 3697.320 1503.550 3698.250 ;
        RECT 1504.390 3697.320 1580.830 3698.250 ;
        RECT 1581.670 3697.320 1658.110 3698.250 ;
        RECT 1658.950 3697.320 1734.930 3698.250 ;
        RECT 1735.770 3697.320 1812.210 3698.250 ;
        RECT 1813.050 3697.320 1889.490 3698.250 ;
        RECT 1890.330 3697.320 1966.310 3698.250 ;
        RECT 1967.150 3697.320 2043.590 3698.250 ;
        RECT 2044.430 3697.320 2120.870 3698.250 ;
        RECT 2121.710 3697.320 2198.150 3698.250 ;
        RECT 2198.990 3697.320 2274.970 3698.250 ;
        RECT 2275.810 3697.320 2352.250 3698.250 ;
        RECT 2353.090 3697.320 2429.530 3698.250 ;
        RECT 2430.370 3697.320 2506.350 3698.250 ;
        RECT 2507.190 3697.320 2583.630 3698.250 ;
        RECT 2584.470 3697.320 2660.910 3698.250 ;
        RECT 2661.750 3697.320 2689.070 3698.250 ;
        RECT 2.400 2.680 2689.070 3697.320 ;
        RECT 2.950 2.390 7.170 2.680 ;
        RECT 8.010 2.390 12.690 2.680 ;
        RECT 13.530 2.390 18.210 2.680 ;
        RECT 19.050 2.390 23.730 2.680 ;
        RECT 24.570 2.390 29.250 2.680 ;
        RECT 30.090 2.390 34.770 2.680 ;
        RECT 35.610 2.390 39.830 2.680 ;
        RECT 40.670 2.390 45.350 2.680 ;
        RECT 46.190 2.390 50.870 2.680 ;
        RECT 51.710 2.390 56.390 2.680 ;
        RECT 57.230 2.390 61.910 2.680 ;
        RECT 62.750 2.390 67.430 2.680 ;
        RECT 68.270 2.390 72.490 2.680 ;
        RECT 73.330 2.390 78.010 2.680 ;
        RECT 78.850 2.390 83.530 2.680 ;
        RECT 84.370 2.390 89.050 2.680 ;
        RECT 89.890 2.390 94.570 2.680 ;
        RECT 95.410 2.390 100.090 2.680 ;
        RECT 100.930 2.390 105.150 2.680 ;
        RECT 105.990 2.390 110.670 2.680 ;
        RECT 111.510 2.390 116.190 2.680 ;
        RECT 117.030 2.390 121.710 2.680 ;
        RECT 122.550 2.390 127.230 2.680 ;
        RECT 128.070 2.390 132.750 2.680 ;
        RECT 133.590 2.390 137.810 2.680 ;
        RECT 138.650 2.390 143.330 2.680 ;
        RECT 144.170 2.390 148.850 2.680 ;
        RECT 149.690 2.390 154.370 2.680 ;
        RECT 155.210 2.390 159.890 2.680 ;
        RECT 160.730 2.390 165.410 2.680 ;
        RECT 166.250 2.390 170.470 2.680 ;
        RECT 171.310 2.390 175.990 2.680 ;
        RECT 176.830 2.390 181.510 2.680 ;
        RECT 182.350 2.390 187.030 2.680 ;
        RECT 187.870 2.390 192.550 2.680 ;
        RECT 193.390 2.390 198.070 2.680 ;
        RECT 198.910 2.390 203.130 2.680 ;
        RECT 203.970 2.390 208.650 2.680 ;
        RECT 209.490 2.390 214.170 2.680 ;
        RECT 215.010 2.390 219.690 2.680 ;
        RECT 220.530 2.390 225.210 2.680 ;
        RECT 226.050 2.390 230.730 2.680 ;
        RECT 231.570 2.390 235.790 2.680 ;
        RECT 236.630 2.390 241.310 2.680 ;
        RECT 242.150 2.390 246.830 2.680 ;
        RECT 247.670 2.390 252.350 2.680 ;
        RECT 253.190 2.390 257.870 2.680 ;
        RECT 258.710 2.390 263.390 2.680 ;
        RECT 264.230 2.390 268.450 2.680 ;
        RECT 269.290 2.390 273.970 2.680 ;
        RECT 274.810 2.390 279.490 2.680 ;
        RECT 280.330 2.390 285.010 2.680 ;
        RECT 285.850 2.390 290.530 2.680 ;
        RECT 291.370 2.390 296.050 2.680 ;
        RECT 296.890 2.390 301.110 2.680 ;
        RECT 301.950 2.390 306.630 2.680 ;
        RECT 307.470 2.390 312.150 2.680 ;
        RECT 312.990 2.390 317.670 2.680 ;
        RECT 318.510 2.390 323.190 2.680 ;
        RECT 324.030 2.390 328.710 2.680 ;
        RECT 329.550 2.390 333.770 2.680 ;
        RECT 334.610 2.390 339.290 2.680 ;
        RECT 340.130 2.390 344.810 2.680 ;
        RECT 345.650 2.390 350.330 2.680 ;
        RECT 351.170 2.390 355.850 2.680 ;
        RECT 356.690 2.390 361.370 2.680 ;
        RECT 362.210 2.390 366.430 2.680 ;
        RECT 367.270 2.390 371.950 2.680 ;
        RECT 372.790 2.390 377.470 2.680 ;
        RECT 378.310 2.390 382.990 2.680 ;
        RECT 383.830 2.390 388.510 2.680 ;
        RECT 389.350 2.390 394.030 2.680 ;
        RECT 394.870 2.390 399.090 2.680 ;
        RECT 399.930 2.390 404.610 2.680 ;
        RECT 405.450 2.390 410.130 2.680 ;
        RECT 410.970 2.390 415.650 2.680 ;
        RECT 416.490 2.390 421.170 2.680 ;
        RECT 422.010 2.390 426.690 2.680 ;
        RECT 427.530 2.390 431.750 2.680 ;
        RECT 432.590 2.390 437.270 2.680 ;
        RECT 438.110 2.390 442.790 2.680 ;
        RECT 443.630 2.390 448.310 2.680 ;
        RECT 449.150 2.390 453.830 2.680 ;
        RECT 454.670 2.390 459.350 2.680 ;
        RECT 460.190 2.390 464.410 2.680 ;
        RECT 465.250 2.390 469.930 2.680 ;
        RECT 470.770 2.390 475.450 2.680 ;
        RECT 476.290 2.390 480.970 2.680 ;
        RECT 481.810 2.390 486.490 2.680 ;
        RECT 487.330 2.390 492.010 2.680 ;
        RECT 492.850 2.390 497.070 2.680 ;
        RECT 497.910 2.390 502.590 2.680 ;
        RECT 503.430 2.390 508.110 2.680 ;
        RECT 508.950 2.390 513.630 2.680 ;
        RECT 514.470 2.390 519.150 2.680 ;
        RECT 519.990 2.390 524.670 2.680 ;
        RECT 525.510 2.390 529.730 2.680 ;
        RECT 530.570 2.390 535.250 2.680 ;
        RECT 536.090 2.390 540.770 2.680 ;
        RECT 541.610 2.390 546.290 2.680 ;
        RECT 547.130 2.390 551.810 2.680 ;
        RECT 552.650 2.390 557.330 2.680 ;
        RECT 558.170 2.390 562.390 2.680 ;
        RECT 563.230 2.390 567.910 2.680 ;
        RECT 568.750 2.390 573.430 2.680 ;
        RECT 574.270 2.390 578.950 2.680 ;
        RECT 579.790 2.390 584.470 2.680 ;
        RECT 585.310 2.390 589.990 2.680 ;
        RECT 590.830 2.390 595.050 2.680 ;
        RECT 595.890 2.390 600.570 2.680 ;
        RECT 601.410 2.390 606.090 2.680 ;
        RECT 606.930 2.390 611.610 2.680 ;
        RECT 612.450 2.390 617.130 2.680 ;
        RECT 617.970 2.390 622.650 2.680 ;
        RECT 623.490 2.390 627.710 2.680 ;
        RECT 628.550 2.390 633.230 2.680 ;
        RECT 634.070 2.390 638.750 2.680 ;
        RECT 639.590 2.390 644.270 2.680 ;
        RECT 645.110 2.390 649.790 2.680 ;
        RECT 650.630 2.390 655.310 2.680 ;
        RECT 656.150 2.390 660.370 2.680 ;
        RECT 661.210 2.390 665.890 2.680 ;
        RECT 666.730 2.390 671.410 2.680 ;
        RECT 672.250 2.390 676.930 2.680 ;
        RECT 677.770 2.390 682.450 2.680 ;
        RECT 683.290 2.390 687.970 2.680 ;
        RECT 688.810 2.390 693.490 2.680 ;
        RECT 694.330 2.390 698.550 2.680 ;
        RECT 699.390 2.390 704.070 2.680 ;
        RECT 704.910 2.390 709.590 2.680 ;
        RECT 710.430 2.390 715.110 2.680 ;
        RECT 715.950 2.390 720.630 2.680 ;
        RECT 721.470 2.390 726.150 2.680 ;
        RECT 726.990 2.390 731.210 2.680 ;
        RECT 732.050 2.390 736.730 2.680 ;
        RECT 737.570 2.390 742.250 2.680 ;
        RECT 743.090 2.390 747.770 2.680 ;
        RECT 748.610 2.390 753.290 2.680 ;
        RECT 754.130 2.390 758.810 2.680 ;
        RECT 759.650 2.390 763.870 2.680 ;
        RECT 764.710 2.390 769.390 2.680 ;
        RECT 770.230 2.390 774.910 2.680 ;
        RECT 775.750 2.390 780.430 2.680 ;
        RECT 781.270 2.390 785.950 2.680 ;
        RECT 786.790 2.390 791.470 2.680 ;
        RECT 792.310 2.390 796.530 2.680 ;
        RECT 797.370 2.390 802.050 2.680 ;
        RECT 802.890 2.390 807.570 2.680 ;
        RECT 808.410 2.390 813.090 2.680 ;
        RECT 813.930 2.390 818.610 2.680 ;
        RECT 819.450 2.390 824.130 2.680 ;
        RECT 824.970 2.390 829.190 2.680 ;
        RECT 830.030 2.390 834.710 2.680 ;
        RECT 835.550 2.390 840.230 2.680 ;
        RECT 841.070 2.390 845.750 2.680 ;
        RECT 846.590 2.390 851.270 2.680 ;
        RECT 852.110 2.390 856.790 2.680 ;
        RECT 857.630 2.390 861.850 2.680 ;
        RECT 862.690 2.390 867.370 2.680 ;
        RECT 868.210 2.390 872.890 2.680 ;
        RECT 873.730 2.390 878.410 2.680 ;
        RECT 879.250 2.390 883.930 2.680 ;
        RECT 884.770 2.390 889.450 2.680 ;
        RECT 890.290 2.390 894.510 2.680 ;
        RECT 895.350 2.390 900.030 2.680 ;
        RECT 900.870 2.390 905.550 2.680 ;
        RECT 906.390 2.390 911.070 2.680 ;
        RECT 911.910 2.390 916.590 2.680 ;
        RECT 917.430 2.390 922.110 2.680 ;
        RECT 922.950 2.390 927.170 2.680 ;
        RECT 928.010 2.390 932.690 2.680 ;
        RECT 933.530 2.390 938.210 2.680 ;
        RECT 939.050 2.390 943.730 2.680 ;
        RECT 944.570 2.390 949.250 2.680 ;
        RECT 950.090 2.390 954.770 2.680 ;
        RECT 955.610 2.390 959.830 2.680 ;
        RECT 960.670 2.390 965.350 2.680 ;
        RECT 966.190 2.390 970.870 2.680 ;
        RECT 971.710 2.390 976.390 2.680 ;
        RECT 977.230 2.390 981.910 2.680 ;
        RECT 982.750 2.390 987.430 2.680 ;
        RECT 988.270 2.390 992.490 2.680 ;
        RECT 993.330 2.390 998.010 2.680 ;
        RECT 998.850 2.390 1003.530 2.680 ;
        RECT 1004.370 2.390 1009.050 2.680 ;
        RECT 1009.890 2.390 1014.570 2.680 ;
        RECT 1015.410 2.390 1020.090 2.680 ;
        RECT 1020.930 2.390 1025.150 2.680 ;
        RECT 1025.990 2.390 1030.670 2.680 ;
        RECT 1031.510 2.390 1036.190 2.680 ;
        RECT 1037.030 2.390 1041.710 2.680 ;
        RECT 1042.550 2.390 1047.230 2.680 ;
        RECT 1048.070 2.390 1052.750 2.680 ;
        RECT 1053.590 2.390 1057.810 2.680 ;
        RECT 1058.650 2.390 1063.330 2.680 ;
        RECT 1064.170 2.390 1068.850 2.680 ;
        RECT 1069.690 2.390 1074.370 2.680 ;
        RECT 1075.210 2.390 1079.890 2.680 ;
        RECT 1080.730 2.390 1085.410 2.680 ;
        RECT 1086.250 2.390 1090.470 2.680 ;
        RECT 1091.310 2.390 1095.990 2.680 ;
        RECT 1096.830 2.390 1101.510 2.680 ;
        RECT 1102.350 2.390 1107.030 2.680 ;
        RECT 1107.870 2.390 1112.550 2.680 ;
        RECT 1113.390 2.390 1118.070 2.680 ;
        RECT 1118.910 2.390 1123.130 2.680 ;
        RECT 1123.970 2.390 1128.650 2.680 ;
        RECT 1129.490 2.390 1134.170 2.680 ;
        RECT 1135.010 2.390 1139.690 2.680 ;
        RECT 1140.530 2.390 1145.210 2.680 ;
        RECT 1146.050 2.390 1150.730 2.680 ;
        RECT 1151.570 2.390 1155.790 2.680 ;
        RECT 1156.630 2.390 1161.310 2.680 ;
        RECT 1162.150 2.390 1166.830 2.680 ;
        RECT 1167.670 2.390 1172.350 2.680 ;
        RECT 1173.190 2.390 1177.870 2.680 ;
        RECT 1178.710 2.390 1183.390 2.680 ;
        RECT 1184.230 2.390 1188.450 2.680 ;
        RECT 1189.290 2.390 1193.970 2.680 ;
        RECT 1194.810 2.390 1199.490 2.680 ;
        RECT 1200.330 2.390 1205.010 2.680 ;
        RECT 1205.850 2.390 1210.530 2.680 ;
        RECT 1211.370 2.390 1216.050 2.680 ;
        RECT 1216.890 2.390 1221.110 2.680 ;
        RECT 1221.950 2.390 1226.630 2.680 ;
        RECT 1227.470 2.390 1232.150 2.680 ;
        RECT 1232.990 2.390 1237.670 2.680 ;
        RECT 1238.510 2.390 1243.190 2.680 ;
        RECT 1244.030 2.390 1248.710 2.680 ;
        RECT 1249.550 2.390 1253.770 2.680 ;
        RECT 1254.610 2.390 1259.290 2.680 ;
        RECT 1260.130 2.390 1264.810 2.680 ;
        RECT 1265.650 2.390 1270.330 2.680 ;
        RECT 1271.170 2.390 1275.850 2.680 ;
        RECT 1276.690 2.390 1281.370 2.680 ;
        RECT 1282.210 2.390 1286.430 2.680 ;
        RECT 1287.270 2.390 1291.950 2.680 ;
        RECT 1292.790 2.390 1297.470 2.680 ;
        RECT 1298.310 2.390 1302.990 2.680 ;
        RECT 1303.830 2.390 1308.510 2.680 ;
        RECT 1309.350 2.390 1314.030 2.680 ;
        RECT 1314.870 2.390 1319.090 2.680 ;
        RECT 1319.930 2.390 1324.610 2.680 ;
        RECT 1325.450 2.390 1330.130 2.680 ;
        RECT 1330.970 2.390 1335.650 2.680 ;
        RECT 1336.490 2.390 1341.170 2.680 ;
        RECT 1342.010 2.390 1346.690 2.680 ;
        RECT 1347.530 2.390 1352.210 2.680 ;
        RECT 1353.050 2.390 1357.270 2.680 ;
        RECT 1358.110 2.390 1362.790 2.680 ;
        RECT 1363.630 2.390 1368.310 2.680 ;
        RECT 1369.150 2.390 1373.830 2.680 ;
        RECT 1374.670 2.390 1379.350 2.680 ;
        RECT 1380.190 2.390 1384.870 2.680 ;
        RECT 1385.710 2.390 1389.930 2.680 ;
        RECT 1390.770 2.390 1395.450 2.680 ;
        RECT 1396.290 2.390 1400.970 2.680 ;
        RECT 1401.810 2.390 1406.490 2.680 ;
        RECT 1407.330 2.390 1412.010 2.680 ;
        RECT 1412.850 2.390 1417.530 2.680 ;
        RECT 1418.370 2.390 1422.590 2.680 ;
        RECT 1423.430 2.390 1428.110 2.680 ;
        RECT 1428.950 2.390 1433.630 2.680 ;
        RECT 1434.470 2.390 1439.150 2.680 ;
        RECT 1439.990 2.390 1444.670 2.680 ;
        RECT 1445.510 2.390 1450.190 2.680 ;
        RECT 1451.030 2.390 1455.250 2.680 ;
        RECT 1456.090 2.390 1460.770 2.680 ;
        RECT 1461.610 2.390 1466.290 2.680 ;
        RECT 1467.130 2.390 1471.810 2.680 ;
        RECT 1472.650 2.390 1477.330 2.680 ;
        RECT 1478.170 2.390 1482.850 2.680 ;
        RECT 1483.690 2.390 1487.910 2.680 ;
        RECT 1488.750 2.390 1493.430 2.680 ;
        RECT 1494.270 2.390 1498.950 2.680 ;
        RECT 1499.790 2.390 1504.470 2.680 ;
        RECT 1505.310 2.390 1509.990 2.680 ;
        RECT 1510.830 2.390 1515.510 2.680 ;
        RECT 1516.350 2.390 1520.570 2.680 ;
        RECT 1521.410 2.390 1526.090 2.680 ;
        RECT 1526.930 2.390 1531.610 2.680 ;
        RECT 1532.450 2.390 1537.130 2.680 ;
        RECT 1537.970 2.390 1542.650 2.680 ;
        RECT 1543.490 2.390 1548.170 2.680 ;
        RECT 1549.010 2.390 1553.230 2.680 ;
        RECT 1554.070 2.390 1558.750 2.680 ;
        RECT 1559.590 2.390 1564.270 2.680 ;
        RECT 1565.110 2.390 1569.790 2.680 ;
        RECT 1570.630 2.390 1575.310 2.680 ;
        RECT 1576.150 2.390 1580.830 2.680 ;
        RECT 1581.670 2.390 1585.890 2.680 ;
        RECT 1586.730 2.390 1591.410 2.680 ;
        RECT 1592.250 2.390 1596.930 2.680 ;
        RECT 1597.770 2.390 1602.450 2.680 ;
        RECT 1603.290 2.390 1607.970 2.680 ;
        RECT 1608.810 2.390 1613.490 2.680 ;
        RECT 1614.330 2.390 1618.550 2.680 ;
        RECT 1619.390 2.390 1624.070 2.680 ;
        RECT 1624.910 2.390 1629.590 2.680 ;
        RECT 1630.430 2.390 1635.110 2.680 ;
        RECT 1635.950 2.390 1640.630 2.680 ;
        RECT 1641.470 2.390 1646.150 2.680 ;
        RECT 1646.990 2.390 1651.210 2.680 ;
        RECT 1652.050 2.390 1656.730 2.680 ;
        RECT 1657.570 2.390 1662.250 2.680 ;
        RECT 1663.090 2.390 1667.770 2.680 ;
        RECT 1668.610 2.390 1673.290 2.680 ;
        RECT 1674.130 2.390 1678.810 2.680 ;
        RECT 1679.650 2.390 1683.870 2.680 ;
        RECT 1684.710 2.390 1689.390 2.680 ;
        RECT 1690.230 2.390 1694.910 2.680 ;
        RECT 1695.750 2.390 1700.430 2.680 ;
        RECT 1701.270 2.390 1705.950 2.680 ;
        RECT 1706.790 2.390 1711.470 2.680 ;
        RECT 1712.310 2.390 1716.530 2.680 ;
        RECT 1717.370 2.390 1722.050 2.680 ;
        RECT 1722.890 2.390 1727.570 2.680 ;
        RECT 1728.410 2.390 1733.090 2.680 ;
        RECT 1733.930 2.390 1738.610 2.680 ;
        RECT 1739.450 2.390 1744.130 2.680 ;
        RECT 1744.970 2.390 1749.190 2.680 ;
        RECT 1750.030 2.390 1754.710 2.680 ;
        RECT 1755.550 2.390 1760.230 2.680 ;
        RECT 1761.070 2.390 1765.750 2.680 ;
        RECT 1766.590 2.390 1771.270 2.680 ;
        RECT 1772.110 2.390 1776.790 2.680 ;
        RECT 1777.630 2.390 1781.850 2.680 ;
        RECT 1782.690 2.390 1787.370 2.680 ;
        RECT 1788.210 2.390 1792.890 2.680 ;
        RECT 1793.730 2.390 1798.410 2.680 ;
        RECT 1799.250 2.390 1803.930 2.680 ;
        RECT 1804.770 2.390 1809.450 2.680 ;
        RECT 1810.290 2.390 1814.510 2.680 ;
        RECT 1815.350 2.390 1820.030 2.680 ;
        RECT 1820.870 2.390 1825.550 2.680 ;
        RECT 1826.390 2.390 1831.070 2.680 ;
        RECT 1831.910 2.390 1836.590 2.680 ;
        RECT 1837.430 2.390 1842.110 2.680 ;
        RECT 1842.950 2.390 1847.170 2.680 ;
        RECT 1848.010 2.390 1852.690 2.680 ;
        RECT 1853.530 2.390 1858.210 2.680 ;
        RECT 1859.050 2.390 1863.730 2.680 ;
        RECT 1864.570 2.390 1869.250 2.680 ;
        RECT 1870.090 2.390 1874.770 2.680 ;
        RECT 1875.610 2.390 1879.830 2.680 ;
        RECT 1880.670 2.390 1885.350 2.680 ;
        RECT 1886.190 2.390 1890.870 2.680 ;
        RECT 1891.710 2.390 1896.390 2.680 ;
        RECT 1897.230 2.390 1901.910 2.680 ;
        RECT 1902.750 2.390 1907.430 2.680 ;
        RECT 1908.270 2.390 1912.490 2.680 ;
        RECT 1913.330 2.390 1918.010 2.680 ;
        RECT 1918.850 2.390 1923.530 2.680 ;
        RECT 1924.370 2.390 1929.050 2.680 ;
        RECT 1929.890 2.390 1934.570 2.680 ;
        RECT 1935.410 2.390 1940.090 2.680 ;
        RECT 1940.930 2.390 1945.150 2.680 ;
        RECT 1945.990 2.390 1950.670 2.680 ;
        RECT 1951.510 2.390 1956.190 2.680 ;
        RECT 1957.030 2.390 1961.710 2.680 ;
        RECT 1962.550 2.390 1967.230 2.680 ;
        RECT 1968.070 2.390 1972.750 2.680 ;
        RECT 1973.590 2.390 1977.810 2.680 ;
        RECT 1978.650 2.390 1983.330 2.680 ;
        RECT 1984.170 2.390 1988.850 2.680 ;
        RECT 1989.690 2.390 1994.370 2.680 ;
        RECT 1995.210 2.390 1999.890 2.680 ;
        RECT 2000.730 2.390 2005.410 2.680 ;
        RECT 2006.250 2.390 2010.470 2.680 ;
        RECT 2011.310 2.390 2015.990 2.680 ;
        RECT 2016.830 2.390 2021.510 2.680 ;
        RECT 2022.350 2.390 2027.030 2.680 ;
        RECT 2027.870 2.390 2032.550 2.680 ;
        RECT 2033.390 2.390 2038.070 2.680 ;
        RECT 2038.910 2.390 2043.590 2.680 ;
        RECT 2044.430 2.390 2048.650 2.680 ;
        RECT 2049.490 2.390 2054.170 2.680 ;
        RECT 2055.010 2.390 2059.690 2.680 ;
        RECT 2060.530 2.390 2065.210 2.680 ;
        RECT 2066.050 2.390 2070.730 2.680 ;
        RECT 2071.570 2.390 2076.250 2.680 ;
        RECT 2077.090 2.390 2081.310 2.680 ;
        RECT 2082.150 2.390 2086.830 2.680 ;
        RECT 2087.670 2.390 2092.350 2.680 ;
        RECT 2093.190 2.390 2097.870 2.680 ;
        RECT 2098.710 2.390 2103.390 2.680 ;
        RECT 2104.230 2.390 2108.910 2.680 ;
        RECT 2109.750 2.390 2113.970 2.680 ;
        RECT 2114.810 2.390 2119.490 2.680 ;
        RECT 2120.330 2.390 2125.010 2.680 ;
        RECT 2125.850 2.390 2130.530 2.680 ;
        RECT 2131.370 2.390 2136.050 2.680 ;
        RECT 2136.890 2.390 2141.570 2.680 ;
        RECT 2142.410 2.390 2146.630 2.680 ;
        RECT 2147.470 2.390 2152.150 2.680 ;
        RECT 2152.990 2.390 2157.670 2.680 ;
        RECT 2158.510 2.390 2163.190 2.680 ;
        RECT 2164.030 2.390 2168.710 2.680 ;
        RECT 2169.550 2.390 2174.230 2.680 ;
        RECT 2175.070 2.390 2179.290 2.680 ;
        RECT 2180.130 2.390 2184.810 2.680 ;
        RECT 2185.650 2.390 2190.330 2.680 ;
        RECT 2191.170 2.390 2195.850 2.680 ;
        RECT 2196.690 2.390 2201.370 2.680 ;
        RECT 2202.210 2.390 2206.890 2.680 ;
        RECT 2207.730 2.390 2211.950 2.680 ;
        RECT 2212.790 2.390 2217.470 2.680 ;
        RECT 2218.310 2.390 2222.990 2.680 ;
        RECT 2223.830 2.390 2228.510 2.680 ;
        RECT 2229.350 2.390 2234.030 2.680 ;
        RECT 2234.870 2.390 2239.550 2.680 ;
        RECT 2240.390 2.390 2244.610 2.680 ;
        RECT 2245.450 2.390 2250.130 2.680 ;
        RECT 2250.970 2.390 2255.650 2.680 ;
        RECT 2256.490 2.390 2261.170 2.680 ;
        RECT 2262.010 2.390 2266.690 2.680 ;
        RECT 2267.530 2.390 2272.210 2.680 ;
        RECT 2273.050 2.390 2277.270 2.680 ;
        RECT 2278.110 2.390 2282.790 2.680 ;
        RECT 2283.630 2.390 2288.310 2.680 ;
        RECT 2289.150 2.390 2293.830 2.680 ;
        RECT 2294.670 2.390 2299.350 2.680 ;
        RECT 2300.190 2.390 2304.870 2.680 ;
        RECT 2305.710 2.390 2309.930 2.680 ;
        RECT 2310.770 2.390 2315.450 2.680 ;
        RECT 2316.290 2.390 2320.970 2.680 ;
        RECT 2321.810 2.390 2326.490 2.680 ;
        RECT 2327.330 2.390 2332.010 2.680 ;
        RECT 2332.850 2.390 2337.530 2.680 ;
        RECT 2338.370 2.390 2342.590 2.680 ;
        RECT 2343.430 2.390 2348.110 2.680 ;
        RECT 2348.950 2.390 2353.630 2.680 ;
        RECT 2354.470 2.390 2359.150 2.680 ;
        RECT 2359.990 2.390 2364.670 2.680 ;
        RECT 2365.510 2.390 2370.190 2.680 ;
        RECT 2371.030 2.390 2375.250 2.680 ;
        RECT 2376.090 2.390 2380.770 2.680 ;
        RECT 2381.610 2.390 2386.290 2.680 ;
        RECT 2387.130 2.390 2391.810 2.680 ;
        RECT 2392.650 2.390 2397.330 2.680 ;
        RECT 2398.170 2.390 2402.850 2.680 ;
        RECT 2403.690 2.390 2407.910 2.680 ;
        RECT 2408.750 2.390 2413.430 2.680 ;
        RECT 2414.270 2.390 2418.950 2.680 ;
        RECT 2419.790 2.390 2424.470 2.680 ;
        RECT 2425.310 2.390 2429.990 2.680 ;
        RECT 2430.830 2.390 2435.510 2.680 ;
        RECT 2436.350 2.390 2440.570 2.680 ;
        RECT 2441.410 2.390 2446.090 2.680 ;
        RECT 2446.930 2.390 2451.610 2.680 ;
        RECT 2452.450 2.390 2457.130 2.680 ;
        RECT 2457.970 2.390 2462.650 2.680 ;
        RECT 2463.490 2.390 2468.170 2.680 ;
        RECT 2469.010 2.390 2473.230 2.680 ;
        RECT 2474.070 2.390 2478.750 2.680 ;
        RECT 2479.590 2.390 2484.270 2.680 ;
        RECT 2485.110 2.390 2489.790 2.680 ;
        RECT 2490.630 2.390 2495.310 2.680 ;
        RECT 2496.150 2.390 2500.830 2.680 ;
        RECT 2501.670 2.390 2505.890 2.680 ;
        RECT 2506.730 2.390 2511.410 2.680 ;
        RECT 2512.250 2.390 2516.930 2.680 ;
        RECT 2517.770 2.390 2522.450 2.680 ;
        RECT 2523.290 2.390 2527.970 2.680 ;
        RECT 2528.810 2.390 2533.490 2.680 ;
        RECT 2534.330 2.390 2538.550 2.680 ;
        RECT 2539.390 2.390 2544.070 2.680 ;
        RECT 2544.910 2.390 2549.590 2.680 ;
        RECT 2550.430 2.390 2555.110 2.680 ;
        RECT 2555.950 2.390 2560.630 2.680 ;
        RECT 2561.470 2.390 2566.150 2.680 ;
        RECT 2566.990 2.390 2571.210 2.680 ;
        RECT 2572.050 2.390 2576.730 2.680 ;
        RECT 2577.570 2.390 2582.250 2.680 ;
        RECT 2583.090 2.390 2587.770 2.680 ;
        RECT 2588.610 2.390 2593.290 2.680 ;
        RECT 2594.130 2.390 2598.810 2.680 ;
        RECT 2599.650 2.390 2603.870 2.680 ;
        RECT 2604.710 2.390 2609.390 2.680 ;
        RECT 2610.230 2.390 2614.910 2.680 ;
        RECT 2615.750 2.390 2620.430 2.680 ;
        RECT 2621.270 2.390 2625.950 2.680 ;
        RECT 2626.790 2.390 2631.470 2.680 ;
        RECT 2632.310 2.390 2636.530 2.680 ;
        RECT 2637.370 2.390 2642.050 2.680 ;
        RECT 2642.890 2.390 2647.570 2.680 ;
        RECT 2648.410 2.390 2653.090 2.680 ;
        RECT 2653.930 2.390 2658.610 2.680 ;
        RECT 2659.450 2.390 2664.130 2.680 ;
        RECT 2664.970 2.390 2669.190 2.680 ;
        RECT 2670.030 2.390 2674.710 2.680 ;
        RECT 2675.550 2.390 2680.230 2.680 ;
        RECT 2681.070 2.390 2685.750 2.680 ;
        RECT 2686.590 2.390 2689.070 2.680 ;
      LAYER met3 ;
        RECT 2.400 3667.600 2697.600 3688.485 ;
        RECT 2.800 3666.920 2697.600 3667.600 ;
        RECT 2.800 3666.200 2697.200 3666.920 ;
        RECT 2.400 3665.520 2697.200 3666.200 ;
        RECT 2.400 3603.000 2697.600 3665.520 ;
        RECT 2.800 3601.600 2697.600 3603.000 ;
        RECT 2.400 3600.960 2697.600 3601.600 ;
        RECT 2.400 3599.560 2697.200 3600.960 ;
        RECT 2.400 3537.720 2697.600 3599.560 ;
        RECT 2.800 3536.320 2697.600 3537.720 ;
        RECT 2.400 3535.000 2697.600 3536.320 ;
        RECT 2.400 3533.600 2697.200 3535.000 ;
        RECT 2.400 3473.120 2697.600 3533.600 ;
        RECT 2.800 3471.720 2697.600 3473.120 ;
        RECT 2.400 3469.040 2697.600 3471.720 ;
        RECT 2.400 3467.640 2697.200 3469.040 ;
        RECT 2.400 3407.840 2697.600 3467.640 ;
        RECT 2.800 3406.440 2697.600 3407.840 ;
        RECT 2.400 3403.080 2697.600 3406.440 ;
        RECT 2.400 3401.680 2697.200 3403.080 ;
        RECT 2.400 3343.240 2697.600 3401.680 ;
        RECT 2.800 3341.840 2697.600 3343.240 ;
        RECT 2.400 3337.120 2697.600 3341.840 ;
        RECT 2.400 3335.720 2697.200 3337.120 ;
        RECT 2.400 3277.960 2697.600 3335.720 ;
        RECT 2.800 3276.560 2697.600 3277.960 ;
        RECT 2.400 3270.480 2697.600 3276.560 ;
        RECT 2.400 3269.080 2697.200 3270.480 ;
        RECT 2.400 3213.360 2697.600 3269.080 ;
        RECT 2.800 3211.960 2697.600 3213.360 ;
        RECT 2.400 3204.520 2697.600 3211.960 ;
        RECT 2.400 3203.120 2697.200 3204.520 ;
        RECT 2.400 3148.080 2697.600 3203.120 ;
        RECT 2.800 3146.680 2697.600 3148.080 ;
        RECT 2.400 3138.560 2697.600 3146.680 ;
        RECT 2.400 3137.160 2697.200 3138.560 ;
        RECT 2.400 3083.480 2697.600 3137.160 ;
        RECT 2.800 3082.080 2697.600 3083.480 ;
        RECT 2.400 3072.600 2697.600 3082.080 ;
        RECT 2.400 3071.200 2697.200 3072.600 ;
        RECT 2.400 3018.200 2697.600 3071.200 ;
        RECT 2.800 3016.800 2697.600 3018.200 ;
        RECT 2.400 3006.640 2697.600 3016.800 ;
        RECT 2.400 3005.240 2697.200 3006.640 ;
        RECT 2.400 2953.600 2697.600 3005.240 ;
        RECT 2.800 2952.200 2697.600 2953.600 ;
        RECT 2.400 2940.680 2697.600 2952.200 ;
        RECT 2.400 2939.280 2697.200 2940.680 ;
        RECT 2.400 2889.000 2697.600 2939.280 ;
        RECT 2.800 2887.600 2697.600 2889.000 ;
        RECT 2.400 2874.040 2697.600 2887.600 ;
        RECT 2.400 2872.640 2697.200 2874.040 ;
        RECT 2.400 2823.720 2697.600 2872.640 ;
        RECT 2.800 2822.320 2697.600 2823.720 ;
        RECT 2.400 2808.080 2697.600 2822.320 ;
        RECT 2.400 2806.680 2697.200 2808.080 ;
        RECT 2.400 2759.120 2697.600 2806.680 ;
        RECT 2.800 2757.720 2697.600 2759.120 ;
        RECT 2.400 2742.120 2697.600 2757.720 ;
        RECT 2.400 2740.720 2697.200 2742.120 ;
        RECT 2.400 2693.840 2697.600 2740.720 ;
        RECT 2.800 2692.440 2697.600 2693.840 ;
        RECT 2.400 2676.160 2697.600 2692.440 ;
        RECT 2.400 2674.760 2697.200 2676.160 ;
        RECT 2.400 2629.240 2697.600 2674.760 ;
        RECT 2.800 2627.840 2697.600 2629.240 ;
        RECT 2.400 2610.200 2697.600 2627.840 ;
        RECT 2.400 2608.800 2697.200 2610.200 ;
        RECT 2.400 2563.960 2697.600 2608.800 ;
        RECT 2.800 2562.560 2697.600 2563.960 ;
        RECT 2.400 2544.240 2697.600 2562.560 ;
        RECT 2.400 2542.840 2697.200 2544.240 ;
        RECT 2.400 2499.360 2697.600 2542.840 ;
        RECT 2.800 2497.960 2697.600 2499.360 ;
        RECT 2.400 2477.600 2697.600 2497.960 ;
        RECT 2.400 2476.200 2697.200 2477.600 ;
        RECT 2.400 2434.080 2697.600 2476.200 ;
        RECT 2.800 2432.680 2697.600 2434.080 ;
        RECT 2.400 2411.640 2697.600 2432.680 ;
        RECT 2.400 2410.240 2697.200 2411.640 ;
        RECT 2.400 2369.480 2697.600 2410.240 ;
        RECT 2.800 2368.080 2697.600 2369.480 ;
        RECT 2.400 2345.680 2697.600 2368.080 ;
        RECT 2.400 2344.280 2697.200 2345.680 ;
        RECT 2.400 2304.200 2697.600 2344.280 ;
        RECT 2.800 2302.800 2697.600 2304.200 ;
        RECT 2.400 2279.720 2697.600 2302.800 ;
        RECT 2.400 2278.320 2697.200 2279.720 ;
        RECT 2.400 2239.600 2697.600 2278.320 ;
        RECT 2.800 2238.200 2697.600 2239.600 ;
        RECT 2.400 2213.760 2697.600 2238.200 ;
        RECT 2.400 2212.360 2697.200 2213.760 ;
        RECT 2.400 2175.000 2697.600 2212.360 ;
        RECT 2.800 2173.600 2697.600 2175.000 ;
        RECT 2.400 2147.800 2697.600 2173.600 ;
        RECT 2.400 2146.400 2697.200 2147.800 ;
        RECT 2.400 2109.720 2697.600 2146.400 ;
        RECT 2.800 2108.320 2697.600 2109.720 ;
        RECT 2.400 2081.160 2697.600 2108.320 ;
        RECT 2.400 2079.760 2697.200 2081.160 ;
        RECT 2.400 2045.120 2697.600 2079.760 ;
        RECT 2.800 2043.720 2697.600 2045.120 ;
        RECT 2.400 2015.200 2697.600 2043.720 ;
        RECT 2.400 2013.800 2697.200 2015.200 ;
        RECT 2.400 1979.840 2697.600 2013.800 ;
        RECT 2.800 1978.440 2697.600 1979.840 ;
        RECT 2.400 1949.240 2697.600 1978.440 ;
        RECT 2.400 1947.840 2697.200 1949.240 ;
        RECT 2.400 1915.240 2697.600 1947.840 ;
        RECT 2.800 1913.840 2697.600 1915.240 ;
        RECT 2.400 1883.280 2697.600 1913.840 ;
        RECT 2.400 1881.880 2697.200 1883.280 ;
        RECT 2.400 1849.960 2697.600 1881.880 ;
        RECT 2.800 1848.560 2697.600 1849.960 ;
        RECT 2.400 1817.320 2697.600 1848.560 ;
        RECT 2.400 1815.920 2697.200 1817.320 ;
        RECT 2.400 1785.360 2697.600 1815.920 ;
        RECT 2.800 1783.960 2697.600 1785.360 ;
        RECT 2.400 1751.360 2697.600 1783.960 ;
        RECT 2.400 1749.960 2697.200 1751.360 ;
        RECT 2.400 1720.080 2697.600 1749.960 ;
        RECT 2.800 1718.680 2697.600 1720.080 ;
        RECT 2.400 1685.400 2697.600 1718.680 ;
        RECT 2.400 1684.000 2697.200 1685.400 ;
        RECT 2.400 1655.480 2697.600 1684.000 ;
        RECT 2.800 1654.080 2697.600 1655.480 ;
        RECT 2.400 1618.760 2697.600 1654.080 ;
        RECT 2.400 1617.360 2697.200 1618.760 ;
        RECT 2.400 1590.200 2697.600 1617.360 ;
        RECT 2.800 1588.800 2697.600 1590.200 ;
        RECT 2.400 1552.800 2697.600 1588.800 ;
        RECT 2.400 1551.400 2697.200 1552.800 ;
        RECT 2.400 1525.600 2697.600 1551.400 ;
        RECT 2.800 1524.200 2697.600 1525.600 ;
        RECT 2.400 1486.840 2697.600 1524.200 ;
        RECT 2.400 1485.440 2697.200 1486.840 ;
        RECT 2.400 1461.000 2697.600 1485.440 ;
        RECT 2.800 1459.600 2697.600 1461.000 ;
        RECT 2.400 1420.880 2697.600 1459.600 ;
        RECT 2.400 1419.480 2697.200 1420.880 ;
        RECT 2.400 1395.720 2697.600 1419.480 ;
        RECT 2.800 1394.320 2697.600 1395.720 ;
        RECT 2.400 1354.920 2697.600 1394.320 ;
        RECT 2.400 1353.520 2697.200 1354.920 ;
        RECT 2.400 1331.120 2697.600 1353.520 ;
        RECT 2.800 1329.720 2697.600 1331.120 ;
        RECT 2.400 1288.960 2697.600 1329.720 ;
        RECT 2.400 1287.560 2697.200 1288.960 ;
        RECT 2.400 1265.840 2697.600 1287.560 ;
        RECT 2.800 1264.440 2697.600 1265.840 ;
        RECT 2.400 1222.320 2697.600 1264.440 ;
        RECT 2.400 1220.920 2697.200 1222.320 ;
        RECT 2.400 1201.240 2697.600 1220.920 ;
        RECT 2.800 1199.840 2697.600 1201.240 ;
        RECT 2.400 1156.360 2697.600 1199.840 ;
        RECT 2.400 1154.960 2697.200 1156.360 ;
        RECT 2.400 1135.960 2697.600 1154.960 ;
        RECT 2.800 1134.560 2697.600 1135.960 ;
        RECT 2.400 1090.400 2697.600 1134.560 ;
        RECT 2.400 1089.000 2697.200 1090.400 ;
        RECT 2.400 1071.360 2697.600 1089.000 ;
        RECT 2.800 1069.960 2697.600 1071.360 ;
        RECT 2.400 1024.440 2697.600 1069.960 ;
        RECT 2.400 1023.040 2697.200 1024.440 ;
        RECT 2.400 1006.080 2697.600 1023.040 ;
        RECT 2.800 1004.680 2697.600 1006.080 ;
        RECT 2.400 958.480 2697.600 1004.680 ;
        RECT 2.400 957.080 2697.200 958.480 ;
        RECT 2.400 941.480 2697.600 957.080 ;
        RECT 2.800 940.080 2697.600 941.480 ;
        RECT 2.400 892.520 2697.600 940.080 ;
        RECT 2.400 891.120 2697.200 892.520 ;
        RECT 2.400 876.200 2697.600 891.120 ;
        RECT 2.800 874.800 2697.600 876.200 ;
        RECT 2.400 825.880 2697.600 874.800 ;
        RECT 2.400 824.480 2697.200 825.880 ;
        RECT 2.400 811.600 2697.600 824.480 ;
        RECT 2.800 810.200 2697.600 811.600 ;
        RECT 2.400 759.920 2697.600 810.200 ;
        RECT 2.400 758.520 2697.200 759.920 ;
        RECT 2.400 747.000 2697.600 758.520 ;
        RECT 2.800 745.600 2697.600 747.000 ;
        RECT 2.400 693.960 2697.600 745.600 ;
        RECT 2.400 692.560 2697.200 693.960 ;
        RECT 2.400 681.720 2697.600 692.560 ;
        RECT 2.800 680.320 2697.600 681.720 ;
        RECT 2.400 628.000 2697.600 680.320 ;
        RECT 2.400 626.600 2697.200 628.000 ;
        RECT 2.400 617.120 2697.600 626.600 ;
        RECT 2.800 615.720 2697.600 617.120 ;
        RECT 2.400 562.040 2697.600 615.720 ;
        RECT 2.400 560.640 2697.200 562.040 ;
        RECT 2.400 551.840 2697.600 560.640 ;
        RECT 2.800 550.440 2697.600 551.840 ;
        RECT 2.400 496.080 2697.600 550.440 ;
        RECT 2.400 494.680 2697.200 496.080 ;
        RECT 2.400 487.240 2697.600 494.680 ;
        RECT 2.800 485.840 2697.600 487.240 ;
        RECT 2.400 429.440 2697.600 485.840 ;
        RECT 2.400 428.040 2697.200 429.440 ;
        RECT 2.400 421.960 2697.600 428.040 ;
        RECT 2.800 420.560 2697.600 421.960 ;
        RECT 2.400 363.480 2697.600 420.560 ;
        RECT 2.400 362.080 2697.200 363.480 ;
        RECT 2.400 357.360 2697.600 362.080 ;
        RECT 2.800 355.960 2697.600 357.360 ;
        RECT 2.400 297.520 2697.600 355.960 ;
        RECT 2.400 296.120 2697.200 297.520 ;
        RECT 2.400 292.080 2697.600 296.120 ;
        RECT 2.800 290.680 2697.600 292.080 ;
        RECT 2.400 231.560 2697.600 290.680 ;
        RECT 2.400 230.160 2697.200 231.560 ;
        RECT 2.400 227.480 2697.600 230.160 ;
        RECT 2.800 226.080 2697.600 227.480 ;
        RECT 2.400 165.600 2697.600 226.080 ;
        RECT 2.400 164.200 2697.200 165.600 ;
        RECT 2.400 162.200 2697.600 164.200 ;
        RECT 2.800 160.800 2697.600 162.200 ;
        RECT 2.400 99.640 2697.600 160.800 ;
        RECT 2.400 98.240 2697.200 99.640 ;
        RECT 2.400 97.600 2697.600 98.240 ;
        RECT 2.800 96.200 2697.600 97.600 ;
        RECT 2.400 33.680 2697.600 96.200 ;
        RECT 2.400 33.000 2697.200 33.680 ;
        RECT 2.800 32.280 2697.200 33.000 ;
        RECT 2.800 31.600 2697.600 32.280 ;
        RECT 2.400 10.715 2697.600 31.600 ;
      LAYER met4 ;
        RECT 21.040 10.640 2633.840 3688.560 ;
      LAYER met5 ;
        RECT 5.520 179.670 2694.220 3627.820 ;
  END
END user_project_wrapper
END LIBRARY

